magic
tech gf180mcuD
magscale 1 10
timestamp 1701971416
<< metal2 >>
rect 11032 595672 11256 597000
rect 33096 595672 33320 597000
rect 55160 595672 55384 597000
rect 11004 595560 11256 595672
rect 33068 595560 33320 595672
rect 55132 595560 55384 595672
rect 77224 595560 77448 597000
rect 99288 595672 99512 597000
rect 121352 595672 121576 597000
rect 143416 595672 143640 597000
rect 99288 595560 99540 595672
rect 121352 595560 121604 595672
rect 4172 460180 4228 460190
rect 4172 420028 4228 460124
rect 4172 419972 4340 420028
rect 4172 417844 4228 417854
rect 4172 415828 4228 417788
rect 4172 415762 4228 415772
rect 4284 410788 4340 419972
rect 4284 410722 4340 410732
rect 10892 389956 10948 389966
rect 4172 333172 4228 333182
rect 4172 322532 4228 333116
rect 4172 322466 4228 322476
rect 4172 297556 4228 297566
rect 4172 291060 4228 297500
rect 4172 290994 4228 291004
rect 4172 208740 4228 208750
rect 4172 121716 4228 208684
rect 4172 121650 4228 121660
rect 4172 79156 4228 79166
rect 4172 50372 4228 79100
rect 4172 50306 4228 50316
rect 4396 49700 4452 49710
rect 4396 36932 4452 49644
rect 4396 36866 4452 36876
rect 10892 22932 10948 389900
rect 11004 311668 11060 595560
rect 12572 488404 12628 488414
rect 12572 402724 12628 488348
rect 15932 415828 15988 415838
rect 15932 407876 15988 415772
rect 15932 407810 15988 407820
rect 12572 402658 12628 402668
rect 33068 390628 33124 595560
rect 55132 409892 55188 595560
rect 77308 570388 77364 595560
rect 99484 590548 99540 595560
rect 121548 590660 121604 595560
rect 143388 595560 143640 595672
rect 165480 595672 165704 597000
rect 187544 595672 187768 597000
rect 209608 595672 209832 597000
rect 231672 595672 231896 597000
rect 253736 595672 253960 597000
rect 275800 595672 276024 597000
rect 297864 595672 298088 597000
rect 319928 595672 320152 597000
rect 341992 595672 342216 597000
rect 364056 595672 364280 597000
rect 386120 595672 386344 597000
rect 165480 595560 165732 595672
rect 187544 595560 187796 595672
rect 121548 590594 121604 590604
rect 136892 590660 136948 590670
rect 99484 590482 99540 590492
rect 77308 570322 77364 570332
rect 55132 409826 55188 409836
rect 56252 530740 56308 530750
rect 56252 404180 56308 530684
rect 136892 409780 136948 590604
rect 136892 409714 136948 409724
rect 56252 404114 56308 404124
rect 111692 402612 111748 402622
rect 106652 393428 106708 393438
rect 103292 393316 103348 393326
rect 33068 390562 33124 390572
rect 40908 393204 40964 393214
rect 31052 386820 31108 386830
rect 11004 311602 11060 311612
rect 14252 386708 14308 386718
rect 10892 22866 10948 22876
rect 13244 222740 13300 222750
rect 11564 5908 11620 5918
rect 11564 480 11620 5852
rect 11368 392 11620 480
rect 13244 480 13300 222684
rect 14252 192052 14308 386652
rect 24668 242676 24724 242686
rect 14252 191986 14308 191996
rect 15148 229348 15204 229358
rect 15148 480 15204 229292
rect 17052 227668 17108 227678
rect 17052 480 17108 227612
rect 22764 224420 22820 224430
rect 18956 222628 19012 222638
rect 18956 480 19012 222572
rect 20860 217588 20916 217598
rect 20860 480 20916 217532
rect 22764 480 22820 224364
rect 24668 480 24724 242620
rect 26572 212548 26628 212558
rect 26572 480 26628 212492
rect 30380 210868 30436 210878
rect 30380 480 30436 210812
rect 31052 107380 31108 386764
rect 34412 385476 34468 385486
rect 34412 276724 34468 385420
rect 34412 276658 34468 276668
rect 40236 383908 40292 383918
rect 40236 238308 40292 383852
rect 40908 242004 40964 393148
rect 100156 391636 100212 391646
rect 99932 391524 99988 391534
rect 41132 384132 41188 384142
rect 40908 241938 40964 241948
rect 41020 384020 41076 384030
rect 41020 238532 41076 383964
rect 41132 255388 41188 384076
rect 62412 383124 62468 383134
rect 62412 299880 62468 383068
rect 77420 303268 77476 303278
rect 77420 299880 77476 303212
rect 92428 301588 92484 301598
rect 92428 299880 92484 301532
rect 47404 299348 47460 299358
rect 47404 299282 47460 299292
rect 41132 255332 41524 255388
rect 41468 240548 41524 255332
rect 41580 242004 41636 242014
rect 41636 241948 41748 242004
rect 41580 241938 41636 241948
rect 41692 240548 41748 241948
rect 50764 240772 50820 240782
rect 50764 240706 50820 240716
rect 44156 240548 44212 240558
rect 54796 240548 54852 240558
rect 41692 240492 42728 240548
rect 44212 240492 44744 240548
rect 41468 240482 41524 240492
rect 44156 240482 44212 240492
rect 54796 240482 54852 240492
rect 58828 240436 58884 240446
rect 58828 240370 58884 240380
rect 62860 240324 62916 240334
rect 62860 240258 62916 240268
rect 52780 240212 52836 240222
rect 52780 240146 52836 240156
rect 60844 240212 60900 240222
rect 60844 240146 60900 240156
rect 56812 240100 56868 240110
rect 41020 238466 41076 238476
rect 46732 238532 46788 240072
rect 46732 238466 46788 238476
rect 40236 238242 40292 238252
rect 48748 238308 48804 240072
rect 56812 240034 56868 240044
rect 64876 239764 64932 240072
rect 64876 239698 64932 239708
rect 48748 238242 48804 238252
rect 66892 236852 66948 240072
rect 66892 236786 66948 236796
rect 38556 236068 38612 236078
rect 31052 107314 31108 107324
rect 32284 234500 32340 234510
rect 32284 480 32340 234444
rect 37996 232820 38052 232830
rect 34188 224308 34244 224318
rect 34188 480 34244 224252
rect 37996 480 38052 232764
rect 38444 227780 38500 227790
rect 38444 4900 38500 227724
rect 38444 4834 38500 4844
rect 38556 4228 38612 236012
rect 68908 235172 68964 240072
rect 70924 236628 70980 240072
rect 70924 236562 70980 236572
rect 68908 235106 68964 235116
rect 72940 235060 72996 240072
rect 74956 238532 75012 240072
rect 74956 238466 75012 238476
rect 76972 238532 77028 240072
rect 78988 239876 79044 240072
rect 78988 239810 79044 239820
rect 76972 238466 77028 238476
rect 81004 237860 81060 240072
rect 81004 237794 81060 237804
rect 83020 237636 83076 240072
rect 85036 237972 85092 240072
rect 87052 238084 87108 240072
rect 89068 238196 89124 240072
rect 91084 238532 91140 240072
rect 91084 238466 91140 238476
rect 93100 238420 93156 240072
rect 93100 238354 93156 238364
rect 95116 238420 95172 240072
rect 95116 238354 95172 238364
rect 89068 238130 89124 238140
rect 97132 238196 97188 240072
rect 99820 238644 99876 238654
rect 99820 238308 99876 238588
rect 99932 238532 99988 391468
rect 99932 238466 99988 238476
rect 99820 238242 99876 238252
rect 97132 238130 97188 238140
rect 87052 238018 87108 238028
rect 85036 237906 85092 237916
rect 100156 237748 100212 391580
rect 100156 237682 100212 237692
rect 100380 390068 100436 390078
rect 83020 237570 83076 237580
rect 100380 237636 100436 390012
rect 102508 257124 102564 257134
rect 102508 255332 102564 257068
rect 102508 255266 102564 255276
rect 103292 238308 103348 393260
rect 104972 390180 105028 390190
rect 103404 286468 103460 286478
rect 103404 266980 103460 286412
rect 103516 285348 103572 285358
rect 103516 272804 103572 285292
rect 103516 272738 103572 272748
rect 103404 266914 103460 266924
rect 103292 238242 103348 238252
rect 104972 238084 105028 390124
rect 106652 238196 106708 393372
rect 106652 238130 106708 238140
rect 110012 384356 110068 384366
rect 104972 238018 105028 238028
rect 110012 237860 110068 384300
rect 111692 284452 111748 402556
rect 120092 391860 120148 391870
rect 116732 389284 116788 389294
rect 111692 284386 111748 284396
rect 113372 321748 113428 321758
rect 113372 278628 113428 321692
rect 113372 278562 113428 278572
rect 115052 320068 115108 320078
rect 115052 261156 115108 320012
rect 115052 261090 115108 261100
rect 116732 239764 116788 389228
rect 116732 239698 116788 239708
rect 120092 237972 120148 391804
rect 126812 388276 126868 388286
rect 126812 240772 126868 388220
rect 138572 386372 138628 386382
rect 138572 361396 138628 386316
rect 138572 361330 138628 361340
rect 143388 287924 143444 595560
rect 165452 590548 165508 590558
rect 148652 570388 148708 570398
rect 148652 289044 148708 570332
rect 165452 399252 165508 590492
rect 165676 590212 165732 595560
rect 165676 590146 165732 590156
rect 168812 590212 168868 590222
rect 165452 399186 165508 399196
rect 168812 397796 168868 590156
rect 187740 590212 187796 595560
rect 209580 595560 209832 595672
rect 231644 595560 231896 595672
rect 253708 595560 253960 595672
rect 275772 595560 276024 595672
rect 297836 595560 298088 595672
rect 319900 595560 320152 595672
rect 341964 595560 342216 595672
rect 364028 595560 364280 595672
rect 386092 595560 386344 595672
rect 408184 595560 408408 597000
rect 430248 595672 430472 597000
rect 430220 595560 430472 595672
rect 452312 595672 452536 597000
rect 474376 595672 474600 597000
rect 452312 595560 452564 595672
rect 190540 591220 190596 591230
rect 190316 590772 190372 590782
rect 187740 590146 187796 590156
rect 188972 590212 189028 590222
rect 182252 587188 182308 587198
rect 177212 573076 177268 573086
rect 175532 446068 175588 446078
rect 175532 400708 175588 446012
rect 175532 400642 175588 400652
rect 168812 397730 168868 397740
rect 177212 390740 177268 573020
rect 181356 410788 181412 410798
rect 181356 408100 181412 410732
rect 182252 409668 182308 587132
rect 182252 409602 182308 409612
rect 188972 409556 189028 590156
rect 188972 409490 189028 409500
rect 190316 409108 190372 590716
rect 190316 409042 190372 409052
rect 190428 572068 190484 572078
rect 181356 408034 181412 408044
rect 190428 393988 190484 572012
rect 190540 408324 190596 591164
rect 190540 408258 190596 408268
rect 190652 590996 190708 591006
rect 190652 407988 190708 590940
rect 209580 590436 209636 595560
rect 209580 590370 209636 590380
rect 231644 572068 231700 595560
rect 253708 591332 253764 595560
rect 253708 591266 253764 591276
rect 275772 591220 275828 595560
rect 275772 591154 275828 591164
rect 297836 591108 297892 595560
rect 297836 591042 297892 591052
rect 319900 590996 319956 595560
rect 319900 590930 319956 590940
rect 341964 590884 342020 595560
rect 341964 590818 342020 590828
rect 364028 590772 364084 595560
rect 364028 590706 364084 590716
rect 386092 590660 386148 595560
rect 408268 591332 408324 595560
rect 408268 591266 408324 591276
rect 386092 590594 386148 590604
rect 430220 590548 430276 595560
rect 430220 590482 430276 590492
rect 452508 590548 452564 595560
rect 474348 595560 474600 595672
rect 496440 595672 496664 597000
rect 518504 595672 518728 597000
rect 496440 595560 496692 595672
rect 474348 591332 474404 595560
rect 474348 591266 474404 591276
rect 496636 590660 496692 595560
rect 496636 590594 496692 590604
rect 518476 595560 518728 595672
rect 540568 595672 540792 597000
rect 562632 595672 562856 597000
rect 584696 595672 584920 597000
rect 540568 595560 540820 595672
rect 452508 590482 452564 590492
rect 231644 572002 231700 572012
rect 518476 570388 518532 595560
rect 540764 590772 540820 595560
rect 562604 595560 562856 595672
rect 584668 595560 584920 595672
rect 560252 591332 560308 591342
rect 540764 590706 540820 590716
rect 549836 590772 549892 590782
rect 518476 570322 518532 570332
rect 549388 550452 549444 550462
rect 548492 410564 548548 410574
rect 190652 407922 190708 407932
rect 195132 406644 195188 410088
rect 195132 406578 195188 406588
rect 197372 408324 197428 408334
rect 190428 393922 190484 393932
rect 177212 390674 177268 390684
rect 196588 346948 196644 346958
rect 181356 313348 181412 313358
rect 148652 288978 148708 288988
rect 163772 297444 163828 297454
rect 163772 290612 163828 297388
rect 143388 287858 143444 287868
rect 163772 285908 163828 290556
rect 172844 289940 172900 289950
rect 163772 285852 164360 285908
rect 172844 285880 172900 289884
rect 181356 285880 181412 313292
rect 192332 289044 192388 289054
rect 192332 253652 192388 288988
rect 196588 285348 196644 346892
rect 196700 343588 196756 343598
rect 196700 286468 196756 343532
rect 197372 302428 197428 408268
rect 198268 406644 198324 406654
rect 198268 349468 198324 406588
rect 198268 349412 198548 349468
rect 198380 336868 198436 336878
rect 197372 302372 197540 302428
rect 196700 286402 196756 286412
rect 197484 285684 197540 302372
rect 197484 285618 197540 285628
rect 196588 285282 196644 285292
rect 197372 284788 197428 284798
rect 192332 253586 192388 253596
rect 196476 257124 196532 257134
rect 196476 245924 196532 257068
rect 197372 257124 197428 284732
rect 198380 284788 198436 336812
rect 198380 284722 198436 284732
rect 198492 329476 198548 349412
rect 199164 339220 199220 339230
rect 197372 257058 197428 257068
rect 196476 245858 196532 245868
rect 198492 243684 198548 329420
rect 199052 333508 199108 333518
rect 199052 249620 199108 333452
rect 199164 320068 199220 339164
rect 200508 333508 200564 410088
rect 204092 391972 204148 391982
rect 200508 333442 200564 333452
rect 202412 368788 202468 368798
rect 199164 320002 199220 320012
rect 200732 331604 200788 331614
rect 199052 249554 199108 249564
rect 198492 243572 199108 243628
rect 126812 240706 126868 240716
rect 120092 237906 120148 237916
rect 110012 237794 110068 237804
rect 100380 237570 100436 237580
rect 72940 234994 72996 235004
rect 41020 232708 41076 232718
rect 40236 229460 40292 229470
rect 40124 217700 40180 217710
rect 40124 4340 40180 217644
rect 40124 4274 40180 4284
rect 38556 4162 38612 4172
rect 39900 4228 39956 4238
rect 39900 480 39956 4172
rect 40236 4228 40292 229404
rect 40236 4162 40292 4172
rect 13244 392 13496 480
rect 15148 392 15400 480
rect 17052 392 17304 480
rect 18956 392 19208 480
rect 20860 392 21112 480
rect 22764 392 23016 480
rect 24668 392 24920 480
rect 26572 392 26824 480
rect 11368 -960 11592 392
rect 13272 -960 13496 392
rect 15176 -960 15400 392
rect 17080 -960 17304 392
rect 18984 -960 19208 392
rect 20888 -960 21112 392
rect 22792 -960 23016 392
rect 24696 -960 24920 392
rect 26600 -960 26824 392
rect 28504 -960 28728 480
rect 30380 392 30632 480
rect 32284 392 32536 480
rect 34188 392 34440 480
rect 30408 -960 30632 392
rect 32312 -960 32536 392
rect 34216 -960 34440 392
rect 36120 -960 36344 480
rect 37996 392 38248 480
rect 39900 392 40152 480
rect 38024 -960 38248 392
rect 39928 -960 40152 392
rect 41020 420 41076 232652
rect 41132 231028 41188 231038
rect 41132 4452 41188 230972
rect 199052 215908 199108 243572
rect 199052 215842 199108 215852
rect 154924 214228 154980 214238
rect 154924 209944 154980 214172
rect 200732 214228 200788 331548
rect 202412 289940 202468 368732
rect 202412 289874 202468 289884
rect 204092 238532 204148 391916
rect 205772 388500 205828 388510
rect 205772 239988 205828 388444
rect 205884 336868 205940 410088
rect 210812 388724 210868 388734
rect 205884 336802 205940 336812
rect 207452 384244 207508 384254
rect 205772 239922 205828 239932
rect 204092 238466 204148 238476
rect 207452 234388 207508 384188
rect 210812 240100 210868 388668
rect 211260 339220 211316 410088
rect 215852 388836 215908 388846
rect 211260 339154 211316 339164
rect 212492 386260 212548 386270
rect 212492 319060 212548 386204
rect 212492 318994 212548 319004
rect 214172 370804 214228 370814
rect 214172 313348 214228 370748
rect 214172 313282 214228 313292
rect 215852 240436 215908 388780
rect 216636 384748 216692 410088
rect 222040 410060 222628 410116
rect 227416 410060 227668 410116
rect 222572 403284 222628 410060
rect 219212 389172 219268 389182
rect 215964 384692 216692 384748
rect 217532 388948 217588 388958
rect 215964 383236 216020 384692
rect 215964 343588 216020 383180
rect 215964 343522 216020 343532
rect 215964 311668 216020 311678
rect 215964 290164 216020 311612
rect 215964 290098 216020 290108
rect 215852 240370 215908 240380
rect 217532 240212 217588 388892
rect 217532 240146 217588 240156
rect 217756 388612 217812 388622
rect 210812 240034 210868 240044
rect 217756 239876 217812 388556
rect 219212 240324 219268 389116
rect 222572 346948 222628 403228
rect 227612 406644 227668 410060
rect 223244 368564 223300 368574
rect 222572 346882 222628 346892
rect 223132 361844 223188 361854
rect 219212 240258 219268 240268
rect 219996 343924 220052 343934
rect 217756 239810 217812 239820
rect 219996 237748 220052 343868
rect 223020 339444 223076 339454
rect 223020 241556 223076 339388
rect 223132 249508 223188 361788
rect 223244 251188 223300 368508
rect 226716 367444 226772 367454
rect 225036 365204 225092 365214
rect 223244 251122 223300 251132
rect 223356 364084 223412 364094
rect 223132 249442 223188 249452
rect 223020 241490 223076 241500
rect 223356 241220 223412 364028
rect 224924 341684 224980 341694
rect 224924 248164 224980 341628
rect 224924 248098 224980 248108
rect 225036 247828 225092 365148
rect 226492 359604 226548 359614
rect 226380 357364 226436 357374
rect 225036 247762 225092 247772
rect 226268 345044 226324 345054
rect 226268 244468 226324 344988
rect 226380 247940 226436 357308
rect 226492 251300 226548 359548
rect 226492 251234 226548 251244
rect 226604 355124 226660 355134
rect 226380 247874 226436 247884
rect 226268 244402 226324 244412
rect 226604 241332 226660 355068
rect 226716 242788 226772 367388
rect 227612 323428 227668 406588
rect 227948 407988 228004 407998
rect 227836 350644 227892 350654
rect 227612 323362 227668 323372
rect 227724 326116 227780 326126
rect 227500 306964 227556 306974
rect 227500 246372 227556 306908
rect 227612 297556 227668 297566
rect 227612 251748 227668 297500
rect 227612 251682 227668 251692
rect 227500 246306 227556 246316
rect 226716 242722 226772 242732
rect 226604 241266 226660 241276
rect 223356 241154 223412 241164
rect 227724 239988 227780 326060
rect 227836 251412 227892 350588
rect 227948 304052 228004 407932
rect 230188 407540 230244 407550
rect 230188 406532 230244 407484
rect 230188 406466 230244 406476
rect 232764 406756 232820 410088
rect 228508 404516 228564 404526
rect 228508 404068 228564 404460
rect 228508 404002 228564 404012
rect 229516 404516 229572 404526
rect 229404 393540 229460 393550
rect 229292 392084 229348 392094
rect 228396 362964 228452 362974
rect 228284 358484 228340 358494
rect 228172 352884 228228 352894
rect 227948 303268 228004 303996
rect 227948 303202 228004 303212
rect 228060 349524 228116 349534
rect 227836 251346 227892 251356
rect 228060 241444 228116 349468
rect 228172 243012 228228 352828
rect 228172 242946 228228 242956
rect 228284 242900 228340 358428
rect 228396 246148 228452 362908
rect 228396 246082 228452 246092
rect 228284 242834 228340 242844
rect 228060 241378 228116 241388
rect 227724 239922 227780 239932
rect 219996 237682 220052 237692
rect 229292 235060 229348 392028
rect 229404 236628 229460 393484
rect 229516 301588 229572 404460
rect 231196 404404 231252 404414
rect 230076 354004 230132 354014
rect 229852 348404 229908 348414
rect 229740 340564 229796 340574
rect 229516 300804 229572 301532
rect 229516 300738 229572 300748
rect 229628 304052 229684 304062
rect 229404 236562 229460 236572
rect 229292 234994 229348 235004
rect 207452 234322 207508 234332
rect 229628 216244 229684 303996
rect 229740 246260 229796 340508
rect 229852 249844 229908 348348
rect 229852 249778 229908 249788
rect 229964 339556 230020 339566
rect 229740 246194 229796 246204
rect 229964 239764 230020 339500
rect 230076 239876 230132 353948
rect 231196 322532 231252 404348
rect 232764 402612 232820 406700
rect 237692 407988 237748 407998
rect 237692 404628 237748 407932
rect 238140 407764 238196 410088
rect 238140 407698 238196 407708
rect 243516 407652 243572 410088
rect 243516 406644 243572 407596
rect 248892 406868 248948 410088
rect 252588 409444 252644 409454
rect 248892 406802 248948 406812
rect 251692 409220 251748 409230
rect 243516 406588 243796 406644
rect 237692 404562 237748 404572
rect 232764 402546 232820 402556
rect 231644 400820 231700 400830
rect 231532 347284 231588 347294
rect 231420 337204 231476 337214
rect 231196 322466 231252 322476
rect 231308 336084 231364 336094
rect 230972 300804 231028 300814
rect 230972 250068 231028 300748
rect 231084 276388 231140 276398
rect 231084 254996 231140 276332
rect 231084 254930 231140 254940
rect 231308 251524 231364 336028
rect 231308 251458 231364 251468
rect 230972 250002 231028 250012
rect 231420 244580 231476 337148
rect 231420 244514 231476 244524
rect 230188 243236 230244 243246
rect 230188 242564 230244 243180
rect 231532 243124 231588 347228
rect 231644 243236 231700 400764
rect 233324 397460 233380 397470
rect 231644 243170 231700 243180
rect 231756 394100 231812 394110
rect 231532 243058 231588 243068
rect 230188 242498 230244 242508
rect 230076 239810 230132 239820
rect 229964 239698 230020 239708
rect 231756 216468 231812 394044
rect 233212 369684 233268 369694
rect 233212 368788 233268 369628
rect 233212 368722 233268 368732
rect 233212 366324 233268 366334
rect 232652 360724 232708 360734
rect 232652 339556 232708 360668
rect 232652 339490 232708 339500
rect 232764 342804 232820 342814
rect 232764 326116 232820 342748
rect 233212 331828 233268 366268
rect 233212 331762 233268 331772
rect 232764 326050 232820 326060
rect 231868 322532 231924 322542
rect 231868 246932 231924 322476
rect 233212 309204 233268 309214
rect 233100 308084 233156 308094
rect 233100 257348 233156 308028
rect 233100 257282 233156 257292
rect 233212 256116 233268 309148
rect 233324 281204 233380 397404
rect 243740 396508 243796 406588
rect 249900 405748 249956 405758
rect 247212 404068 247268 404078
rect 246316 399140 246372 399150
rect 243740 396452 243908 396508
rect 236012 392308 236068 392318
rect 235004 387380 235060 387390
rect 234556 386148 234612 386158
rect 234332 386036 234388 386046
rect 233324 281138 233380 281148
rect 233436 384580 233492 384590
rect 233212 256050 233268 256060
rect 233324 264404 233380 264414
rect 233324 254548 233380 264348
rect 233324 254482 233380 254492
rect 231868 246866 231924 246876
rect 231756 216402 231812 216412
rect 229628 216178 229684 216188
rect 200732 214162 200788 214172
rect 233436 213108 233492 384524
rect 234220 281428 234276 281438
rect 234220 254884 234276 281372
rect 234220 254818 234276 254828
rect 234332 235172 234388 385980
rect 234444 331828 234500 331838
rect 234444 239652 234500 331772
rect 234444 239586 234500 239596
rect 234556 236852 234612 386092
rect 234892 351764 234948 351774
rect 234780 334964 234836 334974
rect 234668 284004 234724 284014
rect 234668 256452 234724 283948
rect 234668 256386 234724 256396
rect 234780 251636 234836 334908
rect 234780 251570 234836 251580
rect 234892 248052 234948 351708
rect 234892 247986 234948 247996
rect 234556 236786 234612 236796
rect 234332 235106 234388 235116
rect 235004 216132 235060 387324
rect 235004 216066 235060 216076
rect 235116 385812 235172 385822
rect 235116 213332 235172 385756
rect 235676 385700 235732 385710
rect 235676 384748 235732 385644
rect 235788 385588 235844 385598
rect 235844 385532 235956 385588
rect 235788 385522 235844 385532
rect 235676 384692 235844 384748
rect 235116 213266 235172 213276
rect 235676 384468 235732 384478
rect 233436 213042 233492 213052
rect 235676 212772 235732 384412
rect 235788 212884 235844 384692
rect 235788 212818 235844 212828
rect 235676 212706 235732 212716
rect 235900 212660 235956 385532
rect 236012 375508 236068 392252
rect 242732 390404 242788 390414
rect 240940 390292 240996 390302
rect 240044 389844 240100 389854
rect 238252 388164 238308 388174
rect 237356 387044 237412 387054
rect 237356 385896 237412 386988
rect 238252 385896 238308 388108
rect 239148 386484 239204 386494
rect 239148 385896 239204 386428
rect 240044 385896 240100 389788
rect 240940 385896 240996 390236
rect 241836 386596 241892 386606
rect 241836 385896 241892 386540
rect 242732 385896 242788 390348
rect 243628 387156 243684 387166
rect 243628 385896 243684 387100
rect 243852 385812 243908 396452
rect 245420 390516 245476 390526
rect 245420 385896 245476 390460
rect 246316 385896 246372 399084
rect 247212 385896 247268 404012
rect 248108 402612 248164 402622
rect 248108 385896 248164 402556
rect 249004 397572 249060 397582
rect 249004 385896 249060 397516
rect 249900 385896 249956 405692
rect 250796 397684 250852 397694
rect 250796 385896 250852 397628
rect 251692 385896 251748 409164
rect 252588 385896 252644 409388
rect 253484 409108 253540 409118
rect 253484 385896 253540 409052
rect 254268 407428 254324 410088
rect 259672 410060 260372 410116
rect 254268 407362 254324 407372
rect 254380 409332 254436 409342
rect 254380 385896 254436 409276
rect 260316 408268 260372 410060
rect 260316 408212 260484 408268
rect 260428 406868 260484 408212
rect 265020 407540 265076 410088
rect 270396 407988 270452 410088
rect 275548 410060 275800 410116
rect 280588 410060 281176 410116
rect 286300 410088 286552 410116
rect 308056 410088 308868 410116
rect 286300 410060 286580 410088
rect 270396 407922 270452 407932
rect 273756 409108 273812 409118
rect 273756 407652 273812 409052
rect 275548 408268 275604 410060
rect 273756 407586 273812 407596
rect 275436 408212 275604 408268
rect 280588 409556 280644 410060
rect 265020 407474 265076 407484
rect 259756 404180 259812 404190
rect 257068 399252 257124 399262
rect 256172 397796 256228 397806
rect 255276 393988 255332 393998
rect 255276 385896 255332 393932
rect 256172 385896 256228 397740
rect 257068 385896 257124 399196
rect 258860 390740 258916 390750
rect 257964 390628 258020 390638
rect 257964 385896 258020 390572
rect 258860 385896 258916 390684
rect 259756 385896 259812 404124
rect 260428 394100 260484 406812
rect 275436 404516 275492 408212
rect 275436 404450 275492 404460
rect 262444 403732 262500 403742
rect 260428 394034 260484 394044
rect 260652 402724 260708 402734
rect 260652 385896 260708 402668
rect 261548 400708 261604 400718
rect 261548 385896 261604 400652
rect 262444 385896 262500 403676
rect 270508 389956 270564 389966
rect 268716 386820 268772 386830
rect 266924 386708 266980 386718
rect 263340 386372 263396 386382
rect 263340 385896 263396 386316
rect 264236 386260 264292 386270
rect 264236 385896 264292 386204
rect 266924 385896 266980 386652
rect 268716 385896 268772 386764
rect 270508 385896 270564 389900
rect 272300 389956 272356 389966
rect 272300 385896 272356 389900
rect 277676 388388 277732 388398
rect 274092 387380 274148 387390
rect 274092 385896 274148 387324
rect 277676 385896 277732 388332
rect 278572 386820 278628 386830
rect 278572 385896 278628 386764
rect 280364 386372 280420 386382
rect 279468 386260 279524 386270
rect 279468 385896 279524 386204
rect 280364 385896 280420 386316
rect 280588 385924 280644 409500
rect 286300 406980 286356 410060
rect 286524 409780 286580 410060
rect 286524 409714 286580 409724
rect 290668 409892 290724 409902
rect 286300 406914 286356 406924
rect 290668 392532 290724 409836
rect 291900 409892 291956 410088
rect 291900 409826 291956 409836
rect 295708 409668 295764 409678
rect 290668 392466 290724 392476
rect 292012 393204 292068 393214
rect 282156 388164 282212 388174
rect 282156 385896 282212 388108
rect 283948 386708 284004 386718
rect 283948 385896 284004 386652
rect 292012 385896 292068 393148
rect 295708 392420 295764 409612
rect 297276 409668 297332 410088
rect 297276 409602 297332 409612
rect 302652 408884 302708 410088
rect 308028 410060 308868 410088
rect 308028 409332 308084 410060
rect 308028 409266 308084 409276
rect 302652 406980 302708 408828
rect 302652 406914 302708 406924
rect 295708 392354 295764 392364
rect 304556 393540 304612 393550
rect 301868 389284 301924 389294
rect 300972 389172 301028 389182
rect 300076 388948 300132 388958
rect 299180 388836 299236 388846
rect 296492 388724 296548 388734
rect 295596 388276 295652 388286
rect 295596 385896 295652 388220
rect 296492 385896 296548 388668
rect 298284 388500 298340 388510
rect 297388 388164 297444 388174
rect 297388 385896 297444 388108
rect 298284 385896 298340 388444
rect 299180 385896 299236 388780
rect 300076 385896 300132 388892
rect 300972 385896 301028 389116
rect 301868 385896 301924 389228
rect 302764 386148 302820 386158
rect 302764 385896 302820 386092
rect 302988 386036 303044 386046
rect 302988 385924 303044 385980
rect 302988 385868 303688 385924
rect 304556 385896 304612 393484
rect 305452 392084 305508 392094
rect 305452 385896 305508 392028
rect 307244 391748 307300 391758
rect 306348 386932 306404 386942
rect 306348 385896 306404 386876
rect 307244 385896 307300 391692
rect 308140 388612 308196 388622
rect 308140 385896 308196 388556
rect 308812 386036 308868 410060
rect 313292 410060 313432 410116
rect 318332 410060 318808 410116
rect 313292 408100 313348 410060
rect 310828 391860 310884 391870
rect 308812 385970 308868 385980
rect 309932 390068 309988 390078
rect 309932 385896 309988 390012
rect 310828 385896 310884 391804
rect 312620 391636 312676 391646
rect 311724 390180 311780 390190
rect 311724 385896 311780 390124
rect 312620 385896 312676 391580
rect 313292 386036 313348 408044
rect 318332 407876 318388 410060
rect 317996 397796 318052 397806
rect 316204 393428 316260 393438
rect 315308 393316 315364 393326
rect 314412 391972 314468 391982
rect 313292 385970 313348 385980
rect 313516 391524 313572 391534
rect 313516 385896 313572 391468
rect 314412 385896 314468 391916
rect 315308 385896 315364 393260
rect 316204 385896 316260 393372
rect 317100 388948 317156 388958
rect 317100 385896 317156 388892
rect 317996 385896 318052 397740
rect 318332 386148 318388 407820
rect 322476 402276 322532 402286
rect 319788 400708 319844 400718
rect 318332 386082 318388 386092
rect 318892 392420 318948 392430
rect 318892 385896 318948 392364
rect 319788 385896 319844 400652
rect 321580 395780 321636 395790
rect 320684 392196 320740 392206
rect 320684 385896 320740 392140
rect 321580 385896 321636 395724
rect 322476 385896 322532 402220
rect 323372 395668 323428 395678
rect 322588 393204 322644 393214
rect 322588 392308 322644 393148
rect 322588 392242 322644 392252
rect 323372 385896 323428 395612
rect 324156 393204 324212 410088
rect 328748 409332 328804 409342
rect 324156 393138 324212 393148
rect 324268 406308 324324 406318
rect 324268 385896 324324 406252
rect 327852 404740 327908 404750
rect 326732 401156 326788 401166
rect 326060 393092 326116 393102
rect 325164 389060 325220 389070
rect 325164 385896 325220 389004
rect 326060 385896 326116 393036
rect 326732 388948 326788 401100
rect 326732 388882 326788 388892
rect 326956 389284 327012 389294
rect 326956 385896 327012 389228
rect 327852 385896 327908 404684
rect 328748 385896 328804 409276
rect 329532 404404 329588 410088
rect 333452 409556 333508 409566
rect 329532 404338 329588 404348
rect 332332 409444 332388 409454
rect 331436 401044 331492 401054
rect 330876 395892 330932 395902
rect 329644 392308 329700 392318
rect 329644 385896 329700 392252
rect 330540 389732 330596 389742
rect 330540 385896 330596 389676
rect 330876 389060 330932 395836
rect 330876 388994 330932 389004
rect 331436 385896 331492 400988
rect 332332 385896 332388 409388
rect 333228 390852 333284 390862
rect 333228 385896 333284 390796
rect 333452 389732 333508 409500
rect 334908 400932 334964 410088
rect 334908 400866 334964 400876
rect 338604 404628 338660 404638
rect 336812 399700 336868 399710
rect 335916 399252 335972 399262
rect 333452 389666 333508 389676
rect 335020 394772 335076 394782
rect 334124 388948 334180 388958
rect 334124 385896 334180 388892
rect 335020 385896 335076 394716
rect 335916 385896 335972 399196
rect 336812 385896 336868 399644
rect 337708 393988 337764 393998
rect 337708 385896 337764 393932
rect 338604 385896 338660 404572
rect 340284 400820 340340 410088
rect 345660 407652 345716 410088
rect 351036 407764 351092 410088
rect 351036 407698 351092 407708
rect 355628 409668 355684 409678
rect 345660 407586 345716 407596
rect 351148 406196 351204 406206
rect 349356 404516 349412 404526
rect 340284 400754 340340 400764
rect 340396 403172 340452 403182
rect 339500 394100 339556 394110
rect 339500 385896 339556 394044
rect 340396 385896 340452 403116
rect 348460 402724 348516 402734
rect 342188 400932 342244 400942
rect 341292 394212 341348 394222
rect 341292 385896 341348 394156
rect 342188 385896 342244 400876
rect 345772 399588 345828 399598
rect 343980 398132 344036 398142
rect 343084 394324 343140 394334
rect 343084 385896 343140 394268
rect 343980 385896 344036 398076
rect 344876 394548 344932 394558
rect 344876 385896 344932 394492
rect 345772 385896 345828 399532
rect 346668 394436 346724 394446
rect 346668 385896 346724 394380
rect 347564 389172 347620 389182
rect 347564 385896 347620 389116
rect 348460 385896 348516 402668
rect 349356 385896 349412 404460
rect 350252 396004 350308 396014
rect 350252 385896 350308 395948
rect 351148 385896 351204 406140
rect 353836 404180 353892 404190
rect 352940 403060 352996 403070
rect 352044 396116 352100 396126
rect 352044 385896 352100 396060
rect 352940 385896 352996 403004
rect 353836 385896 353892 404124
rect 354732 392980 354788 392990
rect 354732 385896 354788 392924
rect 355628 385896 355684 409612
rect 356412 407876 356468 410088
rect 356412 407810 356468 407820
rect 360332 407540 360388 407550
rect 359212 405860 359268 405870
rect 358316 392868 358372 392878
rect 356524 392756 356580 392766
rect 356524 385896 356580 392700
rect 357420 390628 357476 390638
rect 357420 385896 357476 390572
rect 358316 385896 358372 392812
rect 359212 385896 359268 405804
rect 360108 392644 360164 392654
rect 360108 385896 360164 392588
rect 360332 392308 360388 407484
rect 361788 404852 361844 410088
rect 361788 404786 361844 404796
rect 362796 409780 362852 409790
rect 360332 392242 360388 392252
rect 361004 394660 361060 394670
rect 361004 385896 361060 394604
rect 361900 392532 361956 392542
rect 361900 385896 361956 392476
rect 362796 385896 362852 409724
rect 365372 407988 365428 407998
rect 363692 400820 363748 400830
rect 363692 385896 363748 400764
rect 365372 392420 365428 407932
rect 367164 401492 367220 410088
rect 367164 401426 367220 401436
rect 368732 409892 368788 409902
rect 367276 399476 367332 399486
rect 365372 392354 365428 392364
rect 365484 398020 365540 398030
rect 364588 392308 364644 392318
rect 364588 385896 364644 392252
rect 365484 385896 365540 397964
rect 366380 389732 366436 389742
rect 366380 385896 366436 389676
rect 367276 385896 367332 399420
rect 368732 389732 368788 409836
rect 368732 389666 368788 389676
rect 369068 404404 369124 404414
rect 368172 389060 368228 389070
rect 368172 385896 368228 389004
rect 369068 385896 369124 404348
rect 370860 402948 370916 402958
rect 369964 395556 370020 395566
rect 369964 385896 370020 395500
rect 370860 385896 370916 402892
rect 372540 401156 372596 410088
rect 377916 407988 377972 410088
rect 377916 407922 377972 407932
rect 375676 407876 375732 407886
rect 375564 407764 375620 407774
rect 372540 401090 372596 401100
rect 374444 406084 374500 406094
rect 372652 392420 372708 392430
rect 371308 390964 371364 390974
rect 371308 389172 371364 390908
rect 371308 389106 371364 389116
rect 371756 389396 371812 389406
rect 371756 385896 371812 389340
rect 372652 385896 372708 392364
rect 373548 389172 373604 389182
rect 373548 385896 373604 389116
rect 374444 385896 374500 406028
rect 375340 388164 375396 388174
rect 375340 385896 375396 388108
rect 280588 385858 280644 385868
rect 243852 385746 243908 385756
rect 244524 385812 244580 385822
rect 244524 385746 244580 385756
rect 274988 385700 275044 385710
rect 274988 385634 275044 385644
rect 284844 385700 284900 385710
rect 284844 385634 284900 385644
rect 276780 385588 276836 385598
rect 276780 385522 276836 385532
rect 286636 385588 286692 385598
rect 286636 385522 286692 385532
rect 265132 385476 265188 385486
rect 265132 385410 265188 385420
rect 267820 385476 267876 385486
rect 267820 385410 267876 385420
rect 273196 385476 273252 385486
rect 273196 385410 273252 385420
rect 285740 385476 285796 385486
rect 285740 385410 285796 385420
rect 236124 385364 236180 385374
rect 266028 385364 266084 385374
rect 236180 385308 236488 385364
rect 236124 385298 236180 385308
rect 266028 385298 266084 385308
rect 269612 385364 269668 385374
rect 269612 385298 269668 385308
rect 271404 385364 271460 385374
rect 271404 385298 271460 385308
rect 275884 385364 275940 385374
rect 275884 385298 275940 385308
rect 281260 385364 281316 385374
rect 281260 385298 281316 385308
rect 283052 385364 283108 385374
rect 283052 385298 283108 385308
rect 287532 385364 287588 385374
rect 287532 385298 287588 385308
rect 288428 385364 288484 385374
rect 288428 385298 288484 385308
rect 289324 385364 289380 385374
rect 289324 385298 289380 385308
rect 290220 385364 290276 385374
rect 290220 385298 290276 385308
rect 291116 385364 291172 385374
rect 291116 385298 291172 385308
rect 292908 385364 292964 385374
rect 292908 385298 292964 385308
rect 293804 385364 293860 385374
rect 293804 385298 293860 385308
rect 294700 385364 294756 385374
rect 294700 385298 294756 385308
rect 309036 385364 309092 385374
rect 309036 385298 309092 385308
rect 236012 375442 236068 375452
rect 236012 356020 236068 356030
rect 236012 249732 236068 355964
rect 236012 249666 236068 249676
rect 236124 345940 236180 345950
rect 236124 248276 236180 345884
rect 236236 337988 236292 337998
rect 236236 249956 236292 337932
rect 242732 253652 242788 256088
rect 242732 253586 242788 253596
rect 243628 252084 243684 256088
rect 236236 249890 236292 249900
rect 242956 252028 243684 252084
rect 236124 248210 236180 248220
rect 242956 222740 243012 252028
rect 244524 224420 244580 256088
rect 244524 224354 244580 224364
rect 242956 222674 243012 222684
rect 235900 212594 235956 212604
rect 245420 210868 245476 256088
rect 246316 232820 246372 256088
rect 246316 232754 246372 232764
rect 247212 227780 247268 256088
rect 247212 227714 247268 227724
rect 248108 217700 248164 256088
rect 249004 231140 249060 256088
rect 249004 231074 249060 231084
rect 248108 217634 248164 217644
rect 249900 216020 249956 256088
rect 250796 229460 250852 256088
rect 251692 255388 251748 256088
rect 251692 255332 251972 255388
rect 251916 253652 251972 255332
rect 251916 253586 251972 253596
rect 252588 253652 252644 256088
rect 252588 253586 252644 253596
rect 253484 249396 253540 256088
rect 253484 249330 253540 249340
rect 254380 246484 254436 256088
rect 255276 246596 255332 256088
rect 256172 250180 256228 256088
rect 256172 250114 256228 250124
rect 255276 246530 255332 246540
rect 254380 246418 254436 246428
rect 257068 246036 257124 256088
rect 257068 245970 257124 245980
rect 257964 243348 258020 256088
rect 258860 253652 258916 256088
rect 258860 253586 258916 253596
rect 259756 253652 259812 256088
rect 259756 253586 259812 253596
rect 260652 253652 260708 256088
rect 260652 253586 260708 253596
rect 261548 252980 261604 256088
rect 261548 252914 261604 252924
rect 262444 252868 262500 256088
rect 263340 253092 263396 256088
rect 264236 253316 264292 256088
rect 264236 253250 264292 253260
rect 265132 253204 265188 256088
rect 266028 253540 266084 256088
rect 266028 253474 266084 253484
rect 265132 253138 265188 253148
rect 263340 253026 263396 253036
rect 262444 252802 262500 252812
rect 266924 252084 266980 256088
rect 267820 252308 267876 256088
rect 267820 252242 267876 252252
rect 268716 252196 268772 256088
rect 268716 252130 268772 252140
rect 266924 252018 266980 252028
rect 257964 243282 258020 243292
rect 250796 229394 250852 229404
rect 249900 215954 249956 215964
rect 269388 216468 269444 216478
rect 245420 210802 245476 210812
rect 269276 213332 269332 213342
rect 269276 79268 269332 213276
rect 269388 88228 269444 216412
rect 269500 211204 269556 211214
rect 269500 210756 269556 211148
rect 269500 210690 269556 210700
rect 269500 209748 269556 209758
rect 269500 204708 269556 209692
rect 269500 204642 269556 204652
rect 269388 88162 269444 88172
rect 269500 142884 269556 142894
rect 269276 79202 269332 79212
rect 269500 50372 269556 142828
rect 269500 50306 269556 50316
rect 91308 49588 91364 49598
rect 47852 48692 47908 48702
rect 47516 15988 47572 15998
rect 41132 4386 41188 4396
rect 45612 4900 45668 4910
rect 41692 480 41860 532
rect 45612 480 45668 4844
rect 47516 480 47572 15932
rect 47852 5908 47908 48636
rect 87500 47908 87556 47918
rect 68460 41188 68516 41198
rect 57148 37828 57204 37838
rect 47852 5842 47908 5852
rect 55132 17668 55188 17678
rect 49420 4452 49476 4462
rect 49420 480 49476 4396
rect 53228 4340 53284 4350
rect 53228 480 53284 4284
rect 55132 480 55188 17612
rect 57148 480 57204 37772
rect 62748 34468 62804 34478
rect 60844 19348 60900 19358
rect 58940 4564 58996 4574
rect 58940 480 58996 4508
rect 60844 480 60900 19292
rect 62748 480 62804 34412
rect 66780 4676 66836 4686
rect 64652 4452 64708 4462
rect 64652 480 64708 4396
rect 66780 480 66836 4620
rect 41692 476 42056 480
rect 41692 420 41748 476
rect 41020 364 41748 420
rect 41804 392 42056 476
rect 41832 -960 42056 392
rect 43736 -960 43960 480
rect 45612 392 45864 480
rect 47516 392 47768 480
rect 49420 392 49672 480
rect 45640 -960 45864 392
rect 47544 -960 47768 392
rect 49448 -960 49672 392
rect 51352 -960 51576 480
rect 53228 392 53480 480
rect 55132 392 55384 480
rect 53256 -960 53480 392
rect 55160 -960 55384 392
rect 57064 -960 57288 480
rect 58940 392 59192 480
rect 60844 392 61096 480
rect 62748 392 63000 480
rect 64652 392 64904 480
rect 58968 -960 59192 392
rect 60872 -960 61096 392
rect 62776 -960 63000 392
rect 64680 -960 64904 392
rect 66584 392 66836 480
rect 68460 480 68516 41132
rect 76076 36148 76132 36158
rect 74172 34580 74228 34590
rect 72268 24388 72324 24398
rect 68908 9380 68964 9390
rect 68908 4676 68964 9324
rect 68908 4610 68964 4620
rect 70364 4228 70420 4238
rect 70364 480 70420 4172
rect 72268 480 72324 24332
rect 74172 480 74228 34524
rect 76076 480 76132 36092
rect 81788 34692 81844 34702
rect 79884 31108 79940 31118
rect 77980 14308 78036 14318
rect 77980 480 78036 14252
rect 79884 480 79940 31052
rect 81788 480 81844 34636
rect 83692 29428 83748 29438
rect 83692 480 83748 29372
rect 85820 4340 85876 4350
rect 85820 480 85876 4284
rect 68460 392 68712 480
rect 70364 392 70616 480
rect 72268 392 72520 480
rect 74172 392 74424 480
rect 76076 392 76328 480
rect 77980 392 78232 480
rect 79884 392 80136 480
rect 81788 392 82040 480
rect 83692 392 83944 480
rect 66584 -960 66808 392
rect 68488 -960 68712 392
rect 70392 -960 70616 392
rect 72296 -960 72520 392
rect 74200 -960 74424 392
rect 76104 -960 76328 392
rect 78008 -960 78232 392
rect 79912 -960 80136 392
rect 81816 -960 82040 392
rect 83720 -960 83944 392
rect 85624 392 85876 480
rect 87500 480 87556 47852
rect 89404 32900 89460 32910
rect 89404 480 89460 32844
rect 91308 480 91364 49532
rect 97356 48692 97412 50120
rect 180796 49924 180852 49934
rect 97356 48626 97412 48636
rect 167468 49812 167524 49822
rect 127484 48132 127540 48142
rect 93212 48020 93268 48030
rect 93212 480 93268 47964
rect 110348 44996 110404 45006
rect 104636 44884 104692 44894
rect 98924 44772 98980 44782
rect 97020 41300 97076 41310
rect 95116 19460 95172 19470
rect 95116 480 95172 19404
rect 97020 480 97076 41244
rect 98924 480 98980 44716
rect 102732 32788 102788 32798
rect 101052 5908 101108 5918
rect 101052 480 101108 5852
rect 87500 392 87752 480
rect 89404 392 89656 480
rect 91308 392 91560 480
rect 93212 392 93464 480
rect 95116 392 95368 480
rect 97020 392 97272 480
rect 98924 392 99176 480
rect 85624 -960 85848 392
rect 87528 -960 87752 392
rect 89432 -960 89656 392
rect 91336 -960 91560 392
rect 93240 -960 93464 392
rect 95144 -960 95368 392
rect 97048 -960 97272 392
rect 98952 -960 99176 392
rect 100856 392 101108 480
rect 102732 480 102788 32732
rect 104636 480 104692 44828
rect 108444 37940 108500 37950
rect 106764 7588 106820 7598
rect 106764 480 106820 7532
rect 102732 392 102984 480
rect 104636 392 104888 480
rect 100856 -960 101080 392
rect 102760 -960 102984 392
rect 104664 -960 104888 392
rect 106568 392 106820 480
rect 108444 480 108500 37884
rect 110348 480 110404 44940
rect 116060 41524 116116 41534
rect 112476 7700 112532 7710
rect 112476 480 112532 7644
rect 114380 4228 114436 4238
rect 114380 480 114436 4172
rect 108444 392 108696 480
rect 110348 392 110600 480
rect 106568 -960 106792 392
rect 108472 -960 108696 392
rect 110376 -960 110600 392
rect 112280 392 112532 480
rect 114184 392 114436 480
rect 116060 480 116116 41468
rect 119868 38052 119924 38062
rect 118188 7812 118244 7822
rect 118188 480 118244 7756
rect 116060 392 116312 480
rect 112280 -960 112504 392
rect 114184 -960 114408 392
rect 116088 -960 116312 392
rect 117992 392 118244 480
rect 119868 480 119924 37996
rect 121772 34916 121828 34926
rect 121772 480 121828 34860
rect 123676 17780 123732 17790
rect 123676 480 123732 17724
rect 125804 4900 125860 4910
rect 125804 480 125860 4844
rect 119868 392 120120 480
rect 121772 392 122024 480
rect 123676 392 123928 480
rect 117992 -960 118216 392
rect 119896 -960 120120 392
rect 121800 -960 122024 392
rect 123704 -960 123928 392
rect 125608 392 125860 480
rect 127484 480 127540 48076
rect 138908 45108 138964 45118
rect 133196 33012 133252 33022
rect 129388 16100 129444 16110
rect 129388 480 129444 16044
rect 131516 9268 131572 9278
rect 131516 480 131572 9212
rect 127484 392 127736 480
rect 129388 392 129640 480
rect 125608 -960 125832 392
rect 127512 -960 127736 392
rect 129416 -960 129640 392
rect 131320 392 131572 480
rect 133196 480 133252 32956
rect 135100 24500 135156 24510
rect 135100 480 135156 24444
rect 137228 4116 137284 4126
rect 137228 480 137284 4060
rect 133196 392 133448 480
rect 135100 392 135352 480
rect 131320 -960 131544 392
rect 133224 -960 133448 392
rect 135128 -960 135352 392
rect 137032 392 137284 480
rect 138908 480 138964 45052
rect 148428 44660 148484 44670
rect 142828 44548 142884 44558
rect 140812 14420 140868 14430
rect 140812 480 140868 14364
rect 142828 480 142884 44492
rect 144620 31332 144676 31342
rect 144620 480 144676 31276
rect 146524 26068 146580 26078
rect 146524 480 146580 26012
rect 148428 480 148484 44604
rect 156044 42980 156100 42990
rect 152236 31220 152292 31230
rect 150556 10948 150612 10958
rect 150556 480 150612 10892
rect 138908 392 139160 480
rect 140812 392 141064 480
rect 137032 -960 137256 392
rect 138936 -960 139160 392
rect 140840 -960 141064 392
rect 142744 -960 142968 480
rect 144620 392 144872 480
rect 146524 392 146776 480
rect 148428 392 148680 480
rect 144648 -960 144872 392
rect 146552 -960 146776 392
rect 148456 -960 148680 392
rect 150360 392 150612 480
rect 152236 480 152292 31164
rect 154364 4452 154420 4462
rect 154364 480 154420 4396
rect 152236 392 152488 480
rect 150360 -960 150584 392
rect 152264 -960 152488 392
rect 154168 392 154420 480
rect 156044 480 156100 42924
rect 159852 41412 159908 41422
rect 158172 6020 158228 6030
rect 158172 480 158228 5964
rect 156044 392 156296 480
rect 154168 -960 154392 392
rect 156072 -960 156296 392
rect 157976 392 158228 480
rect 159852 480 159908 41356
rect 161756 39508 161812 39518
rect 161756 480 161812 39452
rect 163660 12628 163716 12638
rect 163660 480 163716 12572
rect 165788 4564 165844 4574
rect 165788 480 165844 4508
rect 159852 392 160104 480
rect 161756 392 162008 480
rect 163660 392 163912 480
rect 157976 -960 158200 392
rect 159880 -960 160104 392
rect 161784 -960 162008 392
rect 163688 -960 163912 392
rect 165592 392 165844 480
rect 167468 480 167524 49756
rect 178892 48244 178948 48254
rect 175084 41636 175140 41646
rect 171388 38164 171444 38174
rect 169372 29540 169428 29550
rect 169372 480 169428 29484
rect 171388 480 171444 38108
rect 173180 26180 173236 26190
rect 173180 480 173236 26124
rect 175084 480 175140 41580
rect 177212 4676 177268 4686
rect 177212 480 177268 4620
rect 167468 392 167720 480
rect 169372 392 169624 480
rect 165592 -960 165816 392
rect 167496 -960 167720 392
rect 169400 -960 169624 392
rect 171304 -960 171528 480
rect 173180 392 173432 480
rect 175084 392 175336 480
rect 173208 -960 173432 392
rect 175112 -960 175336 392
rect 177016 392 177268 480
rect 178892 480 178948 48188
rect 180796 480 180852 49868
rect 212268 48580 212324 50120
rect 212268 48514 212324 48524
rect 197932 48356 197988 48366
rect 184604 46228 184660 46238
rect 182700 38276 182756 38286
rect 182700 480 182756 38220
rect 184604 480 184660 46172
rect 188412 42868 188468 42878
rect 186508 21028 186564 21038
rect 186508 480 186564 20972
rect 188412 480 188468 42812
rect 192220 38388 192276 38398
rect 190540 6132 190596 6142
rect 190540 480 190596 6076
rect 178892 392 179144 480
rect 180796 392 181048 480
rect 182700 392 182952 480
rect 184604 392 184856 480
rect 186508 392 186760 480
rect 188412 392 188664 480
rect 177016 -960 177240 392
rect 178920 -960 179144 392
rect 180824 -960 181048 392
rect 182728 -960 182952 392
rect 184632 -960 184856 392
rect 186536 -960 186760 392
rect 188440 -960 188664 392
rect 190344 392 190596 480
rect 192220 480 192276 38332
rect 194124 34804 194180 34814
rect 194124 480 194180 34748
rect 196028 24612 196084 24622
rect 196028 480 196084 24556
rect 197932 480 197988 48300
rect 207452 45220 207508 45230
rect 203644 41748 203700 41758
rect 201740 14532 201796 14542
rect 200060 4788 200116 4798
rect 200060 480 200116 4732
rect 192220 392 192472 480
rect 194124 392 194376 480
rect 196028 392 196280 480
rect 197932 392 198184 480
rect 190344 -960 190568 392
rect 192248 -960 192472 392
rect 194152 -960 194376 392
rect 196056 -960 196280 392
rect 197960 -960 198184 392
rect 199864 392 200116 480
rect 201740 480 201796 14476
rect 203644 480 203700 41692
rect 205772 5012 205828 5022
rect 205772 480 205828 4956
rect 201740 392 201992 480
rect 203644 392 203896 480
rect 199864 -960 200088 392
rect 201768 -960 201992 392
rect 203672 -960 203896 392
rect 205576 392 205828 480
rect 207452 480 207508 45164
rect 209356 36260 209412 36270
rect 209356 480 209412 36204
rect 211260 35028 211316 35038
rect 211260 480 211316 34972
rect 269612 6132 269668 256088
rect 269724 252084 269780 252094
rect 269724 26180 269780 252028
rect 269836 211428 269892 211438
rect 269836 207956 269892 211372
rect 269836 207890 269892 207900
rect 269724 26114 269780 26124
rect 270508 24612 270564 256088
rect 270620 250180 270676 250190
rect 270620 44884 270676 250124
rect 270844 246596 270900 246606
rect 270620 44818 270676 44828
rect 270732 243348 270788 243358
rect 270732 41524 270788 243292
rect 270844 44772 270900 246540
rect 271068 246484 271124 246494
rect 270956 246036 271012 246046
rect 270956 44996 271012 245980
rect 271068 48020 271124 246428
rect 271180 145348 271236 145358
rect 271180 49700 271236 145292
rect 271180 49634 271236 49644
rect 271068 47954 271124 47964
rect 270956 44930 271012 44940
rect 270844 44706 270900 44716
rect 270732 41458 270788 41468
rect 270508 24546 270564 24556
rect 271404 14532 271460 256088
rect 272300 252084 272356 256088
rect 272300 252018 272356 252028
rect 272188 251748 272244 251758
rect 272188 154084 272244 251692
rect 272972 245364 273028 245374
rect 272748 210196 272804 210206
rect 272524 210084 272580 210094
rect 272412 209860 272468 209870
rect 272188 154018 272244 154028
rect 272300 208740 272356 208750
rect 272300 140756 272356 208684
rect 272412 180852 272468 209804
rect 272412 180786 272468 180796
rect 272300 140690 272356 140700
rect 272524 153524 272580 210028
rect 272524 137172 272580 153468
rect 272524 137106 272580 137116
rect 272748 154420 272804 210140
rect 272748 134260 272804 154364
rect 272748 134194 272804 134204
rect 272972 153076 273028 245308
rect 273196 242676 273252 256088
rect 273868 255892 273924 255902
rect 273196 242610 273252 242620
rect 273420 243236 273476 243246
rect 272972 125524 273028 153020
rect 272972 125458 273028 125468
rect 273084 216244 273140 216254
rect 271404 14466 271460 14476
rect 272972 120148 273028 120158
rect 269612 6066 269668 6076
rect 272972 4900 273028 120092
rect 273084 109172 273140 216188
rect 273308 155428 273364 155438
rect 273084 93492 273140 109116
rect 273084 93426 273140 93436
rect 273196 154420 273252 154430
rect 273196 81844 273252 154364
rect 273308 96404 273364 155372
rect 273420 153188 273476 243180
rect 273420 131348 273476 153132
rect 273420 131282 273476 131292
rect 273644 154532 273700 154542
rect 273308 96338 273364 96348
rect 273644 90580 273700 154476
rect 273868 151732 273924 255836
rect 273980 250068 274036 250078
rect 273980 155428 274036 250012
rect 274092 234500 274148 256088
rect 274988 236068 275044 256088
rect 275660 253540 275716 253550
rect 274988 236002 275044 236012
rect 275548 253316 275604 253326
rect 274092 234434 274148 234444
rect 274876 213108 274932 213118
rect 273980 155362 274036 155372
rect 274652 211540 274708 211550
rect 273868 151666 273924 151676
rect 274652 152852 274708 211484
rect 274876 161308 274932 213052
rect 274876 161252 275380 161308
rect 275324 156436 275380 161252
rect 275324 154420 275380 156380
rect 275436 156324 275492 156334
rect 275436 154532 275492 156268
rect 275436 154466 275492 154476
rect 275324 154354 275380 154364
rect 274652 149548 274708 152796
rect 274652 149492 274820 149548
rect 273756 136164 273812 136174
rect 273756 128436 273812 136108
rect 273756 128370 273812 128380
rect 273644 90514 273700 90524
rect 274652 123508 274708 123518
rect 273196 81778 273252 81788
rect 273084 73108 273140 73118
rect 273084 52836 273140 73052
rect 273308 70196 273364 70206
rect 273084 52770 273140 52780
rect 273196 67284 273252 67294
rect 273196 50708 273252 67228
rect 273308 52724 273364 70140
rect 273308 52658 273364 52668
rect 273196 50642 273252 50652
rect 272972 4834 273028 4844
rect 274652 4340 274708 123452
rect 274764 99316 274820 149492
rect 274764 99250 274820 99260
rect 274876 121828 274932 121838
rect 274652 4274 274708 4284
rect 274876 4116 274932 121772
rect 275548 42980 275604 253260
rect 275660 49812 275716 253484
rect 275660 49746 275716 49756
rect 275548 42914 275604 42924
rect 275884 15988 275940 256088
rect 276332 152180 276388 152190
rect 276332 76020 276388 152124
rect 276332 75954 276388 75964
rect 276332 58548 276388 58558
rect 276332 50596 276388 58492
rect 276332 50530 276388 50540
rect 276780 17668 276836 256088
rect 276780 17602 276836 17612
rect 277228 253092 277284 253102
rect 275884 15922 275940 15932
rect 277228 10948 277284 253036
rect 277340 252980 277396 252990
rect 277340 45108 277396 252924
rect 277564 252308 277620 252318
rect 277452 252196 277508 252206
rect 277452 46228 277508 252140
rect 277564 48244 277620 252252
rect 277564 48178 277620 48188
rect 277452 46162 277508 46172
rect 277340 45042 277396 45052
rect 277676 19348 277732 256088
rect 278012 61460 278068 61470
rect 278012 50372 278068 61404
rect 278012 50306 278068 50316
rect 277676 19282 277732 19292
rect 277228 10882 277284 10892
rect 278572 9380 278628 256088
rect 279020 253204 279076 253214
rect 278908 252868 278964 252878
rect 278908 31332 278964 252812
rect 279020 39508 279076 253148
rect 279132 252084 279188 252094
rect 279132 45220 279188 252028
rect 279132 45154 279188 45164
rect 279020 39442 279076 39452
rect 278908 31266 278964 31276
rect 279468 24388 279524 256088
rect 279468 24322 279524 24332
rect 280364 14308 280420 256088
rect 281260 29428 281316 256088
rect 281372 252868 281428 252878
rect 281372 48356 281428 252812
rect 281372 48290 281428 48300
rect 282156 32900 282212 256088
rect 282156 32834 282212 32844
rect 281260 29362 281316 29372
rect 283052 19460 283108 256088
rect 283388 252980 283444 252990
rect 283164 252532 283220 252542
rect 283164 26068 283220 252476
rect 283388 41748 283444 252924
rect 283836 156548 283892 156558
rect 283836 152964 283892 156492
rect 283836 152898 283892 152908
rect 283388 41682 283444 41692
rect 283164 26002 283220 26012
rect 283052 19394 283108 19404
rect 280364 14242 280420 14252
rect 278572 9314 278628 9324
rect 283948 5908 284004 256088
rect 284732 253092 284788 253102
rect 284732 36260 284788 253036
rect 284732 36194 284788 36204
rect 284844 7588 284900 256088
rect 284956 253204 285012 253214
rect 284956 41636 285012 253148
rect 284956 41570 285012 41580
rect 285740 7700 285796 256088
rect 286412 210980 286468 210990
rect 286412 154532 286468 210924
rect 286412 102228 286468 154476
rect 286412 102162 286468 102172
rect 286636 7812 286692 256088
rect 287532 17780 287588 256088
rect 288316 253316 288372 253326
rect 288092 252084 288148 252094
rect 287980 55636 288036 55646
rect 287980 50484 288036 55580
rect 287980 50418 288036 50428
rect 288092 24500 288148 252028
rect 288316 49924 288372 253260
rect 288316 49858 288372 49868
rect 288092 24434 288148 24444
rect 287532 17714 287588 17724
rect 288428 16100 288484 256088
rect 289324 252084 289380 256088
rect 289324 252018 289380 252028
rect 289772 252756 289828 252766
rect 289772 29540 289828 252700
rect 289996 252308 290052 252318
rect 289884 216132 289940 216142
rect 289884 48580 289940 216076
rect 289884 48514 289940 48524
rect 289996 31220 290052 252252
rect 290108 64372 290164 64382
rect 290108 51828 290164 64316
rect 290108 51762 290164 51772
rect 289996 31154 290052 31164
rect 289772 29474 289828 29484
rect 288428 16034 288484 16044
rect 290220 14420 290276 256088
rect 290332 253428 290388 253438
rect 290332 38388 290388 253372
rect 291116 252532 291172 256088
rect 291116 252466 291172 252476
rect 292012 252420 292068 256088
rect 292012 252354 292068 252364
rect 290332 38322 290388 38332
rect 290892 252308 290948 252318
rect 290892 21028 290948 252252
rect 290892 20962 290948 20972
rect 291116 252196 291172 252206
rect 290220 14354 290276 14364
rect 291116 12628 291172 252140
rect 292908 252084 292964 256088
rect 293804 252196 293860 256088
rect 294700 252756 294756 256088
rect 295596 253204 295652 256088
rect 296492 253316 296548 256088
rect 296492 253250 296548 253260
rect 295596 253138 295652 253148
rect 294700 252690 294756 252700
rect 297388 252308 297444 256088
rect 298284 253428 298340 256088
rect 298284 253362 298340 253372
rect 299180 252868 299236 256088
rect 300076 252980 300132 256088
rect 300972 253092 301028 256088
rect 300972 253026 301028 253036
rect 300076 252914 300132 252924
rect 299180 252802 299236 252812
rect 297388 252242 297444 252252
rect 293804 252130 293860 252140
rect 301868 252196 301924 256088
rect 301868 252130 301924 252140
rect 292908 252018 292964 252028
rect 295148 154756 295204 154766
rect 295148 154308 295204 154700
rect 295148 154242 295204 154252
rect 293132 150388 293188 150398
rect 293132 110964 293188 150332
rect 302764 125412 302820 256088
rect 302764 125346 302820 125356
rect 303660 125300 303716 256088
rect 304556 252084 304612 256088
rect 304556 252018 304612 252028
rect 304892 252196 304948 252206
rect 303996 152964 304052 152974
rect 303996 150388 304052 152908
rect 303996 150322 304052 150332
rect 304892 133588 304948 252140
rect 305452 197428 305508 256088
rect 306348 217812 306404 256088
rect 306348 217746 306404 217756
rect 305452 197362 305508 197372
rect 304892 133522 304948 133532
rect 307244 126980 307300 256088
rect 307356 160692 307412 160702
rect 307356 152964 307412 160636
rect 307356 152898 307412 152908
rect 307244 126914 307300 126924
rect 308140 126868 308196 256088
rect 309036 231252 309092 256088
rect 309036 231186 309092 231196
rect 309932 192388 309988 256088
rect 310828 252868 310884 256088
rect 310828 252802 310884 252812
rect 309932 192322 309988 192332
rect 310044 252084 310100 252094
rect 308140 126802 308196 126812
rect 308252 154532 308308 154542
rect 303660 125234 303716 125244
rect 308252 113876 308308 154476
rect 308252 113810 308308 113820
rect 309932 151396 309988 151406
rect 293132 110898 293188 110908
rect 309932 84756 309988 151340
rect 310044 150612 310100 252028
rect 310940 160804 310996 160814
rect 310940 154532 310996 160748
rect 310940 154466 310996 154476
rect 310044 150546 310100 150556
rect 311724 131908 311780 256088
rect 312620 252980 312676 256088
rect 312620 252914 312676 252924
rect 313516 252084 313572 256088
rect 313516 252018 313572 252028
rect 314412 204148 314468 256088
rect 314972 252084 315028 252094
rect 314972 234500 315028 252028
rect 314972 234434 315028 234444
rect 314412 204082 314468 204092
rect 315308 138628 315364 256088
rect 316204 252084 316260 256088
rect 317100 252196 317156 256088
rect 317100 252130 317156 252140
rect 316204 252018 316260 252028
rect 315308 138562 315364 138572
rect 311724 131842 311780 131852
rect 317996 125188 318052 256088
rect 318332 252084 318388 252094
rect 318332 232932 318388 252028
rect 318892 252084 318948 256088
rect 319788 252420 319844 256088
rect 319788 252354 319844 252364
rect 320012 252980 320068 252990
rect 318892 252018 318948 252028
rect 318332 232866 318388 232876
rect 317996 125122 318052 125132
rect 318332 153748 318388 153758
rect 318332 119700 318388 153692
rect 320012 141988 320068 252924
rect 320236 252196 320292 252206
rect 320236 231140 320292 252140
rect 320236 231074 320292 231084
rect 320684 227780 320740 256088
rect 321580 252308 321636 256088
rect 321580 252242 321636 252252
rect 321692 252868 321748 252878
rect 320684 227714 320740 227724
rect 320012 141922 320068 141932
rect 321692 128548 321748 252812
rect 321916 252084 321972 252094
rect 321916 205828 321972 252028
rect 322476 234388 322532 256088
rect 322476 234322 322532 234332
rect 323372 222740 323428 256088
rect 323484 252420 323540 252430
rect 323484 229460 323540 252364
rect 323484 229394 323540 229404
rect 323372 222674 323428 222684
rect 324268 217700 324324 256088
rect 325164 252196 325220 256088
rect 325164 252130 325220 252140
rect 325388 252308 325444 252318
rect 325388 224420 325444 252252
rect 326060 252084 326116 256088
rect 326060 252018 326116 252028
rect 326732 254548 326788 254558
rect 325388 224354 325444 224364
rect 324268 217634 324324 217644
rect 325052 217812 325108 217822
rect 321916 205762 321972 205772
rect 321692 128482 321748 128492
rect 323372 153860 323428 153870
rect 323372 122612 323428 153804
rect 325052 123732 325108 217756
rect 325052 123666 325108 123676
rect 323372 122546 323428 122556
rect 318332 119634 318388 119644
rect 309932 84690 309988 84700
rect 307468 50260 307524 50270
rect 314188 50260 314244 50270
rect 321356 50260 321412 50270
rect 307524 50204 307944 50260
rect 314244 50204 315112 50260
rect 321412 50204 322280 50260
rect 307468 50194 307524 50204
rect 314188 50194 314244 50204
rect 321356 50194 321412 50204
rect 293580 50148 293636 50158
rect 293580 48692 293636 50092
rect 293580 48626 293636 48636
rect 300748 48580 300804 50120
rect 300748 48514 300804 48524
rect 326732 33684 326788 254492
rect 326844 252196 326900 252206
rect 326844 232820 326900 252140
rect 326844 232754 326900 232764
rect 326956 194180 327012 256088
rect 326956 194114 327012 194124
rect 327852 182420 327908 256088
rect 327852 182354 327908 182364
rect 328412 254548 328468 254558
rect 326732 33618 326788 33628
rect 291116 12562 291172 12572
rect 286636 7746 286692 7756
rect 285740 7634 285796 7644
rect 284844 7522 284900 7532
rect 283948 5842 284004 5852
rect 328412 4228 328468 254492
rect 328748 170660 328804 256088
rect 328748 170594 328804 170604
rect 329644 159012 329700 256088
rect 329644 158946 329700 158956
rect 330092 254660 330148 254670
rect 330092 4564 330148 254604
rect 330540 199220 330596 256088
rect 330540 199154 330596 199164
rect 331436 189028 331492 256088
rect 331436 188962 331492 188972
rect 331772 256004 331828 256014
rect 331772 4676 331828 255948
rect 331884 252084 331940 252094
rect 331884 210868 331940 252028
rect 332332 252084 332388 256088
rect 332332 252018 332388 252028
rect 331884 210802 331940 210812
rect 331884 192388 331940 192398
rect 331884 123620 331940 192332
rect 333228 158900 333284 256088
rect 333452 252084 333508 252094
rect 333452 162260 333508 252028
rect 334124 252084 334180 256088
rect 334124 252018 334180 252028
rect 333452 162194 333508 162204
rect 333228 158834 333284 158844
rect 335020 158788 335076 256088
rect 335132 252084 335188 252094
rect 335132 179060 335188 252028
rect 335916 192500 335972 256088
rect 336812 255388 336868 256088
rect 336812 255332 336980 255388
rect 335916 192434 335972 192444
rect 336812 254436 336868 254446
rect 335132 178994 335188 179004
rect 335020 158722 335076 158732
rect 331884 123554 331940 123564
rect 331772 4610 331828 4620
rect 330092 4498 330148 4508
rect 336812 4452 336868 254380
rect 336924 155764 336980 255332
rect 336924 155698 336980 155708
rect 337708 155652 337764 256088
rect 337708 155586 337764 155596
rect 338604 155540 338660 256088
rect 339500 187460 339556 256088
rect 339500 187394 339556 187404
rect 340396 163940 340452 256088
rect 341292 185668 341348 256088
rect 341292 185602 341348 185612
rect 342188 168868 342244 256088
rect 343084 252084 343140 256088
rect 343084 252018 343140 252028
rect 343980 236852 344036 256088
rect 343980 236786 344036 236796
rect 344876 199108 344932 256088
rect 345212 252084 345268 252094
rect 345212 200564 345268 252028
rect 345212 200498 345268 200508
rect 344876 199042 344932 199052
rect 345772 180628 345828 256088
rect 345772 180562 345828 180572
rect 342188 168802 342244 168812
rect 340396 163874 340452 163884
rect 346668 157332 346724 256088
rect 346668 157266 346724 157276
rect 347564 157220 347620 256088
rect 347564 157154 347620 157164
rect 348460 157108 348516 256088
rect 349356 195748 349412 256088
rect 349356 195682 349412 195692
rect 350252 177268 350308 256088
rect 350252 177202 350308 177212
rect 350476 256004 350532 256014
rect 348460 157042 348516 157052
rect 338604 155474 338660 155484
rect 350476 5012 350532 255948
rect 351148 175588 351204 256088
rect 351148 175522 351204 175532
rect 352044 173908 352100 256088
rect 352940 194068 352996 256088
rect 352940 194002 352996 194012
rect 353836 192388 353892 256088
rect 353836 192322 353892 192332
rect 354732 187348 354788 256088
rect 354732 187282 354788 187292
rect 355292 253316 355348 253326
rect 352044 173842 352100 173852
rect 355292 38276 355348 253260
rect 355628 252084 355684 256088
rect 355628 252018 355684 252028
rect 355740 248500 355796 248510
rect 355516 248388 355572 248398
rect 355292 38210 355348 38220
rect 355404 244692 355460 244702
rect 355404 31108 355460 244636
rect 355516 34580 355572 248332
rect 355740 35028 355796 248444
rect 356524 160580 356580 256088
rect 356972 252084 357028 252094
rect 356972 200676 357028 252028
rect 356972 200610 357028 200620
rect 357420 163828 357476 256088
rect 357420 163762 357476 163772
rect 358316 162148 358372 256088
rect 359212 255388 359268 256088
rect 359212 255332 359380 255388
rect 358316 162082 358372 162092
rect 358652 253428 358708 253438
rect 356524 160514 356580 160524
rect 356972 154308 357028 154318
rect 356972 141092 357028 154252
rect 356972 141026 357028 141036
rect 357756 151508 357812 151518
rect 357644 120260 357700 120270
rect 357644 84980 357700 120204
rect 357756 108948 357812 151452
rect 357756 108882 357812 108892
rect 357644 84914 357700 84924
rect 357756 61684 357812 61694
rect 356188 51940 356244 51950
rect 356188 50148 356244 51884
rect 357756 51940 357812 61628
rect 357756 51874 357812 51884
rect 356188 50082 356244 50092
rect 355740 34962 355796 34972
rect 358652 34804 358708 253372
rect 358988 251860 359044 251870
rect 358764 251748 358820 251758
rect 358764 44548 358820 251692
rect 358764 44482 358820 44492
rect 358988 38052 359044 251804
rect 358988 37986 359044 37996
rect 359212 251076 359268 251086
rect 359212 37940 359268 251020
rect 359324 182308 359380 255332
rect 359324 182242 359380 182252
rect 360108 160468 360164 256088
rect 361004 252868 361060 256088
rect 361004 252802 361060 252812
rect 361900 252196 361956 256088
rect 361900 252130 361956 252140
rect 360108 160402 360164 160412
rect 360332 248612 360388 248622
rect 359212 37874 359268 37884
rect 358652 34738 358708 34748
rect 355516 34514 355572 34524
rect 360332 34468 360388 248556
rect 360556 247716 360612 247726
rect 360556 37828 360612 247660
rect 362796 167188 362852 256088
rect 363692 252084 363748 256088
rect 364588 253092 364644 256088
rect 364588 253026 364644 253036
rect 363692 252018 363748 252028
rect 362796 167122 362852 167132
rect 362012 153636 362068 153646
rect 362012 142996 362068 153580
rect 365484 150388 365540 256088
rect 366380 252308 366436 256088
rect 367276 253204 367332 256088
rect 367276 253138 367332 253148
rect 366380 252242 366436 252252
rect 365484 150322 365540 150332
rect 367052 154532 367108 154542
rect 367052 145348 367108 154476
rect 368172 150500 368228 256088
rect 369068 252980 369124 256088
rect 369068 252914 369124 252924
rect 370412 252196 370468 252206
rect 370412 170548 370468 252140
rect 372092 252084 372148 252094
rect 370412 170482 370468 170492
rect 370748 197428 370804 197438
rect 368172 150434 368228 150444
rect 368732 150612 368788 150622
rect 367052 145282 367108 145292
rect 362012 142930 362068 142940
rect 362684 133588 362740 133598
rect 362684 119896 362740 133532
rect 364700 125412 364756 125422
rect 364700 119896 364756 125356
rect 366716 125300 366772 125310
rect 366716 119896 366772 125244
rect 368732 119896 368788 150556
rect 370748 119896 370804 197372
rect 372092 168980 372148 252028
rect 372092 168914 372148 168924
rect 375452 231252 375508 231262
rect 374780 126980 374836 126990
rect 372764 123732 372820 123742
rect 372764 119896 372820 123676
rect 374780 119896 374836 126924
rect 375452 122724 375508 231196
rect 375564 153524 375620 407708
rect 375676 154308 375732 407820
rect 375788 404852 375844 404862
rect 375788 154308 375844 404796
rect 375900 401492 375956 401502
rect 375900 154532 375956 401436
rect 383292 392196 383348 410088
rect 388668 402276 388724 410088
rect 394044 406308 394100 410088
rect 394044 406242 394100 406252
rect 388668 402210 388724 402220
rect 399420 393092 399476 410088
rect 404796 404740 404852 410088
rect 410172 407540 410228 410088
rect 410172 407474 410228 407484
rect 410732 407540 410788 407550
rect 404796 404674 404852 404684
rect 410732 394772 410788 407484
rect 415548 401044 415604 410088
rect 415548 400978 415604 400988
rect 410732 394706 410788 394716
rect 399420 393026 399476 393036
rect 383292 392130 383348 392140
rect 409276 391188 409332 391198
rect 409276 390964 409332 391132
rect 420924 391188 420980 410088
rect 426300 407540 426356 410088
rect 426300 407474 426356 407484
rect 431676 399700 431732 410088
rect 437052 404628 437108 410088
rect 437052 404562 437108 404572
rect 442428 403172 442484 410088
rect 442428 403106 442484 403116
rect 447804 400932 447860 410088
rect 451948 407540 452004 407550
rect 451948 406868 452004 407484
rect 451948 406802 452004 406812
rect 447804 400866 447860 400876
rect 431676 399634 431732 399644
rect 453180 398132 453236 410088
rect 453180 398066 453236 398076
rect 453516 407540 453572 407550
rect 420924 391122 420980 391132
rect 409276 390898 409332 390908
rect 421596 390852 421652 390862
rect 379820 390740 379876 390750
rect 377132 390516 377188 390526
rect 376348 383124 376404 383134
rect 376348 381332 376404 383068
rect 376348 381266 376404 381276
rect 377132 377188 377188 390460
rect 377132 377122 377188 377132
rect 377244 388388 377300 388398
rect 377132 297332 377188 297342
rect 376572 296212 376628 296222
rect 376348 276052 376404 276062
rect 376012 252084 376068 252094
rect 376012 175700 376068 252028
rect 376348 251860 376404 275996
rect 376348 251794 376404 251804
rect 376460 273812 376516 273822
rect 376460 251076 376516 273756
rect 376460 251010 376516 251020
rect 376572 227668 376628 296156
rect 376684 293972 376740 293982
rect 376684 248500 376740 293916
rect 376796 290612 376852 290622
rect 376796 253428 376852 290556
rect 377020 280532 377076 280542
rect 376796 253362 376852 253372
rect 376908 260372 376964 260382
rect 376684 248434 376740 248444
rect 376572 227602 376628 227612
rect 376908 224308 376964 260316
rect 377020 251748 377076 280476
rect 377020 251682 377076 251692
rect 376908 224242 376964 224252
rect 377132 222628 377188 297276
rect 377132 222562 377188 222572
rect 376012 175634 376068 175644
rect 375900 154466 375956 154476
rect 376124 154420 376180 154430
rect 376124 154308 376180 154364
rect 375788 154252 376180 154308
rect 375676 154242 375732 154252
rect 375564 153458 375620 153468
rect 376012 153860 376068 153870
rect 376012 153524 376068 153804
rect 376124 153636 376180 154252
rect 376236 154308 376292 154318
rect 376236 153748 376292 154252
rect 376236 153682 376292 153692
rect 376124 153570 376180 153580
rect 376012 153458 376068 153468
rect 375452 122658 375508 122668
rect 376796 126868 376852 126878
rect 376796 119896 376852 126812
rect 377244 120260 377300 388332
rect 379820 388164 379876 390684
rect 382172 390404 382228 390414
rect 379820 388098 379876 388108
rect 380492 390292 380548 390302
rect 379036 311892 379092 311902
rect 378924 310772 378980 310782
rect 378812 307412 378868 307422
rect 378364 292852 378420 292862
rect 378252 285012 378308 285022
rect 378028 282772 378084 282782
rect 378028 254436 378084 282716
rect 378140 274932 378196 274942
rect 378140 254548 378196 274876
rect 378252 254660 378308 284956
rect 378364 256116 378420 292796
rect 378476 291732 378532 291742
rect 378476 257348 378532 291676
rect 378476 257282 378532 257292
rect 378588 287252 378644 287262
rect 378588 256228 378644 287196
rect 378588 256162 378644 256172
rect 378700 279412 378756 279422
rect 378364 256050 378420 256060
rect 378252 254594 378308 254604
rect 378140 254482 378196 254492
rect 378028 254370 378084 254380
rect 378700 121828 378756 279356
rect 378812 275604 378868 307356
rect 378924 282212 378980 310716
rect 379036 284564 379092 311836
rect 379036 284498 379092 284508
rect 379708 295092 379764 295102
rect 378924 282146 378980 282156
rect 378812 275538 378868 275548
rect 378924 277172 378980 277182
rect 378700 121762 378756 121772
rect 378812 122724 378868 122734
rect 377244 120194 377300 120204
rect 378812 119896 378868 122668
rect 378924 120148 378980 277116
rect 379036 269332 379092 269342
rect 379036 123508 379092 269276
rect 379708 217588 379764 295036
rect 379820 284564 379876 284574
rect 379820 284004 379876 284508
rect 379820 256452 379876 283948
rect 379820 256386 379876 256396
rect 379932 282212 379988 282222
rect 379932 280644 379988 282156
rect 379932 254884 379988 280588
rect 380044 275604 380100 275614
rect 380044 254996 380100 275548
rect 380044 254930 380100 254940
rect 379932 254818 379988 254828
rect 379708 217522 379764 217532
rect 380492 178948 380548 390236
rect 380604 385812 380660 385822
rect 380604 337540 380660 385756
rect 380604 337474 380660 337484
rect 381388 268212 381444 268222
rect 381388 244692 381444 268156
rect 382172 258244 382228 390348
rect 421596 389396 421652 390796
rect 421596 389330 421652 389340
rect 429212 389956 429268 389966
rect 383852 387156 383908 387166
rect 383852 297892 383908 387100
rect 424172 387044 424228 387054
rect 383852 297826 383908 297836
rect 385532 386820 385588 386830
rect 382172 258178 382228 258188
rect 381388 244626 381444 244636
rect 385532 197204 385588 386764
rect 387212 386372 387268 386382
rect 387212 197316 387268 386316
rect 397292 386260 397348 386270
rect 387212 197250 387268 197260
rect 388892 234500 388948 234510
rect 385532 197138 385588 197148
rect 380492 178882 380548 178892
rect 386876 141988 386932 141998
rect 384860 131908 384916 131918
rect 382844 128548 382900 128558
rect 379036 123442 379092 123452
rect 380828 123620 380884 123630
rect 378924 120082 378980 120092
rect 380828 119896 380884 123564
rect 382844 119896 382900 128492
rect 384860 119896 384916 131852
rect 386876 119896 386932 141932
rect 388892 119896 388948 234444
rect 394940 232932 394996 232942
rect 390908 204148 390964 204158
rect 390908 119896 390964 204092
rect 392924 138628 392980 138638
rect 392924 119896 392980 138572
rect 394940 119896 394996 232876
rect 396956 231140 397012 231150
rect 396956 119896 397012 231084
rect 397292 197764 397348 386204
rect 398972 384580 399028 384590
rect 398972 197876 399028 384524
rect 400652 384468 400708 384478
rect 398972 197810 399028 197820
rect 399084 227780 399140 227790
rect 397292 197698 397348 197708
rect 398972 125188 399028 125198
rect 398972 119896 399028 125132
rect 399084 122724 399140 227724
rect 400652 197428 400708 384412
rect 414092 380212 414148 380222
rect 412412 253204 412468 253214
rect 407372 234388 407428 234398
rect 403004 229460 403060 229470
rect 400652 197362 400708 197372
rect 400988 205828 401044 205838
rect 399084 122658 399140 122668
rect 400988 119896 401044 205772
rect 403004 119896 403060 229404
rect 407036 224420 407092 224430
rect 405020 122724 405076 122734
rect 405020 119896 405076 122668
rect 407036 119896 407092 224364
rect 407372 124292 407428 234332
rect 411068 222740 411124 222750
rect 407372 124226 407428 124236
rect 409052 124292 409108 124302
rect 409052 119896 409108 124236
rect 411068 119896 411124 222684
rect 412412 150612 412468 253148
rect 412412 150546 412468 150556
rect 413084 217700 413140 217710
rect 413084 119896 413140 217644
rect 414092 199892 414148 380156
rect 415772 379092 415828 379102
rect 414092 199826 414148 199836
rect 415100 232820 415156 232830
rect 415100 119896 415156 232764
rect 415772 200004 415828 379036
rect 417452 376852 417508 376862
rect 415772 199938 415828 199948
rect 417116 210868 417172 210878
rect 417116 119896 417172 210812
rect 417452 199780 417508 376796
rect 417452 199714 417508 199724
rect 420028 101556 420084 101566
rect 420028 52836 420084 101500
rect 420028 52770 420084 52780
rect 420140 94948 420196 94958
rect 420140 52724 420196 94892
rect 420140 52658 420196 52668
rect 420252 88228 420308 88238
rect 420252 50708 420308 88172
rect 421708 81508 421764 81518
rect 421708 51828 421764 81452
rect 421708 51762 421764 51772
rect 421820 74788 421876 74798
rect 420252 50642 420308 50652
rect 421820 50372 421876 74732
rect 421932 68068 421988 68078
rect 421932 50596 421988 68012
rect 421932 50530 421988 50540
rect 422044 61348 422100 61358
rect 422044 50484 422100 61292
rect 422044 50418 422100 50428
rect 421820 50306 421876 50316
rect 360556 37762 360612 37772
rect 360332 34402 360388 34412
rect 355404 31042 355460 31052
rect 424172 20356 424228 386988
rect 424172 20290 424228 20300
rect 350476 4946 350532 4956
rect 336812 4386 336868 4396
rect 328412 4162 328468 4172
rect 429212 4228 429268 389900
rect 453516 195972 453572 407484
rect 458556 399588 458612 410088
rect 458556 399522 458612 399532
rect 463932 390964 463988 410088
rect 468748 410060 469336 410116
rect 468748 408268 468804 410060
rect 468636 408212 468804 408268
rect 468636 404516 468692 408212
rect 468636 404450 468692 404460
rect 472892 407876 472948 407886
rect 472892 392980 472948 407820
rect 474684 406196 474740 410088
rect 478380 407764 478436 407774
rect 474684 406130 474740 406140
rect 476252 407652 476308 407662
rect 472892 392914 472948 392924
rect 463932 390898 463988 390908
rect 474572 386708 474628 386718
rect 472892 385700 472948 385710
rect 467852 377972 467908 377982
rect 457772 375732 457828 375742
rect 457772 200228 457828 375676
rect 457772 200162 457828 200172
rect 459452 374612 459508 374622
rect 459452 199444 459508 374556
rect 461132 373492 461188 373502
rect 461132 200340 461188 373436
rect 461132 200274 461188 200284
rect 462812 372372 462868 372382
rect 459452 199378 459508 199388
rect 462812 198996 462868 372316
rect 464492 215908 464548 215918
rect 464492 206724 464548 215852
rect 464492 206658 464548 206668
rect 465948 206724 466004 206734
rect 465948 199668 466004 206668
rect 467852 200452 467908 377916
rect 467852 200386 467908 200396
rect 467964 249620 468020 249630
rect 465948 199602 466004 199612
rect 466284 199668 466340 199678
rect 462812 198930 462868 198940
rect 453516 195906 453572 195916
rect 456092 151956 456148 151966
rect 451052 151732 451108 151742
rect 437612 151620 437668 151630
rect 437612 94948 437668 151564
rect 437612 94882 437668 94892
rect 449372 149492 449428 149502
rect 449372 81508 449428 149436
rect 451052 88228 451108 151676
rect 451052 88162 451108 88172
rect 452732 149268 452788 149278
rect 449372 81442 449428 81452
rect 452732 68068 452788 149212
rect 452732 68002 452788 68012
rect 454412 148708 454468 148718
rect 454412 52948 454468 148652
rect 456092 61348 456148 151900
rect 456316 151844 456372 151854
rect 456316 101668 456372 151788
rect 456316 101602 456372 101612
rect 459452 151284 459508 151294
rect 459452 74788 459508 151228
rect 466284 149940 466340 199612
rect 467964 199556 468020 249564
rect 467964 196588 468020 199500
rect 472892 197540 472948 385644
rect 472892 197474 472948 197484
rect 473004 200900 473060 200910
rect 467852 196532 468020 196588
rect 467852 151956 467908 196532
rect 471660 195860 471716 195870
rect 467852 149940 467908 151900
rect 465724 149912 466340 149940
rect 465724 149884 466312 149912
rect 467656 149884 467908 149940
rect 468972 162372 469028 162382
rect 465724 149492 465780 149884
rect 468972 149716 469028 162316
rect 470316 160916 470372 160926
rect 470316 151284 470372 160860
rect 471660 156268 471716 195804
rect 471660 156212 471940 156268
rect 470316 149912 470372 151228
rect 468972 149650 469028 149660
rect 465724 149426 465780 149436
rect 471884 149492 471940 156212
rect 473004 151732 473060 200844
rect 474572 197652 474628 386652
rect 474572 197586 474628 197596
rect 474684 199332 474740 199342
rect 473004 149912 473060 151676
rect 474684 151620 474740 199276
rect 474684 149940 474740 151564
rect 474376 149884 474740 149940
rect 475692 161028 475748 161038
rect 475692 151844 475748 160972
rect 475692 149912 475748 151788
rect 476252 152180 476308 407596
rect 477932 385588 477988 385598
rect 477932 197988 477988 385532
rect 477932 197922 477988 197932
rect 476252 149940 476308 152124
rect 476252 149884 477064 149940
rect 478380 149912 478436 407708
rect 480060 403060 480116 410088
rect 484652 407988 484708 407998
rect 480060 402994 480116 403004
rect 480508 407428 480564 407438
rect 479612 385476 479668 385486
rect 479612 198212 479668 385420
rect 479612 198146 479668 198156
rect 479724 156436 479780 156446
rect 479724 149912 479780 156380
rect 480508 151396 480564 407372
rect 484652 392868 484708 407932
rect 485436 407876 485492 410088
rect 485436 407810 485492 407820
rect 484652 392802 484708 392812
rect 484876 392868 484932 392878
rect 484876 389284 484932 392812
rect 490812 392756 490868 410088
rect 496188 407988 496244 410088
rect 496188 407922 496244 407932
rect 490812 392690 490868 392700
rect 499772 406868 499828 406878
rect 499772 392644 499828 406812
rect 501564 406868 501620 410088
rect 501564 406802 501620 406812
rect 499772 392578 499828 392588
rect 506940 392532 506996 410088
rect 512316 400820 512372 410088
rect 512316 400754 512372 400764
rect 517692 398020 517748 410088
rect 519820 407988 519876 407998
rect 519708 407876 519764 407886
rect 519372 406756 519428 406766
rect 519260 406644 519316 406654
rect 517692 397954 517748 397964
rect 519148 403620 519204 403630
rect 506940 392466 506996 392476
rect 484876 389218 484932 389228
rect 517468 384244 517524 384254
rect 481628 251636 481684 251646
rect 481628 236936 481684 251580
rect 482748 251524 482804 251534
rect 482748 236936 482804 251468
rect 497308 251412 497364 251422
rect 484988 249956 485044 249966
rect 483868 244580 483924 244590
rect 483868 236936 483924 244524
rect 484988 236936 485044 249900
rect 495068 249844 495124 249854
rect 492828 248276 492884 248286
rect 488348 248164 488404 248174
rect 487228 246260 487284 246270
rect 486108 241556 486164 241566
rect 486108 236936 486164 241500
rect 487228 236936 487284 246204
rect 488348 236936 488404 248108
rect 491708 244468 491764 244478
rect 489468 239988 489524 239998
rect 489468 236936 489524 239932
rect 490588 237748 490644 237758
rect 490588 236936 490644 237692
rect 491708 236936 491764 244412
rect 492828 236936 492884 248220
rect 493948 243124 494004 243134
rect 493948 236936 494004 243068
rect 495068 236936 495124 249788
rect 496188 241444 496244 241454
rect 496188 236936 496244 241388
rect 497308 236936 497364 251356
rect 506268 251300 506324 251310
rect 502908 249732 502964 249742
rect 498428 248052 498484 248062
rect 498428 236936 498484 247996
rect 499548 243012 499604 243022
rect 499548 236936 499604 242956
rect 501788 241332 501844 241342
rect 500668 239876 500724 239886
rect 500668 236936 500724 239820
rect 501788 236936 501844 241276
rect 502908 236936 502964 249676
rect 504028 247940 504084 247950
rect 504028 236936 504084 247884
rect 505148 242900 505204 242910
rect 505148 236936 505204 242844
rect 506268 236936 506324 251244
rect 515228 251188 515284 251198
rect 508508 249508 508564 249518
rect 507388 239764 507444 239774
rect 507388 236936 507444 239708
rect 508508 236936 508564 249452
rect 511868 247828 511924 247838
rect 509628 246148 509684 246158
rect 509628 236936 509684 246092
rect 510748 241220 510804 241230
rect 510748 236936 510804 241164
rect 511868 236936 511924 247772
rect 514108 242788 514164 242798
rect 512988 239652 513044 239662
rect 512988 236936 513044 239596
rect 514108 236936 514164 242732
rect 515228 236936 515284 251132
rect 517468 231924 517524 384188
rect 517468 231858 517524 231868
rect 517580 229236 517636 229246
rect 517468 226548 517524 226558
rect 511644 200452 511700 200462
rect 505372 200340 505428 200350
rect 507948 200340 508004 200350
rect 505428 200284 505540 200340
rect 505372 200274 505428 200284
rect 488124 200116 488180 200126
rect 481852 197204 481908 200088
rect 483420 197764 483476 200088
rect 483420 197698 483476 197708
rect 484988 197316 485044 200088
rect 486556 197876 486612 200088
rect 488124 200050 488180 200060
rect 486556 197810 486612 197820
rect 489692 197428 489748 200088
rect 491260 197652 491316 200088
rect 491260 197586 491316 197596
rect 492828 197540 492884 200088
rect 494396 198212 494452 200088
rect 494396 198146 494452 198156
rect 495964 197988 496020 200088
rect 497532 198212 497588 200088
rect 497532 198146 497588 198156
rect 499100 198212 499156 200088
rect 499100 198146 499156 198156
rect 500668 198100 500724 200088
rect 502236 198212 502292 200088
rect 502236 198146 502292 198156
rect 503132 198996 503188 199006
rect 500668 198034 500724 198044
rect 495964 197922 496020 197932
rect 492828 197474 492884 197484
rect 489692 197362 489748 197372
rect 484988 197250 485044 197260
rect 481852 197138 481908 197148
rect 480508 149940 480564 151340
rect 482412 195972 482468 195982
rect 480508 149884 481096 149940
rect 482412 149912 482468 195916
rect 494508 160804 494564 160814
rect 493164 160692 493220 160702
rect 491820 156660 491876 156670
rect 487788 156548 487844 156558
rect 483756 156324 483812 156334
rect 483756 149912 483812 156268
rect 486444 155428 486500 155438
rect 485100 151508 485156 151518
rect 485100 149912 485156 151452
rect 486444 149912 486500 155372
rect 487788 149912 487844 156492
rect 490476 154756 490532 154766
rect 489132 154644 489188 154654
rect 489132 149912 489188 154588
rect 490476 149912 490532 154700
rect 491820 149912 491876 156604
rect 493164 149912 493220 160636
rect 494508 149912 494564 160748
rect 497196 154196 497252 154206
rect 495852 152964 495908 152974
rect 495852 149912 495908 152908
rect 497196 149912 497252 154140
rect 498540 154084 498596 154094
rect 498540 149912 498596 154028
rect 502572 153188 502628 153198
rect 499884 153076 499940 153086
rect 499884 149912 499940 153020
rect 501340 152964 501396 152974
rect 501396 152908 501508 152964
rect 501340 152898 501396 152908
rect 501452 149828 501508 152908
rect 502572 149912 502628 153132
rect 503132 152068 503188 198940
rect 503804 198996 503860 200088
rect 503804 198930 503860 198940
rect 503132 152002 503188 152012
rect 503916 153972 503972 153982
rect 503916 149912 503972 153916
rect 505260 153860 505316 153870
rect 505260 149912 505316 153804
rect 501256 149772 501508 149828
rect 471884 149426 471940 149436
rect 505484 149492 505540 200284
rect 506492 199444 506548 199454
rect 506492 150724 506548 199388
rect 506940 199444 506996 200088
rect 506940 199378 506996 199388
rect 506828 194180 506884 194190
rect 506828 154532 506884 194124
rect 506828 154466 506884 154476
rect 507948 154196 508004 200284
rect 508508 200228 508564 200238
rect 508508 161308 508564 200172
rect 509852 200088 510104 200116
rect 509852 200060 510132 200088
rect 508508 161252 508900 161308
rect 506492 150658 506548 150668
rect 506604 153748 506660 153758
rect 506604 149912 506660 153692
rect 507948 149912 508004 154140
rect 508844 149604 508900 161252
rect 509852 152180 509908 200060
rect 510076 199780 510132 200060
rect 510076 199714 510132 199724
rect 510300 199444 510356 199454
rect 510300 161308 510356 199388
rect 509852 152114 509908 152124
rect 510076 161252 510356 161308
rect 510076 154420 510132 161252
rect 510076 149940 510132 154364
rect 509320 149884 510132 149940
rect 510636 154532 510692 154542
rect 510636 149912 510692 154476
rect 511644 152292 511700 200396
rect 512428 200088 513240 200116
rect 512428 200060 513268 200088
rect 514808 200060 514948 200116
rect 512428 200004 512484 200060
rect 512428 199938 512484 199948
rect 511644 152226 511700 152236
rect 511980 182420 512036 182430
rect 511980 149912 512036 182364
rect 513212 155428 513268 200060
rect 514892 199892 514948 200060
rect 513436 199220 513492 199230
rect 513212 155362 513268 155372
rect 513324 170660 513380 170670
rect 513324 149912 513380 170604
rect 513436 154532 513492 199164
rect 513436 154466 513492 154476
rect 514668 159012 514724 159022
rect 514668 149912 514724 158956
rect 514892 159012 514948 199836
rect 514892 158946 514948 158956
rect 515004 192500 515060 192510
rect 515004 154420 515060 192444
rect 517356 189028 517412 189038
rect 515004 154354 515060 154364
rect 516012 154532 516068 154542
rect 516012 149912 516068 154476
rect 517356 149912 517412 188972
rect 517468 161028 517524 226492
rect 517580 200340 517636 229180
rect 517580 200274 517636 200284
rect 517692 223860 517748 223870
rect 517692 199332 517748 223804
rect 517804 221732 517860 221742
rect 517804 200900 517860 221676
rect 519148 221732 519204 403564
rect 519260 226100 519316 406588
rect 519372 226548 519428 406700
rect 519708 406644 519764 407820
rect 519820 406756 519876 407932
rect 519820 406690 519876 406700
rect 519708 406578 519764 406588
rect 523068 399476 523124 410088
rect 527548 410060 528472 410116
rect 527548 408268 527604 410060
rect 527436 408212 527604 408268
rect 527436 404404 527492 408212
rect 527436 404338 527492 404348
rect 533820 402948 533876 410088
rect 533820 402882 533876 402892
rect 523068 399410 523124 399420
rect 539196 392420 539252 410088
rect 544572 406084 544628 410088
rect 544572 406018 544628 406028
rect 539196 392354 539252 392364
rect 548492 388948 548548 410508
rect 549388 395556 549444 550396
rect 549500 512820 549556 512830
rect 549500 409668 549556 512764
rect 549500 409602 549556 409612
rect 549612 484484 549668 484494
rect 549388 395490 549444 395500
rect 549612 394548 549668 484428
rect 549612 394482 549668 394492
rect 549724 475524 549780 475534
rect 549724 394212 549780 475468
rect 549836 397460 549892 590716
rect 550060 570388 550116 570398
rect 549836 397394 549892 397404
rect 549948 465668 550004 465678
rect 549724 394146 549780 394156
rect 549948 393988 550004 465612
rect 550060 407428 550116 570332
rect 552748 565124 552804 565134
rect 551852 560308 551908 560318
rect 551180 508676 551236 508686
rect 550284 482916 550340 482926
rect 550060 407362 550116 407372
rect 550172 419300 550228 419310
rect 550172 400708 550228 419244
rect 550284 407988 550340 482860
rect 550284 407922 550340 407932
rect 551068 414596 551124 414606
rect 550172 400642 550228 400652
rect 551068 397796 551124 414540
rect 551180 404180 551236 508620
rect 551180 404114 551236 404124
rect 551292 480452 551348 480462
rect 551068 397730 551124 397740
rect 551292 394324 551348 480396
rect 551292 394258 551348 394268
rect 551404 471044 551460 471054
rect 551404 394100 551460 470988
rect 551516 461636 551572 461646
rect 551516 399252 551572 461580
rect 551628 442820 551684 442830
rect 551628 409332 551684 442764
rect 551628 409266 551684 409276
rect 551740 424004 551796 424014
rect 551516 399186 551572 399196
rect 551740 395780 551796 423948
rect 551852 407764 551908 560252
rect 551852 407698 551908 407708
rect 551964 536900 552020 536910
rect 551740 395714 551796 395724
rect 551404 394034 551460 394044
rect 549948 393922 550004 393932
rect 551964 392308 552020 536844
rect 551964 392242 552020 392252
rect 552748 390740 552804 565068
rect 556108 560420 556164 560430
rect 552860 555716 552916 555726
rect 552860 390852 552916 555660
rect 553532 546308 553588 546318
rect 552972 541604 553028 541614
rect 552972 409892 553028 541548
rect 553196 456932 553252 456942
rect 552972 409826 553028 409836
rect 553084 438116 553140 438126
rect 553084 392868 553140 438060
rect 553196 410564 553252 456876
rect 553196 410498 553252 410508
rect 553308 452228 553364 452238
rect 553308 409444 553364 452172
rect 553532 452004 553588 546252
rect 553532 451938 553588 451948
rect 554428 522788 554484 522798
rect 553420 447524 553476 447534
rect 553420 409556 553476 447468
rect 553420 409490 553476 409500
rect 553532 433412 553588 433422
rect 553308 409378 553364 409388
rect 553532 395892 553588 433356
rect 554428 405860 554484 522732
rect 555212 522564 555268 522574
rect 554428 405794 554484 405804
rect 554540 503972 554596 503982
rect 554540 396116 554596 503916
rect 554540 396050 554596 396060
rect 554652 499268 554708 499278
rect 554652 396004 554708 499212
rect 554652 395938 554708 395948
rect 554764 489860 554820 489870
rect 553532 395826 553588 395836
rect 554764 394436 554820 489804
rect 554764 394370 554820 394380
rect 554876 452004 554932 452014
rect 553084 392802 553140 392812
rect 552860 390786 552916 390796
rect 552748 390674 552804 390684
rect 554876 389060 554932 451948
rect 554988 428708 555044 428718
rect 554988 395668 555044 428652
rect 555212 407652 555268 522508
rect 555212 407586 555268 407596
rect 554988 395602 555044 395612
rect 556108 389172 556164 560364
rect 556444 532196 556500 532206
rect 556220 527492 556276 527502
rect 556220 394660 556276 527436
rect 556220 394594 556276 394604
rect 556332 518084 556388 518094
rect 556332 390628 556388 518028
rect 556444 409780 556500 532140
rect 556444 409714 556500 409724
rect 556556 494564 556612 494574
rect 556556 402724 556612 494508
rect 556556 402658 556612 402668
rect 556892 416836 556948 416846
rect 556892 399140 556948 416780
rect 556892 399074 556948 399084
rect 560252 397684 560308 591276
rect 562604 591332 562660 595560
rect 562604 591266 562660 591276
rect 566972 575428 567028 575438
rect 560252 397618 560308 397628
rect 563612 535780 563668 535790
rect 563612 397572 563668 535724
rect 565292 456484 565348 456494
rect 565292 404068 565348 456428
rect 566972 405748 567028 575372
rect 566972 405682 567028 405692
rect 583772 496132 583828 496142
rect 565292 404002 565348 404012
rect 583772 402612 583828 496076
rect 584668 409108 584724 595560
rect 591276 562212 591332 562222
rect 591276 560308 591332 562156
rect 591276 560242 591332 560252
rect 584668 409042 584724 409052
rect 587132 443268 587188 443278
rect 587132 407876 587188 443212
rect 587132 407810 587188 407820
rect 583772 402546 583828 402556
rect 563612 397506 563668 397516
rect 556332 390562 556388 390572
rect 556108 389106 556164 389116
rect 578732 389844 578788 389854
rect 554876 388994 554932 389004
rect 548492 388882 548548 388892
rect 521612 386596 521668 386606
rect 519932 383236 519988 383246
rect 519932 344372 519988 383180
rect 519372 226482 519428 226492
rect 519484 246932 519540 246942
rect 519484 245924 519540 246876
rect 519260 226044 519428 226100
rect 519372 223860 519428 226044
rect 519372 223794 519428 223804
rect 519484 223636 519540 245868
rect 519148 221666 519204 221676
rect 519260 223580 519540 223636
rect 519260 213108 519316 223580
rect 519932 220108 519988 344316
rect 517804 200834 517860 200844
rect 519148 207732 519204 207742
rect 519148 205380 519204 207676
rect 519148 199780 519204 205324
rect 519148 199714 519204 199724
rect 517692 199266 517748 199276
rect 519260 162372 519316 213052
rect 519372 220052 519988 220108
rect 520044 324324 520100 324334
rect 519372 218484 519428 220052
rect 519372 195860 519428 218428
rect 519596 215796 519652 215806
rect 520044 215796 520100 324268
rect 520156 284676 520212 284686
rect 520156 246932 520212 284620
rect 520156 246866 520212 246876
rect 521612 218596 521668 386540
rect 521612 218530 521668 218540
rect 523292 253092 523348 253102
rect 519652 215740 520100 215796
rect 519484 210868 519540 210878
rect 519484 199556 519540 210812
rect 519484 199490 519540 199500
rect 519372 195794 519428 195804
rect 519260 162306 519316 162316
rect 517468 160962 517524 160972
rect 518700 162260 518756 162270
rect 518700 149912 518756 162204
rect 519596 160916 519652 215740
rect 519596 160850 519652 160860
rect 521388 179060 521444 179070
rect 520044 158900 520100 158910
rect 520044 149912 520100 158844
rect 521388 149912 521444 179004
rect 522732 158788 522788 158798
rect 522732 149912 522788 158732
rect 523292 152404 523348 253036
rect 548492 252980 548548 252990
rect 536172 236852 536228 236862
rect 534828 200564 534884 200574
rect 533372 199108 533428 199118
rect 529452 187460 529508 187470
rect 526652 185668 526708 185678
rect 525420 155764 525476 155774
rect 523292 152338 523348 152348
rect 524076 154420 524132 154430
rect 524076 149912 524132 154364
rect 525420 149912 525476 155708
rect 526652 154532 526708 185612
rect 526652 154466 526708 154476
rect 526764 155652 526820 155662
rect 526764 149912 526820 155596
rect 528108 155540 528164 155550
rect 528108 149912 528164 155484
rect 529452 149912 529508 187404
rect 530796 163940 530852 163950
rect 530796 149912 530852 163884
rect 532140 154532 532196 154542
rect 532140 149912 532196 154476
rect 533372 154532 533428 199052
rect 533372 154466 533428 154476
rect 533484 168868 533540 168878
rect 533484 149912 533540 168812
rect 534828 149912 534884 200508
rect 536172 149912 536228 236796
rect 544236 195748 544292 195758
rect 538860 180628 538916 180638
rect 537516 154532 537572 154542
rect 537516 149912 537572 154476
rect 538860 149912 538916 180572
rect 541772 175588 541828 175598
rect 540204 157332 540260 157342
rect 540204 149912 540260 157276
rect 541548 157220 541604 157230
rect 541548 149912 541604 157164
rect 541772 154532 541828 175532
rect 541772 154466 541828 154476
rect 542892 157108 542948 157118
rect 542892 149912 542948 157052
rect 544236 149912 544292 195692
rect 547148 192388 547204 192398
rect 545580 177268 545636 177278
rect 545580 149912 545636 177212
rect 546924 154532 546980 154542
rect 546924 149912 546980 154476
rect 547148 154532 547204 192332
rect 547148 154466 547204 154476
rect 548268 173908 548324 173918
rect 548268 149912 548324 173852
rect 548492 150836 548548 252924
rect 560252 252868 560308 252878
rect 553644 200676 553700 200686
rect 548492 150770 548548 150780
rect 549612 194068 549668 194078
rect 549612 149912 549668 194012
rect 552300 187348 552356 187358
rect 550956 154532 551012 154542
rect 550956 149912 551012 154476
rect 552300 149912 552356 187292
rect 553644 149912 553700 200620
rect 559468 182308 559524 182318
rect 508844 149538 508900 149548
rect 505484 149426 505540 149436
rect 459900 149380 459956 149390
rect 459900 148708 459956 149324
rect 471660 149268 471716 149278
rect 471660 149202 471716 149212
rect 459900 148642 459956 148652
rect 559468 113764 559524 182252
rect 559468 113698 559524 113708
rect 559580 163828 559636 163838
rect 559580 110628 559636 163772
rect 559804 162148 559860 162158
rect 559580 110562 559636 110572
rect 559692 160580 559748 160590
rect 559692 109172 559748 160524
rect 559804 112196 559860 162092
rect 559916 150500 559972 150510
rect 559916 127652 559972 150444
rect 559916 127586 559972 127596
rect 560252 122500 560308 252812
rect 565292 236628 565348 236638
rect 562828 175700 562884 175710
rect 561708 159012 561764 159022
rect 561372 155428 561428 155438
rect 561148 152180 561204 152190
rect 561148 136724 561204 152124
rect 561148 136658 561204 136668
rect 561260 149492 561316 149502
rect 561260 132020 561316 149436
rect 561372 139860 561428 155372
rect 561596 152292 561652 152302
rect 561372 139794 561428 139804
rect 561484 149268 561540 149278
rect 561484 135156 561540 149212
rect 561596 138292 561652 152236
rect 561708 141428 561764 158956
rect 561708 141362 561764 141372
rect 561596 138226 561652 138236
rect 561484 135090 561540 135100
rect 561260 131954 561316 131964
rect 562828 124180 562884 175644
rect 563164 170548 563220 170558
rect 562828 124114 562884 124124
rect 562940 168980 562996 168990
rect 560252 122434 560308 122444
rect 562828 122500 562884 122510
rect 562828 116340 562884 122444
rect 562940 119476 562996 168924
rect 563052 152404 563108 152414
rect 563052 121044 563108 152348
rect 563164 142996 563220 170492
rect 564508 160468 564564 160478
rect 563388 150836 563444 150846
rect 563164 142930 563220 142940
rect 563276 150612 563332 150622
rect 563276 125748 563332 150556
rect 563388 128884 563444 150780
rect 563388 128818 563444 128828
rect 563276 125682 563332 125692
rect 563052 120978 563108 120988
rect 562940 119410 562996 119420
rect 562828 116274 562884 116284
rect 564508 114772 564564 160412
rect 564732 150724 564788 150734
rect 564620 150388 564676 150398
rect 564620 122612 564676 150332
rect 564732 133588 564788 150668
rect 564732 133522 564788 133532
rect 564620 122546 564676 122556
rect 564508 114706 564564 114716
rect 559804 112130 559860 112140
rect 559692 109106 559748 109116
rect 459452 74722 459508 74732
rect 456092 61282 456148 61292
rect 454412 52882 454468 52892
rect 565292 7140 565348 236572
rect 566188 167188 566244 167198
rect 566188 117908 566244 167132
rect 566300 152068 566356 152078
rect 566300 130452 566356 152012
rect 578732 139300 578788 389788
rect 578732 139234 578788 139244
rect 585452 386484 585508 386494
rect 566300 130386 566356 130396
rect 566188 117842 566244 117852
rect 585452 99876 585508 386428
rect 587132 363972 587188 363982
rect 587132 344372 587188 363916
rect 587132 344306 587188 344316
rect 587132 245028 587188 245038
rect 587132 210868 587188 244972
rect 587132 210802 587188 210812
rect 585452 99810 585508 99820
rect 565292 7074 565348 7084
rect 429212 4162 429268 4172
rect 580636 4228 580692 4238
rect 274876 4050 274932 4060
rect 580636 480 580692 4172
rect 584444 4228 584500 4238
rect 582540 4116 582596 4126
rect 582540 480 582596 4060
rect 584444 480 584500 4172
rect 207452 392 207704 480
rect 209356 392 209608 480
rect 211260 392 211512 480
rect 205576 -960 205800 392
rect 207480 -960 207704 392
rect 209384 -960 209608 392
rect 211288 -960 211512 392
rect 213192 -960 213416 480
rect 215096 -960 215320 480
rect 217000 -960 217224 480
rect 218904 -960 219128 480
rect 220808 -960 221032 480
rect 222712 -960 222936 480
rect 224616 -960 224840 480
rect 226520 -960 226744 480
rect 228424 -960 228648 480
rect 230328 -960 230552 480
rect 232232 -960 232456 480
rect 234136 -960 234360 480
rect 236040 -960 236264 480
rect 237944 -960 238168 480
rect 239848 -960 240072 480
rect 241752 -960 241976 480
rect 243656 -960 243880 480
rect 245560 -960 245784 480
rect 247464 -960 247688 480
rect 249368 -960 249592 480
rect 251272 -960 251496 480
rect 253176 -960 253400 480
rect 255080 -960 255304 480
rect 256984 -960 257208 480
rect 258888 -960 259112 480
rect 260792 -960 261016 480
rect 262696 -960 262920 480
rect 264600 -960 264824 480
rect 266504 -960 266728 480
rect 268408 -960 268632 480
rect 270312 -960 270536 480
rect 272216 -960 272440 480
rect 274120 -960 274344 480
rect 276024 -960 276248 480
rect 277928 -960 278152 480
rect 279832 -960 280056 480
rect 281736 -960 281960 480
rect 283640 -960 283864 480
rect 285544 -960 285768 480
rect 287448 -960 287672 480
rect 289352 -960 289576 480
rect 291256 -960 291480 480
rect 293160 -960 293384 480
rect 295064 -960 295288 480
rect 296968 -960 297192 480
rect 298872 -960 299096 480
rect 300776 -960 301000 480
rect 302680 -960 302904 480
rect 304584 -960 304808 480
rect 306488 -960 306712 480
rect 308392 -960 308616 480
rect 310296 -960 310520 480
rect 312200 -960 312424 480
rect 314104 -960 314328 480
rect 316008 -960 316232 480
rect 317912 -960 318136 480
rect 319816 -960 320040 480
rect 321720 -960 321944 480
rect 323624 -960 323848 480
rect 325528 -960 325752 480
rect 327432 -960 327656 480
rect 329336 -960 329560 480
rect 331240 -960 331464 480
rect 333144 -960 333368 480
rect 335048 -960 335272 480
rect 336952 -960 337176 480
rect 338856 -960 339080 480
rect 340760 -960 340984 480
rect 342664 -960 342888 480
rect 344568 -960 344792 480
rect 346472 -960 346696 480
rect 348376 -960 348600 480
rect 350280 -960 350504 480
rect 352184 -960 352408 480
rect 354088 -960 354312 480
rect 355992 -960 356216 480
rect 357896 -960 358120 480
rect 359800 -960 360024 480
rect 361704 -960 361928 480
rect 363608 -960 363832 480
rect 365512 -960 365736 480
rect 367416 -960 367640 480
rect 369320 -960 369544 480
rect 371224 -960 371448 480
rect 373128 -960 373352 480
rect 375032 -960 375256 480
rect 376936 -960 377160 480
rect 378840 -960 379064 480
rect 380744 -960 380968 480
rect 382648 -960 382872 480
rect 384552 -960 384776 480
rect 386456 -960 386680 480
rect 388360 -960 388584 480
rect 390264 -960 390488 480
rect 392168 -960 392392 480
rect 394072 -960 394296 480
rect 395976 -960 396200 480
rect 397880 -960 398104 480
rect 399784 -960 400008 480
rect 401688 -960 401912 480
rect 403592 -960 403816 480
rect 405496 -960 405720 480
rect 407400 -960 407624 480
rect 409304 -960 409528 480
rect 411208 -960 411432 480
rect 413112 -960 413336 480
rect 415016 -960 415240 480
rect 416920 -960 417144 480
rect 418824 -960 419048 480
rect 420728 -960 420952 480
rect 422632 -960 422856 480
rect 424536 -960 424760 480
rect 426440 -960 426664 480
rect 428344 -960 428568 480
rect 430248 -960 430472 480
rect 432152 -960 432376 480
rect 434056 -960 434280 480
rect 435960 -960 436184 480
rect 437864 -960 438088 480
rect 439768 -960 439992 480
rect 441672 -960 441896 480
rect 443576 -960 443800 480
rect 445480 -960 445704 480
rect 447384 -960 447608 480
rect 449288 -960 449512 480
rect 451192 -960 451416 480
rect 453096 -960 453320 480
rect 455000 -960 455224 480
rect 456904 -960 457128 480
rect 458808 -960 459032 480
rect 460712 -960 460936 480
rect 462616 -960 462840 480
rect 464520 -960 464744 480
rect 466424 -960 466648 480
rect 468328 -960 468552 480
rect 470232 -960 470456 480
rect 472136 -960 472360 480
rect 474040 -960 474264 480
rect 475944 -960 476168 480
rect 477848 -960 478072 480
rect 479752 -960 479976 480
rect 481656 -960 481880 480
rect 483560 -960 483784 480
rect 485464 -960 485688 480
rect 487368 -960 487592 480
rect 489272 -960 489496 480
rect 491176 -960 491400 480
rect 493080 -960 493304 480
rect 494984 -960 495208 480
rect 496888 -960 497112 480
rect 498792 -960 499016 480
rect 500696 -960 500920 480
rect 502600 -960 502824 480
rect 504504 -960 504728 480
rect 506408 -960 506632 480
rect 508312 -960 508536 480
rect 510216 -960 510440 480
rect 512120 -960 512344 480
rect 514024 -960 514248 480
rect 515928 -960 516152 480
rect 517832 -960 518056 480
rect 519736 -960 519960 480
rect 521640 -960 521864 480
rect 523544 -960 523768 480
rect 525448 -960 525672 480
rect 527352 -960 527576 480
rect 529256 -960 529480 480
rect 531160 -960 531384 480
rect 533064 -960 533288 480
rect 534968 -960 535192 480
rect 536872 -960 537096 480
rect 538776 -960 539000 480
rect 540680 -960 540904 480
rect 542584 -960 542808 480
rect 544488 -960 544712 480
rect 546392 -960 546616 480
rect 548296 -960 548520 480
rect 550200 -960 550424 480
rect 552104 -960 552328 480
rect 554008 -960 554232 480
rect 555912 -960 556136 480
rect 557816 -960 558040 480
rect 559720 -960 559944 480
rect 561624 -960 561848 480
rect 563528 -960 563752 480
rect 565432 -960 565656 480
rect 567336 -960 567560 480
rect 569240 -960 569464 480
rect 571144 -960 571368 480
rect 573048 -960 573272 480
rect 574952 -960 575176 480
rect 576856 -960 577080 480
rect 578760 -960 578984 480
rect 580636 392 580888 480
rect 582540 392 582792 480
rect 584444 392 584696 480
rect 580664 -960 580888 392
rect 582568 -960 582792 392
rect 584472 -960 584696 392
<< via2 >>
rect 4172 460124 4228 460180
rect 4172 417788 4228 417844
rect 4172 415772 4228 415828
rect 4284 410732 4340 410788
rect 10892 389900 10948 389956
rect 4172 333116 4228 333172
rect 4172 322476 4228 322532
rect 4172 297500 4228 297556
rect 4172 291004 4228 291060
rect 4172 208684 4228 208740
rect 4172 121660 4228 121716
rect 4172 79100 4228 79156
rect 4172 50316 4228 50372
rect 4396 49644 4452 49700
rect 4396 36876 4452 36932
rect 12572 488348 12628 488404
rect 15932 415772 15988 415828
rect 15932 407820 15988 407876
rect 12572 402668 12628 402724
rect 121548 590604 121604 590660
rect 136892 590604 136948 590660
rect 99484 590492 99540 590548
rect 77308 570332 77364 570388
rect 55132 409836 55188 409892
rect 56252 530684 56308 530740
rect 136892 409724 136948 409780
rect 56252 404124 56308 404180
rect 111692 402556 111748 402612
rect 106652 393372 106708 393428
rect 103292 393260 103348 393316
rect 33068 390572 33124 390628
rect 40908 393148 40964 393204
rect 31052 386764 31108 386820
rect 11004 311612 11060 311668
rect 14252 386652 14308 386708
rect 10892 22876 10948 22932
rect 13244 222684 13300 222740
rect 11564 5852 11620 5908
rect 24668 242620 24724 242676
rect 14252 191996 14308 192052
rect 15148 229292 15204 229348
rect 17052 227612 17108 227668
rect 22764 224364 22820 224420
rect 18956 222572 19012 222628
rect 20860 217532 20916 217588
rect 26572 212492 26628 212548
rect 30380 210812 30436 210868
rect 34412 385420 34468 385476
rect 34412 276668 34468 276724
rect 40236 383852 40292 383908
rect 100156 391580 100212 391636
rect 99932 391468 99988 391524
rect 41132 384076 41188 384132
rect 40908 241948 40964 242004
rect 41020 383964 41076 384020
rect 62412 383068 62468 383124
rect 77420 303212 77476 303268
rect 92428 301532 92484 301588
rect 47404 299292 47460 299348
rect 41580 241948 41636 242004
rect 41468 240492 41524 240548
rect 50764 240716 50820 240772
rect 44156 240492 44212 240548
rect 54796 240492 54852 240548
rect 58828 240380 58884 240436
rect 62860 240268 62916 240324
rect 52780 240156 52836 240212
rect 60844 240156 60900 240212
rect 41020 238476 41076 238532
rect 46732 238476 46788 238532
rect 40236 238252 40292 238308
rect 56812 240044 56868 240100
rect 64876 239708 64932 239764
rect 48748 238252 48804 238308
rect 66892 236796 66948 236852
rect 38556 236012 38612 236068
rect 31052 107324 31108 107380
rect 32284 234444 32340 234500
rect 37996 232764 38052 232820
rect 34188 224252 34244 224308
rect 38444 227724 38500 227780
rect 38444 4844 38500 4900
rect 70924 236572 70980 236628
rect 68908 235116 68964 235172
rect 74956 238476 75012 238532
rect 78988 239820 79044 239876
rect 76972 238476 77028 238532
rect 81004 237804 81060 237860
rect 91084 238476 91140 238532
rect 93100 238364 93156 238420
rect 95116 238364 95172 238420
rect 89068 238140 89124 238196
rect 99820 238588 99876 238644
rect 99932 238476 99988 238532
rect 99820 238252 99876 238308
rect 97132 238140 97188 238196
rect 87052 238028 87108 238084
rect 85036 237916 85092 237972
rect 100156 237692 100212 237748
rect 100380 390012 100436 390068
rect 83020 237580 83076 237636
rect 102508 257068 102564 257124
rect 102508 255276 102564 255332
rect 104972 390124 105028 390180
rect 103404 286412 103460 286468
rect 103516 285292 103572 285348
rect 103516 272748 103572 272804
rect 103404 266924 103460 266980
rect 103292 238252 103348 238308
rect 106652 238140 106708 238196
rect 110012 384300 110068 384356
rect 104972 238028 105028 238084
rect 120092 391804 120148 391860
rect 116732 389228 116788 389284
rect 111692 284396 111748 284452
rect 113372 321692 113428 321748
rect 113372 278572 113428 278628
rect 115052 320012 115108 320068
rect 115052 261100 115108 261156
rect 116732 239708 116788 239764
rect 126812 388220 126868 388276
rect 138572 386316 138628 386372
rect 138572 361340 138628 361396
rect 165452 590492 165508 590548
rect 148652 570332 148708 570388
rect 165676 590156 165732 590212
rect 168812 590156 168868 590212
rect 165452 399196 165508 399252
rect 190540 591164 190596 591220
rect 190316 590716 190372 590772
rect 187740 590156 187796 590212
rect 188972 590156 189028 590212
rect 182252 587132 182308 587188
rect 177212 573020 177268 573076
rect 175532 446012 175588 446068
rect 175532 400652 175588 400708
rect 168812 397740 168868 397796
rect 181356 410732 181412 410788
rect 182252 409612 182308 409668
rect 188972 409500 189028 409556
rect 190316 409052 190372 409108
rect 190428 572012 190484 572068
rect 181356 408044 181412 408100
rect 190540 408268 190596 408324
rect 190652 590940 190708 590996
rect 209580 590380 209636 590436
rect 253708 591276 253764 591332
rect 275772 591164 275828 591220
rect 297836 591052 297892 591108
rect 319900 590940 319956 590996
rect 341964 590828 342020 590884
rect 364028 590716 364084 590772
rect 408268 591276 408324 591332
rect 386092 590604 386148 590660
rect 430220 590492 430276 590548
rect 474348 591276 474404 591332
rect 496636 590604 496692 590660
rect 452508 590492 452564 590548
rect 231644 572012 231700 572068
rect 560252 591276 560308 591332
rect 540764 590716 540820 590772
rect 549836 590716 549892 590772
rect 518476 570332 518532 570388
rect 549388 550396 549444 550452
rect 548492 410508 548548 410564
rect 190652 407932 190708 407988
rect 195132 406588 195188 406644
rect 197372 408268 197428 408324
rect 190428 393932 190484 393988
rect 177212 390684 177268 390740
rect 196588 346892 196644 346948
rect 181356 313292 181412 313348
rect 148652 288988 148708 289044
rect 163772 297388 163828 297444
rect 163772 290556 163828 290612
rect 143388 287868 143444 287924
rect 172844 289884 172900 289940
rect 192332 288988 192388 289044
rect 196700 343532 196756 343588
rect 198268 406588 198324 406644
rect 198380 336812 198436 336868
rect 196700 286412 196756 286468
rect 197484 285628 197540 285684
rect 196588 285292 196644 285348
rect 197372 284732 197428 284788
rect 192332 253596 192388 253652
rect 196476 257068 196532 257124
rect 198380 284732 198436 284788
rect 199164 339164 199220 339220
rect 198492 329420 198548 329476
rect 197372 257068 197428 257124
rect 196476 245868 196532 245924
rect 199052 333452 199108 333508
rect 204092 391916 204148 391972
rect 200508 333452 200564 333508
rect 202412 368732 202468 368788
rect 199164 320012 199220 320068
rect 200732 331548 200788 331604
rect 199052 249564 199108 249620
rect 198492 243628 198548 243684
rect 126812 240716 126868 240772
rect 120092 237916 120148 237972
rect 110012 237804 110068 237860
rect 100380 237580 100436 237636
rect 72940 235004 72996 235060
rect 41020 232652 41076 232708
rect 40236 229404 40292 229460
rect 40124 217644 40180 217700
rect 40124 4284 40180 4340
rect 38556 4172 38612 4228
rect 39900 4172 39956 4228
rect 40236 4172 40292 4228
rect 41132 230972 41188 231028
rect 199052 215852 199108 215908
rect 154924 214172 154980 214228
rect 202412 289884 202468 289940
rect 205772 388444 205828 388500
rect 210812 388668 210868 388724
rect 205884 336812 205940 336868
rect 207452 384188 207508 384244
rect 205772 239932 205828 239988
rect 204092 238476 204148 238532
rect 215852 388780 215908 388836
rect 211260 339164 211316 339220
rect 212492 386204 212548 386260
rect 212492 319004 212548 319060
rect 214172 370748 214228 370804
rect 214172 313292 214228 313348
rect 222572 403228 222628 403284
rect 219212 389116 219268 389172
rect 217532 388892 217588 388948
rect 215964 383180 216020 383236
rect 215964 343532 216020 343588
rect 215964 311612 216020 311668
rect 215964 290108 216020 290164
rect 215852 240380 215908 240436
rect 217532 240156 217588 240212
rect 217756 388556 217812 388612
rect 210812 240044 210868 240100
rect 227612 406588 227668 406644
rect 223244 368508 223300 368564
rect 222572 346892 222628 346948
rect 223132 361788 223188 361844
rect 219212 240268 219268 240324
rect 219996 343868 220052 343924
rect 217756 239820 217812 239876
rect 223020 339388 223076 339444
rect 226716 367388 226772 367444
rect 225036 365148 225092 365204
rect 223244 251132 223300 251188
rect 223356 364028 223412 364084
rect 223132 249452 223188 249508
rect 223020 241500 223076 241556
rect 224924 341628 224980 341684
rect 224924 248108 224980 248164
rect 226492 359548 226548 359604
rect 226380 357308 226436 357364
rect 225036 247772 225092 247828
rect 226268 344988 226324 345044
rect 226492 251244 226548 251300
rect 226604 355068 226660 355124
rect 226380 247884 226436 247940
rect 226268 244412 226324 244468
rect 227948 407932 228004 407988
rect 227836 350588 227892 350644
rect 227612 323372 227668 323428
rect 227724 326060 227780 326116
rect 227500 306908 227556 306964
rect 227612 297500 227668 297556
rect 227612 251692 227668 251748
rect 227500 246316 227556 246372
rect 226716 242732 226772 242788
rect 226604 241276 226660 241332
rect 223356 241164 223412 241220
rect 230188 407484 230244 407540
rect 230188 406476 230244 406532
rect 232764 406700 232820 406756
rect 228508 404460 228564 404516
rect 228508 404012 228564 404068
rect 229516 404460 229572 404516
rect 229404 393484 229460 393540
rect 229292 392028 229348 392084
rect 228396 362908 228452 362964
rect 228284 358428 228340 358484
rect 228172 352828 228228 352884
rect 227948 303996 228004 304052
rect 227948 303212 228004 303268
rect 228060 349468 228116 349524
rect 227836 251356 227892 251412
rect 228172 242956 228228 243012
rect 228396 246092 228452 246148
rect 228284 242844 228340 242900
rect 228060 241388 228116 241444
rect 227724 239932 227780 239988
rect 219996 237692 220052 237748
rect 231196 404348 231252 404404
rect 230076 353948 230132 354004
rect 229852 348348 229908 348404
rect 229740 340508 229796 340564
rect 229516 301532 229572 301588
rect 229516 300748 229572 300804
rect 229628 303996 229684 304052
rect 229404 236572 229460 236628
rect 229292 235004 229348 235060
rect 207452 234332 207508 234388
rect 229852 249788 229908 249844
rect 229964 339500 230020 339556
rect 229740 246204 229796 246260
rect 237692 407932 237748 407988
rect 238140 407708 238196 407764
rect 243516 407596 243572 407652
rect 252588 409388 252644 409444
rect 248892 406812 248948 406868
rect 251692 409164 251748 409220
rect 237692 404572 237748 404628
rect 232764 402556 232820 402612
rect 231644 400764 231700 400820
rect 231532 347228 231588 347284
rect 231420 337148 231476 337204
rect 231196 322476 231252 322532
rect 231308 336028 231364 336084
rect 230972 300748 231028 300804
rect 231084 276332 231140 276388
rect 231084 254940 231140 254996
rect 231308 251468 231364 251524
rect 230972 250012 231028 250068
rect 231420 244524 231476 244580
rect 230188 243180 230244 243236
rect 233324 397404 233380 397460
rect 231644 243180 231700 243236
rect 231756 394044 231812 394100
rect 231532 243068 231588 243124
rect 230188 242508 230244 242564
rect 230076 239820 230132 239876
rect 229964 239708 230020 239764
rect 233212 369628 233268 369684
rect 233212 368732 233268 368788
rect 233212 366268 233268 366324
rect 232652 360668 232708 360724
rect 232652 339500 232708 339556
rect 232764 342748 232820 342804
rect 233212 331772 233268 331828
rect 232764 326060 232820 326116
rect 231868 322476 231924 322532
rect 233212 309148 233268 309204
rect 233100 308028 233156 308084
rect 233100 257292 233156 257348
rect 249900 405692 249956 405748
rect 247212 404012 247268 404068
rect 246316 399084 246372 399140
rect 236012 392252 236068 392308
rect 235004 387324 235060 387380
rect 234556 386092 234612 386148
rect 234332 385980 234388 386036
rect 233324 281148 233380 281204
rect 233436 384524 233492 384580
rect 233212 256060 233268 256116
rect 233324 264348 233380 264404
rect 233324 254492 233380 254548
rect 231868 246876 231924 246932
rect 231756 216412 231812 216468
rect 229628 216188 229684 216244
rect 200732 214172 200788 214228
rect 234220 281372 234276 281428
rect 234220 254828 234276 254884
rect 234444 331772 234500 331828
rect 234444 239596 234500 239652
rect 234892 351708 234948 351764
rect 234780 334908 234836 334964
rect 234668 283948 234724 284004
rect 234668 256396 234724 256452
rect 234780 251580 234836 251636
rect 234892 247996 234948 248052
rect 234556 236796 234612 236852
rect 234332 235116 234388 235172
rect 235004 216076 235060 216132
rect 235116 385756 235172 385812
rect 235676 385644 235732 385700
rect 235788 385532 235844 385588
rect 235116 213276 235172 213332
rect 235676 384412 235732 384468
rect 233436 213052 233492 213108
rect 235788 212828 235844 212884
rect 235676 212716 235732 212772
rect 242732 390348 242788 390404
rect 240940 390236 240996 390292
rect 240044 389788 240100 389844
rect 238252 388108 238308 388164
rect 237356 386988 237412 387044
rect 239148 386428 239204 386484
rect 241836 386540 241892 386596
rect 243628 387100 243684 387156
rect 245420 390460 245476 390516
rect 248108 402556 248164 402612
rect 249004 397516 249060 397572
rect 250796 397628 250852 397684
rect 253484 409052 253540 409108
rect 254268 407372 254324 407428
rect 254380 409276 254436 409332
rect 270396 407932 270452 407988
rect 273756 409052 273812 409108
rect 273756 407596 273812 407652
rect 280588 409500 280644 409556
rect 265020 407484 265076 407540
rect 260428 406812 260484 406868
rect 259756 404124 259812 404180
rect 257068 399196 257124 399252
rect 256172 397740 256228 397796
rect 255276 393932 255332 393988
rect 258860 390684 258916 390740
rect 257964 390572 258020 390628
rect 275436 404460 275492 404516
rect 262444 403676 262500 403732
rect 260428 394044 260484 394100
rect 260652 402668 260708 402724
rect 261548 400652 261604 400708
rect 270508 389900 270564 389956
rect 268716 386764 268772 386820
rect 266924 386652 266980 386708
rect 263340 386316 263396 386372
rect 264236 386204 264292 386260
rect 272300 389900 272356 389956
rect 277676 388332 277732 388388
rect 274092 387324 274148 387380
rect 278572 386764 278628 386820
rect 280364 386316 280420 386372
rect 279468 386204 279524 386260
rect 286524 409724 286580 409780
rect 290668 409836 290724 409892
rect 286300 406924 286356 406980
rect 291900 409836 291956 409892
rect 295708 409612 295764 409668
rect 290668 392476 290724 392532
rect 292012 393148 292068 393204
rect 280588 385868 280644 385924
rect 282156 388108 282212 388164
rect 283948 386652 284004 386708
rect 297276 409612 297332 409668
rect 308028 409276 308084 409332
rect 302652 408828 302708 408884
rect 302652 406924 302708 406980
rect 295708 392364 295764 392420
rect 304556 393484 304612 393540
rect 301868 389228 301924 389284
rect 300972 389116 301028 389172
rect 300076 388892 300132 388948
rect 299180 388780 299236 388836
rect 296492 388668 296548 388724
rect 295596 388220 295652 388276
rect 298284 388444 298340 388500
rect 297388 388108 297444 388164
rect 302764 386092 302820 386148
rect 302988 385980 303044 386036
rect 305452 392028 305508 392084
rect 307244 391692 307300 391748
rect 306348 386876 306404 386932
rect 308140 388556 308196 388612
rect 313292 408044 313348 408100
rect 310828 391804 310884 391860
rect 308812 385980 308868 386036
rect 309932 390012 309988 390068
rect 312620 391580 312676 391636
rect 311724 390124 311780 390180
rect 318332 407820 318388 407876
rect 317996 397740 318052 397796
rect 316204 393372 316260 393428
rect 315308 393260 315364 393316
rect 314412 391916 314468 391972
rect 313292 385980 313348 386036
rect 313516 391468 313572 391524
rect 317100 388892 317156 388948
rect 322476 402220 322532 402276
rect 319788 400652 319844 400708
rect 318332 386092 318388 386148
rect 318892 392364 318948 392420
rect 321580 395724 321636 395780
rect 320684 392140 320740 392196
rect 323372 395612 323428 395668
rect 322588 393148 322644 393204
rect 322588 392252 322644 392308
rect 328748 409276 328804 409332
rect 324156 393148 324212 393204
rect 324268 406252 324324 406308
rect 327852 404684 327908 404740
rect 326732 401100 326788 401156
rect 326060 393036 326116 393092
rect 325164 389004 325220 389060
rect 326732 388892 326788 388948
rect 326956 389228 327012 389284
rect 333452 409500 333508 409556
rect 329532 404348 329588 404404
rect 332332 409388 332388 409444
rect 331436 400988 331492 401044
rect 330876 395836 330932 395892
rect 329644 392252 329700 392308
rect 330540 389676 330596 389732
rect 330876 389004 330932 389060
rect 333228 390796 333284 390852
rect 334908 400876 334964 400932
rect 338604 404572 338660 404628
rect 336812 399644 336868 399700
rect 335916 399196 335972 399252
rect 333452 389676 333508 389732
rect 335020 394716 335076 394772
rect 334124 388892 334180 388948
rect 337708 393932 337764 393988
rect 351036 407708 351092 407764
rect 355628 409612 355684 409668
rect 345660 407596 345716 407652
rect 351148 406140 351204 406196
rect 349356 404460 349412 404516
rect 340284 400764 340340 400820
rect 340396 403116 340452 403172
rect 339500 394044 339556 394100
rect 348460 402668 348516 402724
rect 342188 400876 342244 400932
rect 341292 394156 341348 394212
rect 345772 399532 345828 399588
rect 343980 398076 344036 398132
rect 343084 394268 343140 394324
rect 344876 394492 344932 394548
rect 346668 394380 346724 394436
rect 347564 389116 347620 389172
rect 350252 395948 350308 396004
rect 353836 404124 353892 404180
rect 352940 403004 352996 403060
rect 352044 396060 352100 396116
rect 354732 392924 354788 392980
rect 356412 407820 356468 407876
rect 360332 407484 360388 407540
rect 359212 405804 359268 405860
rect 358316 392812 358372 392868
rect 356524 392700 356580 392756
rect 357420 390572 357476 390628
rect 360108 392588 360164 392644
rect 361788 404796 361844 404852
rect 362796 409724 362852 409780
rect 360332 392252 360388 392308
rect 361004 394604 361060 394660
rect 361900 392476 361956 392532
rect 365372 407932 365428 407988
rect 363692 400764 363748 400820
rect 367164 401436 367220 401492
rect 368732 409836 368788 409892
rect 367276 399420 367332 399476
rect 365372 392364 365428 392420
rect 365484 397964 365540 398020
rect 364588 392252 364644 392308
rect 366380 389676 366436 389732
rect 368732 389676 368788 389732
rect 369068 404348 369124 404404
rect 368172 389004 368228 389060
rect 370860 402892 370916 402948
rect 369964 395500 370020 395556
rect 377916 407932 377972 407988
rect 375676 407820 375732 407876
rect 375564 407708 375620 407764
rect 372540 401100 372596 401156
rect 374444 406028 374500 406084
rect 372652 392364 372708 392420
rect 371308 390908 371364 390964
rect 371308 389116 371364 389172
rect 371756 389340 371812 389396
rect 373548 389116 373604 389172
rect 375340 388108 375396 388164
rect 243852 385756 243908 385812
rect 244524 385756 244580 385812
rect 274988 385644 275044 385700
rect 284844 385644 284900 385700
rect 276780 385532 276836 385588
rect 286636 385532 286692 385588
rect 265132 385420 265188 385476
rect 267820 385420 267876 385476
rect 273196 385420 273252 385476
rect 285740 385420 285796 385476
rect 236124 385308 236180 385364
rect 266028 385308 266084 385364
rect 269612 385308 269668 385364
rect 271404 385308 271460 385364
rect 275884 385308 275940 385364
rect 281260 385308 281316 385364
rect 283052 385308 283108 385364
rect 287532 385308 287588 385364
rect 288428 385308 288484 385364
rect 289324 385308 289380 385364
rect 290220 385308 290276 385364
rect 291116 385308 291172 385364
rect 292908 385308 292964 385364
rect 293804 385308 293860 385364
rect 294700 385308 294756 385364
rect 309036 385308 309092 385364
rect 236012 375452 236068 375508
rect 236012 355964 236068 356020
rect 236012 249676 236068 249732
rect 236124 345884 236180 345940
rect 236236 337932 236292 337988
rect 242732 253596 242788 253652
rect 236236 249900 236292 249956
rect 236124 248220 236180 248276
rect 244524 224364 244580 224420
rect 242956 222684 243012 222740
rect 235900 212604 235956 212660
rect 246316 232764 246372 232820
rect 247212 227724 247268 227780
rect 249004 231084 249060 231140
rect 248108 217644 248164 217700
rect 251916 253596 251972 253652
rect 252588 253596 252644 253652
rect 253484 249340 253540 249396
rect 256172 250124 256228 250180
rect 255276 246540 255332 246596
rect 254380 246428 254436 246484
rect 257068 245980 257124 246036
rect 258860 253596 258916 253652
rect 259756 253596 259812 253652
rect 260652 253596 260708 253652
rect 261548 252924 261604 252980
rect 264236 253260 264292 253316
rect 266028 253484 266084 253540
rect 265132 253148 265188 253204
rect 263340 253036 263396 253092
rect 262444 252812 262500 252868
rect 267820 252252 267876 252308
rect 268716 252140 268772 252196
rect 266924 252028 266980 252084
rect 257964 243292 258020 243348
rect 250796 229404 250852 229460
rect 249900 215964 249956 216020
rect 269388 216412 269444 216468
rect 245420 210812 245476 210868
rect 269276 213276 269332 213332
rect 269500 211148 269556 211204
rect 269500 210700 269556 210756
rect 269500 209692 269556 209748
rect 269500 204652 269556 204708
rect 269388 88172 269444 88228
rect 269500 142828 269556 142884
rect 269276 79212 269332 79268
rect 269500 50316 269556 50372
rect 91308 49532 91364 49588
rect 47852 48636 47908 48692
rect 47516 15932 47572 15988
rect 41132 4396 41188 4452
rect 45612 4844 45668 4900
rect 87500 47852 87556 47908
rect 68460 41132 68516 41188
rect 57148 37772 57204 37828
rect 47852 5852 47908 5908
rect 55132 17612 55188 17668
rect 49420 4396 49476 4452
rect 53228 4284 53284 4340
rect 62748 34412 62804 34468
rect 60844 19292 60900 19348
rect 58940 4508 58996 4564
rect 66780 4620 66836 4676
rect 64652 4396 64708 4452
rect 76076 36092 76132 36148
rect 74172 34524 74228 34580
rect 72268 24332 72324 24388
rect 68908 9324 68964 9380
rect 68908 4620 68964 4676
rect 70364 4172 70420 4228
rect 81788 34636 81844 34692
rect 79884 31052 79940 31108
rect 77980 14252 78036 14308
rect 83692 29372 83748 29428
rect 85820 4284 85876 4340
rect 89404 32844 89460 32900
rect 180796 49868 180852 49924
rect 97356 48636 97412 48692
rect 167468 49756 167524 49812
rect 127484 48076 127540 48132
rect 93212 47964 93268 48020
rect 110348 44940 110404 44996
rect 104636 44828 104692 44884
rect 98924 44716 98980 44772
rect 97020 41244 97076 41300
rect 95116 19404 95172 19460
rect 102732 32732 102788 32788
rect 101052 5852 101108 5908
rect 108444 37884 108500 37940
rect 106764 7532 106820 7588
rect 116060 41468 116116 41524
rect 112476 7644 112532 7700
rect 114380 4172 114436 4228
rect 119868 37996 119924 38052
rect 118188 7756 118244 7812
rect 121772 34860 121828 34916
rect 123676 17724 123732 17780
rect 125804 4844 125860 4900
rect 138908 45052 138964 45108
rect 133196 32956 133252 33012
rect 129388 16044 129444 16100
rect 131516 9212 131572 9268
rect 135100 24444 135156 24500
rect 137228 4060 137284 4116
rect 148428 44604 148484 44660
rect 142828 44492 142884 44548
rect 140812 14364 140868 14420
rect 144620 31276 144676 31332
rect 146524 26012 146580 26068
rect 156044 42924 156100 42980
rect 152236 31164 152292 31220
rect 150556 10892 150612 10948
rect 154364 4396 154420 4452
rect 159852 41356 159908 41412
rect 158172 5964 158228 6020
rect 161756 39452 161812 39508
rect 163660 12572 163716 12628
rect 165788 4508 165844 4564
rect 178892 48188 178948 48244
rect 175084 41580 175140 41636
rect 171388 38108 171444 38164
rect 169372 29484 169428 29540
rect 173180 26124 173236 26180
rect 177212 4620 177268 4676
rect 212268 48524 212324 48580
rect 197932 48300 197988 48356
rect 184604 46172 184660 46228
rect 182700 38220 182756 38276
rect 188412 42812 188468 42868
rect 186508 20972 186564 21028
rect 192220 38332 192276 38388
rect 190540 6076 190596 6132
rect 194124 34748 194180 34804
rect 196028 24556 196084 24612
rect 207452 45164 207508 45220
rect 203644 41692 203700 41748
rect 201740 14476 201796 14532
rect 200060 4732 200116 4788
rect 205772 4956 205828 5012
rect 209356 36204 209412 36260
rect 211260 34972 211316 35028
rect 269724 252028 269780 252084
rect 269836 211372 269892 211428
rect 269836 207900 269892 207956
rect 269724 26124 269780 26180
rect 270620 250124 270676 250180
rect 270844 246540 270900 246596
rect 270620 44828 270676 44884
rect 270732 243292 270788 243348
rect 271068 246428 271124 246484
rect 270956 245980 271012 246036
rect 271180 145292 271236 145348
rect 271180 49644 271236 49700
rect 271068 47964 271124 48020
rect 270956 44940 271012 44996
rect 270844 44716 270900 44772
rect 270732 41468 270788 41524
rect 270508 24556 270564 24612
rect 272300 252028 272356 252084
rect 272188 251692 272244 251748
rect 272972 245308 273028 245364
rect 272748 210140 272804 210196
rect 272524 210028 272580 210084
rect 272412 209804 272468 209860
rect 272188 154028 272244 154084
rect 272300 208684 272356 208740
rect 272412 180796 272468 180852
rect 272300 140700 272356 140756
rect 272524 153468 272580 153524
rect 272524 137116 272580 137172
rect 272748 154364 272804 154420
rect 272748 134204 272804 134260
rect 273868 255836 273924 255892
rect 273196 242620 273252 242676
rect 273420 243180 273476 243236
rect 272972 153020 273028 153076
rect 272972 125468 273028 125524
rect 273084 216188 273140 216244
rect 271404 14476 271460 14532
rect 272972 120092 273028 120148
rect 269612 6076 269668 6132
rect 273308 155372 273364 155428
rect 273084 109116 273140 109172
rect 273084 93436 273140 93492
rect 273196 154364 273252 154420
rect 273420 153132 273476 153188
rect 273420 131292 273476 131348
rect 273644 154476 273700 154532
rect 273308 96348 273364 96404
rect 273980 250012 274036 250068
rect 275660 253484 275716 253540
rect 274988 236012 275044 236068
rect 275548 253260 275604 253316
rect 274092 234444 274148 234500
rect 274876 213052 274932 213108
rect 273980 155372 274036 155428
rect 274652 211484 274708 211540
rect 273868 151676 273924 151732
rect 275324 156380 275380 156436
rect 275436 156268 275492 156324
rect 275436 154476 275492 154532
rect 275324 154364 275380 154420
rect 274652 152796 274708 152852
rect 273756 136108 273812 136164
rect 273756 128380 273812 128436
rect 273644 90524 273700 90580
rect 274652 123452 274708 123508
rect 273196 81788 273252 81844
rect 273084 73052 273140 73108
rect 273308 70140 273364 70196
rect 273084 52780 273140 52836
rect 273196 67228 273252 67284
rect 273308 52668 273364 52724
rect 273196 50652 273252 50708
rect 272972 4844 273028 4900
rect 274764 99260 274820 99316
rect 274876 121772 274932 121828
rect 274652 4284 274708 4340
rect 275660 49756 275716 49812
rect 275548 42924 275604 42980
rect 276332 152124 276388 152180
rect 276332 75964 276388 76020
rect 276332 58492 276388 58548
rect 276332 50540 276388 50596
rect 276780 17612 276836 17668
rect 277228 253036 277284 253092
rect 275884 15932 275940 15988
rect 277340 252924 277396 252980
rect 277564 252252 277620 252308
rect 277452 252140 277508 252196
rect 277564 48188 277620 48244
rect 277452 46172 277508 46228
rect 277340 45052 277396 45108
rect 278012 61404 278068 61460
rect 278012 50316 278068 50372
rect 277676 19292 277732 19348
rect 277228 10892 277284 10948
rect 279020 253148 279076 253204
rect 278908 252812 278964 252868
rect 279132 252028 279188 252084
rect 279132 45164 279188 45220
rect 279020 39452 279076 39508
rect 278908 31276 278964 31332
rect 279468 24332 279524 24388
rect 281372 252812 281428 252868
rect 281372 48300 281428 48356
rect 282156 32844 282212 32900
rect 281260 29372 281316 29428
rect 283388 252924 283444 252980
rect 283164 252476 283220 252532
rect 283836 156492 283892 156548
rect 283836 152908 283892 152964
rect 283388 41692 283444 41748
rect 283164 26012 283220 26068
rect 283052 19404 283108 19460
rect 280364 14252 280420 14308
rect 278572 9324 278628 9380
rect 284732 253036 284788 253092
rect 284732 36204 284788 36260
rect 284956 253148 285012 253204
rect 284956 41580 285012 41636
rect 286412 210924 286468 210980
rect 286412 154476 286468 154532
rect 286412 102172 286468 102228
rect 288316 253260 288372 253316
rect 288092 252028 288148 252084
rect 287980 55580 288036 55636
rect 287980 50428 288036 50484
rect 288316 49868 288372 49924
rect 288092 24444 288148 24500
rect 287532 17724 287588 17780
rect 289324 252028 289380 252084
rect 289772 252700 289828 252756
rect 289996 252252 290052 252308
rect 289884 216076 289940 216132
rect 289884 48524 289940 48580
rect 290108 64316 290164 64372
rect 290108 51772 290164 51828
rect 289996 31164 290052 31220
rect 289772 29484 289828 29540
rect 288428 16044 288484 16100
rect 290332 253372 290388 253428
rect 291116 252476 291172 252532
rect 292012 252364 292068 252420
rect 290332 38332 290388 38388
rect 290892 252252 290948 252308
rect 290892 20972 290948 21028
rect 291116 252140 291172 252196
rect 290220 14364 290276 14420
rect 296492 253260 296548 253316
rect 295596 253148 295652 253204
rect 294700 252700 294756 252756
rect 298284 253372 298340 253428
rect 300972 253036 301028 253092
rect 300076 252924 300132 252980
rect 299180 252812 299236 252868
rect 297388 252252 297444 252308
rect 293804 252140 293860 252196
rect 301868 252140 301924 252196
rect 292908 252028 292964 252084
rect 295148 154700 295204 154756
rect 295148 154252 295204 154308
rect 293132 150332 293188 150388
rect 302764 125356 302820 125412
rect 304556 252028 304612 252084
rect 304892 252140 304948 252196
rect 303996 152908 304052 152964
rect 303996 150332 304052 150388
rect 306348 217756 306404 217812
rect 305452 197372 305508 197428
rect 304892 133532 304948 133588
rect 307356 160636 307412 160692
rect 307356 152908 307412 152964
rect 307244 126924 307300 126980
rect 309036 231196 309092 231252
rect 310828 252812 310884 252868
rect 309932 192332 309988 192388
rect 310044 252028 310100 252084
rect 308140 126812 308196 126868
rect 308252 154476 308308 154532
rect 303660 125244 303716 125300
rect 308252 113820 308308 113876
rect 309932 151340 309988 151396
rect 293132 110908 293188 110964
rect 310940 160748 310996 160804
rect 310940 154476 310996 154532
rect 310044 150556 310100 150612
rect 312620 252924 312676 252980
rect 313516 252028 313572 252084
rect 314972 252028 315028 252084
rect 314972 234444 315028 234500
rect 314412 204092 314468 204148
rect 317100 252140 317156 252196
rect 316204 252028 316260 252084
rect 315308 138572 315364 138628
rect 311724 131852 311780 131908
rect 318332 252028 318388 252084
rect 319788 252364 319844 252420
rect 320012 252924 320068 252980
rect 318892 252028 318948 252084
rect 318332 232876 318388 232932
rect 317996 125132 318052 125188
rect 318332 153692 318388 153748
rect 320236 252140 320292 252196
rect 320236 231084 320292 231140
rect 321580 252252 321636 252308
rect 321692 252812 321748 252868
rect 320684 227724 320740 227780
rect 320012 141932 320068 141988
rect 321916 252028 321972 252084
rect 322476 234332 322532 234388
rect 323484 252364 323540 252420
rect 323484 229404 323540 229460
rect 323372 222684 323428 222740
rect 325164 252140 325220 252196
rect 325388 252252 325444 252308
rect 326060 252028 326116 252084
rect 326732 254492 326788 254548
rect 325388 224364 325444 224420
rect 324268 217644 324324 217700
rect 325052 217756 325108 217812
rect 321916 205772 321972 205828
rect 321692 128492 321748 128548
rect 323372 153804 323428 153860
rect 325052 123676 325108 123732
rect 323372 122556 323428 122612
rect 318332 119644 318388 119700
rect 309932 84700 309988 84756
rect 307468 50204 307524 50260
rect 314188 50204 314244 50260
rect 321356 50204 321412 50260
rect 293580 50092 293636 50148
rect 293580 48636 293636 48692
rect 300748 48524 300804 48580
rect 326844 252140 326900 252196
rect 326844 232764 326900 232820
rect 326956 194124 327012 194180
rect 327852 182364 327908 182420
rect 328412 254492 328468 254548
rect 326732 33628 326788 33684
rect 291116 12572 291172 12628
rect 286636 7756 286692 7812
rect 285740 7644 285796 7700
rect 284844 7532 284900 7588
rect 283948 5852 284004 5908
rect 328748 170604 328804 170660
rect 329644 158956 329700 159012
rect 330092 254604 330148 254660
rect 330540 199164 330596 199220
rect 331436 188972 331492 189028
rect 331772 255948 331828 256004
rect 331884 252028 331940 252084
rect 332332 252028 332388 252084
rect 331884 210812 331940 210868
rect 331884 192332 331940 192388
rect 333452 252028 333508 252084
rect 334124 252028 334180 252084
rect 333452 162204 333508 162260
rect 333228 158844 333284 158900
rect 335132 252028 335188 252084
rect 335916 192444 335972 192500
rect 336812 254380 336868 254436
rect 335132 179004 335188 179060
rect 335020 158732 335076 158788
rect 331884 123564 331940 123620
rect 331772 4620 331828 4676
rect 330092 4508 330148 4564
rect 336924 155708 336980 155764
rect 337708 155596 337764 155652
rect 339500 187404 339556 187460
rect 341292 185612 341348 185668
rect 343084 252028 343140 252084
rect 343980 236796 344036 236852
rect 345212 252028 345268 252084
rect 345212 200508 345268 200564
rect 344876 199052 344932 199108
rect 345772 180572 345828 180628
rect 342188 168812 342244 168868
rect 340396 163884 340452 163940
rect 346668 157276 346724 157332
rect 347564 157164 347620 157220
rect 349356 195692 349412 195748
rect 350252 177212 350308 177268
rect 350476 255948 350532 256004
rect 348460 157052 348516 157108
rect 338604 155484 338660 155540
rect 351148 175532 351204 175588
rect 352940 194012 352996 194068
rect 353836 192332 353892 192388
rect 354732 187292 354788 187348
rect 355292 253260 355348 253316
rect 352044 173852 352100 173908
rect 355628 252028 355684 252084
rect 355740 248444 355796 248500
rect 355516 248332 355572 248388
rect 355292 38220 355348 38276
rect 355404 244636 355460 244692
rect 356972 252028 357028 252084
rect 356972 200620 357028 200676
rect 357420 163772 357476 163828
rect 358316 162092 358372 162148
rect 358652 253372 358708 253428
rect 356524 160524 356580 160580
rect 356972 154252 357028 154308
rect 356972 141036 357028 141092
rect 357756 151452 357812 151508
rect 357644 120204 357700 120260
rect 357756 108892 357812 108948
rect 357644 84924 357700 84980
rect 357756 61628 357812 61684
rect 356188 51884 356244 51940
rect 357756 51884 357812 51940
rect 356188 50092 356244 50148
rect 355740 34972 355796 35028
rect 358988 251804 359044 251860
rect 358764 251692 358820 251748
rect 358764 44492 358820 44548
rect 358988 37996 359044 38052
rect 359212 251020 359268 251076
rect 359324 182252 359380 182308
rect 361004 252812 361060 252868
rect 361900 252140 361956 252196
rect 360108 160412 360164 160468
rect 360332 248556 360388 248612
rect 359212 37884 359268 37940
rect 358652 34748 358708 34804
rect 355516 34524 355572 34580
rect 360556 247660 360612 247716
rect 364588 253036 364644 253092
rect 363692 252028 363748 252084
rect 362796 167132 362852 167188
rect 362012 153580 362068 153636
rect 367276 253148 367332 253204
rect 366380 252252 366436 252308
rect 365484 150332 365540 150388
rect 367052 154476 367108 154532
rect 369068 252924 369124 252980
rect 370412 252140 370468 252196
rect 372092 252028 372148 252084
rect 370412 170492 370468 170548
rect 370748 197372 370804 197428
rect 368172 150444 368228 150500
rect 368732 150556 368788 150612
rect 367052 145292 367108 145348
rect 362012 142940 362068 142996
rect 362684 133532 362740 133588
rect 364700 125356 364756 125412
rect 366716 125244 366772 125300
rect 372092 168924 372148 168980
rect 375452 231196 375508 231252
rect 374780 126924 374836 126980
rect 372764 123676 372820 123732
rect 375676 154252 375732 154308
rect 375788 404796 375844 404852
rect 375900 401436 375956 401492
rect 394044 406252 394100 406308
rect 388668 402220 388724 402276
rect 410172 407484 410228 407540
rect 410732 407484 410788 407540
rect 404796 404684 404852 404740
rect 415548 400988 415604 401044
rect 410732 394716 410788 394772
rect 399420 393036 399476 393092
rect 383292 392140 383348 392196
rect 409276 391132 409332 391188
rect 426300 407484 426356 407540
rect 437052 404572 437108 404628
rect 442428 403116 442484 403172
rect 451948 407484 452004 407540
rect 451948 406812 452004 406868
rect 447804 400876 447860 400932
rect 431676 399644 431732 399700
rect 453180 398076 453236 398132
rect 453516 407484 453572 407540
rect 420924 391132 420980 391188
rect 409276 390908 409332 390964
rect 421596 390796 421652 390852
rect 379820 390684 379876 390740
rect 377132 390460 377188 390516
rect 376348 383068 376404 383124
rect 376348 381276 376404 381332
rect 377132 377132 377188 377188
rect 377244 388332 377300 388388
rect 377132 297276 377188 297332
rect 376572 296156 376628 296212
rect 376348 275996 376404 276052
rect 376012 252028 376068 252084
rect 376348 251804 376404 251860
rect 376460 273756 376516 273812
rect 376460 251020 376516 251076
rect 376684 293916 376740 293972
rect 376796 290556 376852 290612
rect 377020 280476 377076 280532
rect 376796 253372 376852 253428
rect 376908 260316 376964 260372
rect 376684 248444 376740 248500
rect 376572 227612 376628 227668
rect 377020 251692 377076 251748
rect 376908 224252 376964 224308
rect 377132 222572 377188 222628
rect 376012 175644 376068 175700
rect 375900 154476 375956 154532
rect 376124 154364 376180 154420
rect 375564 153468 375620 153524
rect 376012 153804 376068 153860
rect 376236 154252 376292 154308
rect 376236 153692 376292 153748
rect 376124 153580 376180 153636
rect 376012 153468 376068 153524
rect 375452 122668 375508 122724
rect 376796 126812 376852 126868
rect 382172 390348 382228 390404
rect 379820 388108 379876 388164
rect 380492 390236 380548 390292
rect 379036 311836 379092 311892
rect 378924 310716 378980 310772
rect 378812 307356 378868 307412
rect 378364 292796 378420 292852
rect 378252 284956 378308 285012
rect 378028 282716 378084 282772
rect 378140 274876 378196 274932
rect 378476 291676 378532 291732
rect 378476 257292 378532 257348
rect 378588 287196 378644 287252
rect 378588 256172 378644 256228
rect 378700 279356 378756 279412
rect 378364 256060 378420 256116
rect 378252 254604 378308 254660
rect 378140 254492 378196 254548
rect 378028 254380 378084 254436
rect 379036 284508 379092 284564
rect 379708 295036 379764 295092
rect 378924 282156 378980 282212
rect 378812 275548 378868 275604
rect 378924 277116 378980 277172
rect 378700 121772 378756 121828
rect 378812 122668 378868 122724
rect 377244 120204 377300 120260
rect 379036 269276 379092 269332
rect 379820 284508 379876 284564
rect 379820 283948 379876 284004
rect 379820 256396 379876 256452
rect 379932 282156 379988 282212
rect 379932 280588 379988 280644
rect 380044 275548 380100 275604
rect 380044 254940 380100 254996
rect 379932 254828 379988 254884
rect 379708 217532 379764 217588
rect 380604 385756 380660 385812
rect 380604 337484 380660 337540
rect 381388 268156 381444 268212
rect 421596 389340 421652 389396
rect 429212 389900 429268 389956
rect 383852 387100 383908 387156
rect 424172 386988 424228 387044
rect 383852 297836 383908 297892
rect 385532 386764 385588 386820
rect 382172 258188 382228 258244
rect 381388 244636 381444 244692
rect 387212 386316 387268 386372
rect 397292 386204 397348 386260
rect 387212 197260 387268 197316
rect 388892 234444 388948 234500
rect 385532 197148 385588 197204
rect 380492 178892 380548 178948
rect 386876 141932 386932 141988
rect 384860 131852 384916 131908
rect 382844 128492 382900 128548
rect 379036 123452 379092 123508
rect 380828 123564 380884 123620
rect 378924 120092 378980 120148
rect 394940 232876 394996 232932
rect 390908 204092 390964 204148
rect 392924 138572 392980 138628
rect 396956 231084 397012 231140
rect 398972 384524 399028 384580
rect 400652 384412 400708 384468
rect 398972 197820 399028 197876
rect 399084 227724 399140 227780
rect 397292 197708 397348 197764
rect 398972 125132 399028 125188
rect 414092 380156 414148 380212
rect 412412 253148 412468 253204
rect 407372 234332 407428 234388
rect 403004 229404 403060 229460
rect 400652 197372 400708 197428
rect 400988 205772 401044 205828
rect 399084 122668 399140 122724
rect 407036 224364 407092 224420
rect 405020 122668 405076 122724
rect 411068 222684 411124 222740
rect 407372 124236 407428 124292
rect 409052 124236 409108 124292
rect 412412 150556 412468 150612
rect 413084 217644 413140 217700
rect 415772 379036 415828 379092
rect 414092 199836 414148 199892
rect 415100 232764 415156 232820
rect 417452 376796 417508 376852
rect 415772 199948 415828 200004
rect 417116 210812 417172 210868
rect 417452 199724 417508 199780
rect 420028 101500 420084 101556
rect 420028 52780 420084 52836
rect 420140 94892 420196 94948
rect 420140 52668 420196 52724
rect 420252 88172 420308 88228
rect 421708 81452 421764 81508
rect 421708 51772 421764 51828
rect 421820 74732 421876 74788
rect 420252 50652 420308 50708
rect 421932 68012 421988 68068
rect 421932 50540 421988 50596
rect 422044 61292 422100 61348
rect 422044 50428 422100 50484
rect 421820 50316 421876 50372
rect 360556 37772 360612 37828
rect 360332 34412 360388 34468
rect 355404 31052 355460 31108
rect 424172 20300 424228 20356
rect 350476 4956 350532 5012
rect 336812 4396 336868 4452
rect 328412 4172 328468 4228
rect 458556 399532 458612 399588
rect 468636 404460 468692 404516
rect 472892 407820 472948 407876
rect 478380 407708 478436 407764
rect 474684 406140 474740 406196
rect 476252 407596 476308 407652
rect 472892 392924 472948 392980
rect 463932 390908 463988 390964
rect 474572 386652 474628 386708
rect 472892 385644 472948 385700
rect 467852 377916 467908 377972
rect 457772 375676 457828 375732
rect 457772 200172 457828 200228
rect 459452 374556 459508 374612
rect 461132 373436 461188 373492
rect 461132 200284 461188 200340
rect 462812 372316 462868 372372
rect 459452 199388 459508 199444
rect 464492 215852 464548 215908
rect 464492 206668 464548 206724
rect 465948 206668 466004 206724
rect 467852 200396 467908 200452
rect 467964 249564 468020 249620
rect 465948 199612 466004 199668
rect 466284 199612 466340 199668
rect 462812 198940 462868 198996
rect 453516 195916 453572 195972
rect 456092 151900 456148 151956
rect 451052 151676 451108 151732
rect 437612 151564 437668 151620
rect 437612 94892 437668 94948
rect 449372 149436 449428 149492
rect 451052 88172 451108 88228
rect 452732 149212 452788 149268
rect 449372 81452 449428 81508
rect 452732 68012 452788 68068
rect 454412 148652 454468 148708
rect 456316 151788 456372 151844
rect 456316 101612 456372 101668
rect 459452 151228 459508 151284
rect 467964 199500 468020 199556
rect 472892 197484 472948 197540
rect 473004 200844 473060 200900
rect 471660 195804 471716 195860
rect 467852 151900 467908 151956
rect 468972 162316 469028 162372
rect 470316 160860 470372 160916
rect 470316 151228 470372 151284
rect 468972 149660 469028 149716
rect 465724 149436 465780 149492
rect 474572 197596 474628 197652
rect 474684 199276 474740 199332
rect 473004 151676 473060 151732
rect 474684 151564 474740 151620
rect 475692 160972 475748 161028
rect 475692 151788 475748 151844
rect 477932 385532 477988 385588
rect 477932 197932 477988 197988
rect 476252 152124 476308 152180
rect 484652 407932 484708 407988
rect 480060 403004 480116 403060
rect 480508 407372 480564 407428
rect 479612 385420 479668 385476
rect 479612 198156 479668 198212
rect 479724 156380 479780 156436
rect 485436 407820 485492 407876
rect 484652 392812 484708 392868
rect 484876 392812 484932 392868
rect 496188 407932 496244 407988
rect 490812 392700 490868 392756
rect 499772 406812 499828 406868
rect 501564 406812 501620 406868
rect 499772 392588 499828 392644
rect 512316 400764 512372 400820
rect 519820 407932 519876 407988
rect 519708 407820 519764 407876
rect 519372 406700 519428 406756
rect 519260 406588 519316 406644
rect 517692 397964 517748 398020
rect 519148 403564 519204 403620
rect 506940 392476 506996 392532
rect 484876 389228 484932 389284
rect 517468 384188 517524 384244
rect 481628 251580 481684 251636
rect 482748 251468 482804 251524
rect 497308 251356 497364 251412
rect 484988 249900 485044 249956
rect 483868 244524 483924 244580
rect 495068 249788 495124 249844
rect 492828 248220 492884 248276
rect 488348 248108 488404 248164
rect 487228 246204 487284 246260
rect 486108 241500 486164 241556
rect 491708 244412 491764 244468
rect 489468 239932 489524 239988
rect 490588 237692 490644 237748
rect 493948 243068 494004 243124
rect 496188 241388 496244 241444
rect 506268 251244 506324 251300
rect 502908 249676 502964 249732
rect 498428 247996 498484 248052
rect 499548 242956 499604 243012
rect 501788 241276 501844 241332
rect 500668 239820 500724 239876
rect 504028 247884 504084 247940
rect 505148 242844 505204 242900
rect 515228 251132 515284 251188
rect 508508 249452 508564 249508
rect 507388 239708 507444 239764
rect 511868 247772 511924 247828
rect 509628 246092 509684 246148
rect 510748 241164 510804 241220
rect 514108 242732 514164 242788
rect 512988 239596 513044 239652
rect 517468 231868 517524 231924
rect 517580 229180 517636 229236
rect 517468 226492 517524 226548
rect 511644 200396 511700 200452
rect 505372 200284 505428 200340
rect 483420 197708 483476 197764
rect 488124 200060 488180 200116
rect 486556 197820 486612 197876
rect 491260 197596 491316 197652
rect 494396 198156 494452 198212
rect 497532 198156 497588 198212
rect 499100 198156 499156 198212
rect 502236 198156 502292 198212
rect 503132 198940 503188 198996
rect 500668 198044 500724 198100
rect 495964 197932 496020 197988
rect 492828 197484 492884 197540
rect 489692 197372 489748 197428
rect 484988 197260 485044 197316
rect 481852 197148 481908 197204
rect 480508 151340 480564 151396
rect 482412 195916 482468 195972
rect 494508 160748 494564 160804
rect 493164 160636 493220 160692
rect 491820 156604 491876 156660
rect 487788 156492 487844 156548
rect 483756 156268 483812 156324
rect 486444 155372 486500 155428
rect 485100 151452 485156 151508
rect 490476 154700 490532 154756
rect 489132 154588 489188 154644
rect 497196 154140 497252 154196
rect 495852 152908 495908 152964
rect 498540 154028 498596 154084
rect 502572 153132 502628 153188
rect 499884 153020 499940 153076
rect 501340 152908 501396 152964
rect 503804 198940 503860 198996
rect 503132 152012 503188 152068
rect 503916 153916 503972 153972
rect 505260 153804 505316 153860
rect 471884 149436 471940 149492
rect 507948 200284 508004 200340
rect 506492 199388 506548 199444
rect 506940 199388 506996 199444
rect 506828 194124 506884 194180
rect 506828 154476 506884 154532
rect 508508 200172 508564 200228
rect 507948 154140 508004 154196
rect 506492 150668 506548 150724
rect 506604 153692 506660 153748
rect 510076 199724 510132 199780
rect 510300 199388 510356 199444
rect 509852 152124 509908 152180
rect 510076 154364 510132 154420
rect 510636 154476 510692 154532
rect 512428 199948 512484 200004
rect 511644 152236 511700 152292
rect 511980 182364 512036 182420
rect 514892 199836 514948 199892
rect 513436 199164 513492 199220
rect 513212 155372 513268 155428
rect 513324 170604 513380 170660
rect 513436 154476 513492 154532
rect 514668 158956 514724 159012
rect 514892 158956 514948 159012
rect 515004 192444 515060 192500
rect 517356 188972 517412 189028
rect 515004 154364 515060 154420
rect 516012 154476 516068 154532
rect 517580 200284 517636 200340
rect 517692 223804 517748 223860
rect 517804 221676 517860 221732
rect 519820 406700 519876 406756
rect 519708 406588 519764 406644
rect 527436 404348 527492 404404
rect 533820 402892 533876 402948
rect 523068 399420 523124 399476
rect 544572 406028 544628 406084
rect 539196 392364 539252 392420
rect 549500 512764 549556 512820
rect 549500 409612 549556 409668
rect 549612 484428 549668 484484
rect 549388 395500 549444 395556
rect 549612 394492 549668 394548
rect 549724 475468 549780 475524
rect 550060 570332 550116 570388
rect 549836 397404 549892 397460
rect 549948 465612 550004 465668
rect 549724 394156 549780 394212
rect 552748 565068 552804 565124
rect 551852 560252 551908 560308
rect 551180 508620 551236 508676
rect 550284 482860 550340 482916
rect 550060 407372 550116 407428
rect 550172 419244 550228 419300
rect 550284 407932 550340 407988
rect 551068 414540 551124 414596
rect 550172 400652 550228 400708
rect 551180 404124 551236 404180
rect 551292 480396 551348 480452
rect 551068 397740 551124 397796
rect 551292 394268 551348 394324
rect 551404 470988 551460 471044
rect 551516 461580 551572 461636
rect 551628 442764 551684 442820
rect 551628 409276 551684 409332
rect 551740 423948 551796 424004
rect 551516 399196 551572 399252
rect 551852 407708 551908 407764
rect 551964 536844 552020 536900
rect 551740 395724 551796 395780
rect 551404 394044 551460 394100
rect 549948 393932 550004 393988
rect 551964 392252 552020 392308
rect 556108 560364 556164 560420
rect 552860 555660 552916 555716
rect 553532 546252 553588 546308
rect 552972 541548 553028 541604
rect 553196 456876 553252 456932
rect 552972 409836 553028 409892
rect 553084 438060 553140 438116
rect 553196 410508 553252 410564
rect 553308 452172 553364 452228
rect 553532 451948 553588 452004
rect 554428 522732 554484 522788
rect 553420 447468 553476 447524
rect 553420 409500 553476 409556
rect 553532 433356 553588 433412
rect 553308 409388 553364 409444
rect 555212 522508 555268 522564
rect 554428 405804 554484 405860
rect 554540 503916 554596 503972
rect 554540 396060 554596 396116
rect 554652 499212 554708 499268
rect 554652 395948 554708 396004
rect 554764 489804 554820 489860
rect 553532 395836 553588 395892
rect 554764 394380 554820 394436
rect 554876 451948 554932 452004
rect 553084 392812 553140 392868
rect 552860 390796 552916 390852
rect 552748 390684 552804 390740
rect 554988 428652 555044 428708
rect 555212 407596 555268 407652
rect 554988 395612 555044 395668
rect 556444 532140 556500 532196
rect 556220 527436 556276 527492
rect 556220 394604 556276 394660
rect 556332 518028 556388 518084
rect 556444 409724 556500 409780
rect 556556 494508 556612 494564
rect 556556 402668 556612 402724
rect 556892 416780 556948 416836
rect 556892 399084 556948 399140
rect 562604 591276 562660 591332
rect 566972 575372 567028 575428
rect 560252 397628 560308 397684
rect 563612 535724 563668 535780
rect 565292 456428 565348 456484
rect 566972 405692 567028 405748
rect 583772 496076 583828 496132
rect 565292 404012 565348 404068
rect 591276 562156 591332 562212
rect 591276 560252 591332 560308
rect 584668 409052 584724 409108
rect 587132 443212 587188 443268
rect 587132 407820 587188 407876
rect 583772 402556 583828 402612
rect 563612 397516 563668 397572
rect 556332 390572 556388 390628
rect 556108 389116 556164 389172
rect 578732 389788 578788 389844
rect 554876 389004 554932 389060
rect 548492 388892 548548 388948
rect 521612 386540 521668 386596
rect 519932 383180 519988 383236
rect 519932 344316 519988 344372
rect 519372 226492 519428 226548
rect 519484 246876 519540 246932
rect 519484 245868 519540 245924
rect 519372 223804 519428 223860
rect 519148 221676 519204 221732
rect 519260 213052 519316 213108
rect 517804 200844 517860 200900
rect 519148 207676 519204 207732
rect 519148 205324 519204 205380
rect 519148 199724 519204 199780
rect 517692 199276 517748 199332
rect 520044 324268 520100 324324
rect 519372 218428 519428 218484
rect 520156 284620 520212 284676
rect 520156 246876 520212 246932
rect 521612 218540 521668 218596
rect 523292 253036 523348 253092
rect 519596 215740 519652 215796
rect 519484 210812 519540 210868
rect 519484 199500 519540 199556
rect 519372 195804 519428 195860
rect 519260 162316 519316 162372
rect 517468 160972 517524 161028
rect 518700 162204 518756 162260
rect 519596 160860 519652 160916
rect 521388 179004 521444 179060
rect 520044 158844 520100 158900
rect 522732 158732 522788 158788
rect 548492 252924 548548 252980
rect 536172 236796 536228 236852
rect 534828 200508 534884 200564
rect 533372 199052 533428 199108
rect 529452 187404 529508 187460
rect 526652 185612 526708 185668
rect 525420 155708 525476 155764
rect 523292 152348 523348 152404
rect 524076 154364 524132 154420
rect 526652 154476 526708 154532
rect 526764 155596 526820 155652
rect 528108 155484 528164 155540
rect 530796 163884 530852 163940
rect 532140 154476 532196 154532
rect 533372 154476 533428 154532
rect 533484 168812 533540 168868
rect 544236 195692 544292 195748
rect 538860 180572 538916 180628
rect 537516 154476 537572 154532
rect 541772 175532 541828 175588
rect 540204 157276 540260 157332
rect 541548 157164 541604 157220
rect 541772 154476 541828 154532
rect 542892 157052 542948 157108
rect 547148 192332 547204 192388
rect 545580 177212 545636 177268
rect 546924 154476 546980 154532
rect 547148 154476 547204 154532
rect 548268 173852 548324 173908
rect 560252 252812 560308 252868
rect 553644 200620 553700 200676
rect 548492 150780 548548 150836
rect 549612 194012 549668 194068
rect 552300 187292 552356 187348
rect 550956 154476 551012 154532
rect 559468 182252 559524 182308
rect 508844 149548 508900 149604
rect 505484 149436 505540 149492
rect 459900 149324 459956 149380
rect 471660 149212 471716 149268
rect 459900 148652 459956 148708
rect 559468 113708 559524 113764
rect 559580 163772 559636 163828
rect 559804 162092 559860 162148
rect 559580 110572 559636 110628
rect 559692 160524 559748 160580
rect 559916 150444 559972 150500
rect 559916 127596 559972 127652
rect 565292 236572 565348 236628
rect 562828 175644 562884 175700
rect 561708 158956 561764 159012
rect 561372 155372 561428 155428
rect 561148 152124 561204 152180
rect 561148 136668 561204 136724
rect 561260 149436 561316 149492
rect 561596 152236 561652 152292
rect 561372 139804 561428 139860
rect 561484 149212 561540 149268
rect 561708 141372 561764 141428
rect 561596 138236 561652 138292
rect 561484 135100 561540 135156
rect 561260 131964 561316 132020
rect 563164 170492 563220 170548
rect 562828 124124 562884 124180
rect 562940 168924 562996 168980
rect 560252 122444 560308 122500
rect 562828 122444 562884 122500
rect 563052 152348 563108 152404
rect 564508 160412 564564 160468
rect 563388 150780 563444 150836
rect 563164 142940 563220 142996
rect 563276 150556 563332 150612
rect 563388 128828 563444 128884
rect 563276 125692 563332 125748
rect 563052 120988 563108 121044
rect 562940 119420 562996 119476
rect 562828 116284 562884 116340
rect 564732 150668 564788 150724
rect 564620 150332 564676 150388
rect 564732 133532 564788 133588
rect 564620 122556 564676 122612
rect 564508 114716 564564 114772
rect 559804 112140 559860 112196
rect 559692 109116 559748 109172
rect 459452 74732 459508 74788
rect 456092 61292 456148 61348
rect 454412 52892 454468 52948
rect 566188 167132 566244 167188
rect 566300 152012 566356 152068
rect 578732 139244 578788 139300
rect 585452 386428 585508 386484
rect 566300 130396 566356 130452
rect 566188 117852 566244 117908
rect 587132 363916 587188 363972
rect 587132 344316 587188 344372
rect 587132 244972 587188 245028
rect 587132 210812 587188 210868
rect 585452 99820 585508 99876
rect 565292 7084 565348 7140
rect 429212 4172 429268 4228
rect 580636 4172 580692 4228
rect 274876 4060 274932 4116
rect 584444 4172 584500 4228
rect 582540 4060 582596 4116
<< metal3 >>
rect 190418 591276 190428 591332
rect 190484 591276 253708 591332
rect 253764 591276 253774 591332
rect 408258 591276 408268 591332
rect 408324 591276 408362 591332
rect 474310 591276 474348 591332
rect 474404 591276 474414 591332
rect 560242 591276 560252 591332
rect 560308 591276 562604 591332
rect 562660 591276 562670 591332
rect 190530 591164 190540 591220
rect 190596 591164 275772 591220
rect 275828 591164 275838 591220
rect 192770 591052 192780 591108
rect 192836 591052 297836 591108
rect 297892 591052 297902 591108
rect 190642 590940 190652 590996
rect 190708 590940 319900 590996
rect 319956 590940 319966 590996
rect 192994 590828 193004 590884
rect 193060 590828 341964 590884
rect 342020 590828 342030 590884
rect 190306 590716 190316 590772
rect 190372 590716 364028 590772
rect 364084 590716 364094 590772
rect 540754 590716 540764 590772
rect 540820 590716 549836 590772
rect 549892 590716 549902 590772
rect 121538 590604 121548 590660
rect 121604 590604 136892 590660
rect 136948 590604 136958 590660
rect 190530 590604 190540 590660
rect 190596 590604 386092 590660
rect 386148 590604 386158 590660
rect 496626 590604 496636 590660
rect 496692 590604 546028 590660
rect 546084 590604 546094 590660
rect 99474 590492 99484 590548
rect 99540 590492 165452 590548
rect 165508 590492 165518 590548
rect 192658 590492 192668 590548
rect 192724 590492 430220 590548
rect 430276 590492 430286 590548
rect 452498 590492 452508 590548
rect 452564 590492 545580 590548
rect 545636 590492 545646 590548
rect 192882 590380 192892 590436
rect 192948 590380 209580 590436
rect 209636 590380 209646 590436
rect 165666 590156 165676 590212
rect 165732 590156 168812 590212
rect 168868 590156 168878 590212
rect 187730 590156 187740 590212
rect 187796 590156 188972 590212
rect 189028 590156 189038 590212
rect 595560 588644 597000 588840
rect 590482 588588 590492 588644
rect 590548 588616 597000 588644
rect 590548 588588 595672 588616
rect -960 587188 480 587384
rect -960 587160 182252 587188
rect 392 587132 182252 587160
rect 182308 587132 182318 587188
rect 595560 575428 597000 575624
rect 566962 575372 566972 575428
rect 567028 575400 597000 575428
rect 567028 575372 595672 575400
rect -960 573076 480 573272
rect -960 573048 177212 573076
rect 392 573020 177212 573048
rect 177268 573020 177278 573076
rect 190418 572012 190428 572068
rect 190484 572012 231644 572068
rect 231700 572012 231710 572068
rect 77298 570332 77308 570388
rect 77364 570332 148652 570388
rect 148708 570332 148718 570388
rect 518466 570332 518476 570388
rect 518532 570332 550060 570388
rect 550116 570332 550126 570388
rect 184706 565068 184716 565124
rect 184772 565068 190120 565124
rect 549864 565068 552748 565124
rect 552804 565068 552814 565124
rect 595560 562212 597000 562408
rect 591266 562156 591276 562212
rect 591332 562184 597000 562212
rect 591332 562156 595672 562184
rect 549864 560364 556108 560420
rect 556164 560364 556174 560420
rect 551842 560252 551852 560308
rect 551908 560252 591276 560308
rect 591332 560252 591342 560308
rect -960 558964 480 559160
rect -960 558936 4172 558964
rect 392 558908 4172 558936
rect 4228 558908 4238 558964
rect 187842 557900 187852 557956
rect 187908 557900 190120 557956
rect 549864 555660 552860 555716
rect 552916 555660 552926 555716
rect 186386 550732 186396 550788
rect 186452 550732 190120 550788
rect 549388 550452 549444 550984
rect 549378 550396 549388 550452
rect 549444 550396 549454 550452
rect 595560 548996 597000 549192
rect 590594 548940 590604 548996
rect 590660 548968 597000 548996
rect 590660 548940 595672 548968
rect 549864 546252 553532 546308
rect 553588 546252 553598 546308
rect -960 544852 480 545048
rect -960 544824 7532 544852
rect 392 544796 7532 544824
rect 7588 544796 7598 544852
rect 187506 543564 187516 543620
rect 187572 543564 190120 543620
rect 549864 541548 552972 541604
rect 553028 541548 553038 541604
rect 549864 536844 551964 536900
rect 552020 536844 552030 536900
rect 186274 536396 186284 536452
rect 186340 536396 190120 536452
rect 595560 535780 597000 535976
rect 563602 535724 563612 535780
rect 563668 535752 597000 535780
rect 563668 535724 595672 535752
rect 549864 532140 556444 532196
rect 556500 532140 556510 532196
rect -960 530740 480 530936
rect -960 530712 56252 530740
rect 392 530684 56252 530712
rect 56308 530684 56318 530740
rect 187730 529228 187740 529284
rect 187796 529228 190120 529284
rect 549864 527436 556220 527492
rect 556276 527436 556286 527492
rect 549864 522732 554428 522788
rect 554484 522732 554494 522788
rect 595560 522564 597000 522760
rect 555202 522508 555212 522564
rect 555268 522536 597000 522564
rect 555268 522508 595672 522536
rect 187618 522060 187628 522116
rect 187684 522060 190120 522116
rect 549864 518028 556332 518084
rect 556388 518028 556398 518084
rect -960 516628 480 516824
rect -960 516600 4284 516628
rect 392 516572 4284 516600
rect 4340 516572 4350 516628
rect 186162 514892 186172 514948
rect 186228 514892 190120 514948
rect 549500 512820 549556 513352
rect 549490 512764 549500 512820
rect 549556 512764 549566 512820
rect 595560 509348 597000 509544
rect 590706 509292 590716 509348
rect 590772 509320 597000 509348
rect 590772 509292 595672 509320
rect 549864 508620 551180 508676
rect 551236 508620 551246 508676
rect 187394 507724 187404 507780
rect 187460 507724 190120 507780
rect 166226 506492 166236 506548
rect 166292 506492 187404 506548
rect 187460 506492 187470 506548
rect 549864 503916 554540 503972
rect 554596 503916 554606 503972
rect -960 502516 480 502712
rect -960 502488 57932 502516
rect 392 502460 57932 502488
rect 57988 502460 57998 502516
rect 167906 500556 167916 500612
rect 167972 500556 190120 500612
rect 549864 499212 554652 499268
rect 554708 499212 554718 499268
rect 595560 496132 597000 496328
rect 583762 496076 583772 496132
rect 583828 496104 597000 496132
rect 583828 496076 595672 496104
rect 549864 494508 556556 494564
rect 556612 494508 556622 494564
rect 188962 493388 188972 493444
rect 189028 493388 190120 493444
rect 549864 489804 554764 489860
rect 554820 489804 554830 489860
rect -960 488404 480 488600
rect -960 488376 12572 488404
rect 392 488348 12572 488376
rect 12628 488348 12638 488404
rect 189522 486220 189532 486276
rect 189588 486220 190120 486276
rect 549612 484484 549668 485128
rect 549602 484428 549612 484484
rect 549668 484428 549678 484484
rect 595560 482916 597000 483112
rect 550274 482860 550284 482916
rect 550340 482888 597000 482916
rect 550340 482860 595672 482888
rect 549864 480396 551292 480452
rect 551348 480396 551358 480452
rect 189410 479052 189420 479108
rect 189476 479052 190120 479108
rect 4162 476252 4172 476308
rect 4228 476252 146972 476308
rect 147028 476252 147038 476308
rect 549724 475524 549780 475720
rect 549714 475468 549724 475524
rect 549780 475468 549790 475524
rect -960 474292 480 474488
rect -960 474264 141932 474292
rect 392 474236 141932 474264
rect 141988 474236 141998 474292
rect 187954 471884 187964 471940
rect 188020 471884 190120 471940
rect 549864 470988 551404 471044
rect 551460 470988 551470 471044
rect 595560 469700 597000 469896
rect 590818 469644 590828 469700
rect 590884 469672 597000 469700
rect 590884 469644 595672 469672
rect 4274 469532 4284 469588
rect 4340 469532 145292 469588
rect 145348 469532 145358 469588
rect 549836 465668 549892 466312
rect 549836 465612 549948 465668
rect 550004 465612 550014 465668
rect 162530 464716 162540 464772
rect 162596 464716 190120 464772
rect 549864 461580 551516 461636
rect 551572 461580 551582 461636
rect -960 460180 480 460376
rect -960 460152 4172 460180
rect 392 460124 4172 460152
rect 4228 460124 4238 460180
rect 187954 457548 187964 457604
rect 188020 457548 190120 457604
rect 549864 456876 553196 456932
rect 553252 456876 553262 456932
rect 595560 456484 597000 456680
rect 565282 456428 565292 456484
rect 565348 456456 597000 456484
rect 565348 456428 595672 456456
rect 549864 452172 553308 452228
rect 553364 452172 553374 452228
rect 553522 451948 553532 452004
rect 553588 451948 554876 452004
rect 554932 451948 554942 452004
rect 166114 450380 166124 450436
rect 166180 450380 190120 450436
rect 549864 447468 553420 447524
rect 553476 447468 553486 447524
rect -960 446068 480 446264
rect -960 446040 175532 446068
rect 392 446012 175532 446040
rect 175588 446012 175598 446068
rect 595560 443268 597000 443464
rect 167794 443212 167804 443268
rect 167860 443212 190120 443268
rect 587122 443212 587132 443268
rect 587188 443240 597000 443268
rect 587188 443212 595672 443240
rect 549864 442764 551628 442820
rect 551684 442764 551694 442820
rect 549864 438060 553084 438116
rect 553140 438060 553150 438116
rect 187282 436044 187292 436100
rect 187348 436044 190120 436100
rect 549864 433356 553532 433412
rect 553588 433356 553598 433412
rect -960 431956 480 432152
rect -960 431928 140252 431956
rect 392 431900 140252 431928
rect 140308 431900 140318 431956
rect 595560 430164 597000 430248
rect 590930 430108 590940 430164
rect 590996 430108 597000 430164
rect 595560 430024 597000 430108
rect 187394 428876 187404 428932
rect 187460 428876 190120 428932
rect 549864 428652 554988 428708
rect 555044 428652 555054 428708
rect 549864 423948 551740 424004
rect 551796 423948 551806 424004
rect 189298 421708 189308 421764
rect 189364 421708 190120 421764
rect 549864 419244 550172 419300
rect 550228 419244 550238 419300
rect -960 417844 480 418040
rect -960 417816 4172 417844
rect 392 417788 4172 417816
rect 4228 417788 4238 417844
rect 595560 416836 597000 417032
rect 556882 416780 556892 416836
rect 556948 416808 597000 416836
rect 556948 416780 595672 416808
rect 4162 415772 4172 415828
rect 4228 415772 15932 415828
rect 15988 415772 15998 415828
rect 188066 414540 188076 414596
rect 188132 414540 190120 414596
rect 549864 414540 551068 414596
rect 551124 414540 551134 414596
rect 4274 410732 4284 410788
rect 4340 410732 181356 410788
rect 181412 410732 181422 410788
rect 548482 410508 548492 410564
rect 548548 410508 553196 410564
rect 553252 410508 553262 410564
rect 55122 409836 55132 409892
rect 55188 409836 290668 409892
rect 290724 409836 291900 409892
rect 291956 409836 291966 409892
rect 368722 409836 368732 409892
rect 368788 409836 552972 409892
rect 553028 409836 553038 409892
rect 136882 409724 136892 409780
rect 136948 409724 286524 409780
rect 286580 409724 286590 409780
rect 362786 409724 362796 409780
rect 362852 409724 556444 409780
rect 556500 409724 556510 409780
rect 182242 409612 182252 409668
rect 182308 409612 295708 409668
rect 295764 409612 297276 409668
rect 297332 409612 297342 409668
rect 355618 409612 355628 409668
rect 355684 409612 549500 409668
rect 549556 409612 549566 409668
rect 188962 409500 188972 409556
rect 189028 409500 280588 409556
rect 280644 409500 280654 409556
rect 333442 409500 333452 409556
rect 333508 409500 553420 409556
rect 553476 409500 553486 409556
rect 192658 409388 192668 409444
rect 192724 409388 252588 409444
rect 252644 409388 252654 409444
rect 332322 409388 332332 409444
rect 332388 409388 553308 409444
rect 553364 409388 553374 409444
rect 192770 409276 192780 409332
rect 192836 409276 254380 409332
rect 254436 409276 254446 409332
rect 307990 409276 308028 409332
rect 308084 409276 308094 409332
rect 328738 409276 328748 409332
rect 328804 409276 551628 409332
rect 551684 409276 551694 409332
rect 251682 409164 251692 409220
rect 251748 409164 546028 409220
rect 546084 409164 546094 409220
rect 190306 409052 190316 409108
rect 190372 409052 253484 409108
rect 253540 409052 253550 409108
rect 273746 409052 273756 409108
rect 273812 409052 584668 409108
rect 584724 409052 584734 409108
rect 187618 408940 187628 408996
rect 187684 408940 376348 408996
rect 376404 408940 376414 408996
rect 302614 408828 302652 408884
rect 302708 408828 302718 408884
rect 190530 408268 190540 408324
rect 190596 408268 197372 408324
rect 197428 408268 197438 408324
rect 181346 408044 181356 408100
rect 181412 408044 313292 408100
rect 313348 408044 313358 408100
rect 190642 407932 190652 407988
rect 190708 407932 227948 407988
rect 228004 407932 237692 407988
rect 237748 407932 237758 407988
rect 261202 407932 261212 407988
rect 261268 407932 270396 407988
rect 270452 407932 270462 407988
rect 365362 407932 365372 407988
rect 365428 407932 377916 407988
rect 377972 407932 377982 407988
rect 484642 407932 484652 407988
rect 484708 407932 496188 407988
rect 496244 407932 496254 407988
rect 519810 407932 519820 407988
rect 519876 407932 550284 407988
rect 550340 407932 550350 407988
rect 15922 407820 15932 407876
rect 15988 407820 318332 407876
rect 318388 407820 318398 407876
rect 356402 407820 356412 407876
rect 356468 407820 375676 407876
rect 375732 407820 375742 407876
rect 472882 407820 472892 407876
rect 472948 407820 485436 407876
rect 485492 407820 485502 407876
rect 519698 407820 519708 407876
rect 519764 407820 587132 407876
rect 587188 407820 587198 407876
rect 238102 407708 238140 407764
rect 238196 407708 238206 407764
rect 351026 407708 351036 407764
rect 351092 407708 375564 407764
rect 375620 407708 375630 407764
rect 477138 407708 477148 407764
rect 477204 407708 478380 407764
rect 478436 407708 551852 407764
rect 551908 407708 551918 407764
rect 243506 407596 243516 407652
rect 243572 407596 245196 407652
rect 245252 407596 245262 407652
rect 250338 407596 250348 407652
rect 250404 407596 273756 407652
rect 273812 407596 273822 407652
rect 345650 407596 345660 407652
rect 345716 407596 375452 407652
rect 375508 407596 375518 407652
rect 475458 407596 475468 407652
rect 475524 407596 476252 407652
rect 476308 407596 555212 407652
rect 555268 407596 555278 407652
rect 230178 407484 230188 407540
rect 230244 407484 265020 407540
rect 265076 407484 265086 407540
rect 360322 407484 360332 407540
rect 360388 407484 410172 407540
rect 410228 407484 410238 407540
rect 410722 407484 410732 407540
rect 410788 407484 426300 407540
rect 426356 407484 426366 407540
rect 451938 407484 451948 407540
rect 452004 407484 453516 407540
rect 453572 407484 545580 407540
rect 545636 407484 545646 407540
rect 254258 407372 254268 407428
rect 254324 407372 480508 407428
rect 480564 407372 550060 407428
rect 550116 407372 550126 407428
rect 286262 406924 286300 406980
rect 286356 406924 286366 406980
rect 302642 406924 302652 406980
rect 302708 406924 303996 406980
rect 304052 406924 304062 406980
rect 248882 406812 248892 406868
rect 248948 406812 250348 406868
rect 250404 406812 250414 406868
rect 260418 406812 260428 406868
rect 260484 406812 451948 406868
rect 452004 406812 452014 406868
rect 499762 406812 499772 406868
rect 499828 406812 501564 406868
rect 501620 406812 501630 406868
rect 232754 406700 232764 406756
rect 232820 406700 519372 406756
rect 519428 406700 519820 406756
rect 519876 406700 519886 406756
rect 195122 406588 195132 406644
rect 195188 406588 198268 406644
rect 198324 406588 198334 406644
rect 227602 406588 227612 406644
rect 227668 406588 519260 406644
rect 519316 406588 519708 406644
rect 519764 406588 519774 406644
rect 190530 406476 190540 406532
rect 190596 406476 230188 406532
rect 230244 406476 230972 406532
rect 231028 406476 231038 406532
rect 324258 406252 324268 406308
rect 324324 406252 394044 406308
rect 394100 406252 394110 406308
rect 351138 406140 351148 406196
rect 351204 406140 474684 406196
rect 474740 406140 474750 406196
rect 374434 406028 374444 406084
rect 374500 406028 544572 406084
rect 544628 406028 544638 406084
rect 186274 405916 186284 405972
rect 186340 405916 378476 405972
rect 378532 405916 378542 405972
rect 359202 405804 359212 405860
rect 359268 405804 554428 405860
rect 554484 405804 554494 405860
rect 249890 405692 249900 405748
rect 249956 405692 566972 405748
rect 567028 405692 567038 405748
rect 243572 404796 261212 404852
rect 261268 404796 261278 404852
rect 361778 404796 361788 404852
rect 361844 404796 375788 404852
rect 375844 404796 375854 404852
rect 243572 404628 243628 404796
rect 327842 404684 327852 404740
rect 327908 404684 404796 404740
rect 404852 404684 404862 404740
rect 237682 404572 237692 404628
rect 237748 404572 243628 404628
rect 338594 404572 338604 404628
rect 338660 404572 437052 404628
rect 437108 404572 437118 404628
rect 228498 404460 228508 404516
rect 228564 404460 229516 404516
rect 229572 404460 275436 404516
rect 275492 404460 275502 404516
rect 349346 404460 349356 404516
rect 349412 404460 468636 404516
rect 468692 404460 468702 404516
rect 231186 404348 231196 404404
rect 231252 404348 329532 404404
rect 329588 404348 329598 404404
rect 369058 404348 369068 404404
rect 369124 404348 527436 404404
rect 527492 404348 527502 404404
rect 187506 404236 187516 404292
rect 187572 404236 376460 404292
rect 376516 404236 376526 404292
rect 56242 404124 56252 404180
rect 56308 404124 259756 404180
rect 259812 404124 259822 404180
rect 353826 404124 353836 404180
rect 353892 404124 551180 404180
rect 551236 404124 551246 404180
rect 190418 404012 190428 404068
rect 190484 404012 228508 404068
rect 228564 404012 228574 404068
rect 247202 404012 247212 404068
rect 247268 404012 565292 404068
rect 565348 404012 565358 404068
rect -960 403732 480 403928
rect -960 403704 262444 403732
rect 392 403676 262444 403704
rect 262500 403676 262510 403732
rect 595560 403620 597000 403816
rect 502292 403564 519148 403620
rect 519204 403592 597000 403620
rect 519204 403564 595672 403592
rect 502292 403284 502348 403564
rect 222562 403228 222572 403284
rect 222628 403228 502348 403284
rect 340386 403116 340396 403172
rect 340452 403116 442428 403172
rect 442484 403116 442494 403172
rect 352930 403004 352940 403060
rect 352996 403004 480060 403060
rect 480116 403004 480126 403060
rect 370850 402892 370860 402948
rect 370916 402892 533820 402948
rect 533876 402892 533886 402948
rect 187842 402780 187852 402836
rect 187908 402780 375676 402836
rect 375732 402780 375742 402836
rect 12562 402668 12572 402724
rect 12628 402668 260652 402724
rect 260708 402668 260718 402724
rect 348450 402668 348460 402724
rect 348516 402668 556556 402724
rect 556612 402668 556622 402724
rect 111682 402556 111692 402612
rect 111748 402556 232764 402612
rect 232820 402556 232830 402612
rect 248098 402556 248108 402612
rect 248164 402556 583772 402612
rect 583828 402556 583838 402612
rect 231522 402444 231532 402500
rect 231588 402444 590604 402500
rect 590660 402444 590670 402500
rect 231634 402332 231644 402388
rect 231700 402332 590940 402388
rect 590996 402332 591006 402388
rect 322466 402220 322476 402276
rect 322532 402220 388668 402276
rect 388724 402220 388734 402276
rect 367154 401436 367164 401492
rect 367220 401436 375900 401492
rect 375956 401436 375966 401492
rect 326722 401100 326732 401156
rect 326788 401100 372540 401156
rect 372596 401100 372606 401156
rect 331426 400988 331436 401044
rect 331492 400988 415548 401044
rect 415604 400988 415614 401044
rect 236002 400876 236012 400932
rect 236068 400876 334908 400932
rect 334964 400876 334974 400932
rect 342178 400876 342188 400932
rect 342244 400876 447804 400932
rect 447860 400876 447870 400932
rect 231634 400764 231644 400820
rect 231700 400764 340284 400820
rect 340340 400764 340350 400820
rect 363682 400764 363692 400820
rect 363748 400764 512316 400820
rect 512372 400764 512382 400820
rect 175522 400652 175532 400708
rect 175588 400652 261548 400708
rect 261604 400652 261614 400708
rect 319778 400652 319788 400708
rect 319844 400652 550172 400708
rect 550228 400652 550238 400708
rect 336802 399644 336812 399700
rect 336868 399644 431676 399700
rect 431732 399644 431742 399700
rect 345762 399532 345772 399588
rect 345828 399532 458556 399588
rect 458612 399532 458622 399588
rect 367266 399420 367276 399476
rect 367332 399420 523068 399476
rect 523124 399420 523134 399476
rect 186386 399308 186396 399364
rect 186452 399308 378700 399364
rect 378756 399308 378766 399364
rect 165442 399196 165452 399252
rect 165508 399196 257068 399252
rect 257124 399196 257134 399252
rect 335906 399196 335916 399252
rect 335972 399196 551516 399252
rect 551572 399196 551582 399252
rect 246306 399084 246316 399140
rect 246372 399084 556892 399140
rect 556948 399084 556958 399140
rect 234882 398972 234892 399028
rect 234948 398972 590492 399028
rect 590548 398972 590558 399028
rect 343970 398076 343980 398132
rect 344036 398076 453180 398132
rect 453236 398076 453246 398132
rect 365474 397964 365484 398020
rect 365540 397964 517692 398020
rect 517748 397964 517758 398020
rect 184706 397852 184716 397908
rect 184772 397852 378812 397908
rect 378868 397852 378878 397908
rect 168802 397740 168812 397796
rect 168868 397740 256172 397796
rect 256228 397740 256238 397796
rect 317986 397740 317996 397796
rect 318052 397740 551068 397796
rect 551124 397740 551134 397796
rect 250786 397628 250796 397684
rect 250852 397628 560252 397684
rect 560308 397628 560318 397684
rect 248994 397516 249004 397572
rect 249060 397516 563612 397572
rect 563668 397516 563678 397572
rect 233314 397404 233324 397460
rect 233380 397404 549836 397460
rect 549892 397404 549902 397460
rect 230066 397292 230076 397348
rect 230132 397292 590716 397348
rect 590772 397292 590782 397348
rect 189298 396396 189308 396452
rect 189364 396396 378924 396452
rect 378980 396396 378990 396452
rect 187730 396284 187740 396340
rect 187796 396284 376572 396340
rect 376628 396284 376638 396340
rect 186162 396172 186172 396228
rect 186228 396172 378588 396228
rect 378644 396172 378654 396228
rect 352034 396060 352044 396116
rect 352100 396060 554540 396116
rect 554596 396060 554606 396116
rect 350242 395948 350252 396004
rect 350308 395948 554652 396004
rect 554708 395948 554718 396004
rect 330866 395836 330876 395892
rect 330932 395836 553532 395892
rect 553588 395836 553598 395892
rect 321570 395724 321580 395780
rect 321636 395724 551740 395780
rect 551796 395724 551806 395780
rect 323362 395612 323372 395668
rect 323428 395612 554988 395668
rect 555044 395612 555054 395668
rect 369954 395500 369964 395556
rect 370020 395500 549388 395556
rect 549444 395500 549454 395556
rect 335010 394716 335020 394772
rect 335076 394716 410732 394772
rect 410788 394716 410798 394772
rect 360994 394604 361004 394660
rect 361060 394604 556220 394660
rect 556276 394604 556286 394660
rect 344866 394492 344876 394548
rect 344932 394492 549612 394548
rect 549668 394492 549678 394548
rect 346658 394380 346668 394436
rect 346724 394380 554764 394436
rect 554820 394380 554830 394436
rect 343074 394268 343084 394324
rect 343140 394268 551292 394324
rect 551348 394268 551358 394324
rect 341282 394156 341292 394212
rect 341348 394156 549724 394212
rect 549780 394156 549790 394212
rect 231746 394044 231756 394100
rect 231812 394044 260428 394100
rect 260484 394044 260494 394100
rect 339490 394044 339500 394100
rect 339556 394044 551404 394100
rect 551460 394044 551470 394100
rect 190418 393932 190428 393988
rect 190484 393932 255276 393988
rect 255332 393932 255342 393988
rect 337698 393932 337708 393988
rect 337764 393932 549948 393988
rect 550004 393932 550014 393988
rect 229394 393484 229404 393540
rect 229460 393484 304556 393540
rect 304612 393484 304622 393540
rect 106642 393372 106652 393428
rect 106708 393372 316204 393428
rect 316260 393372 316270 393428
rect 103282 393260 103292 393316
rect 103348 393260 315308 393316
rect 315364 393260 315374 393316
rect 40898 393148 40908 393204
rect 40964 393148 292012 393204
rect 292068 393148 292078 393204
rect 322578 393148 322588 393204
rect 322644 393148 324156 393204
rect 324212 393148 372988 393204
rect 373044 393148 373054 393204
rect 326050 393036 326060 393092
rect 326116 393036 399420 393092
rect 399476 393036 399486 393092
rect 354722 392924 354732 392980
rect 354788 392924 472892 392980
rect 472948 392924 472958 392980
rect 358306 392812 358316 392868
rect 358372 392812 484652 392868
rect 484708 392812 484718 392868
rect 484866 392812 484876 392868
rect 484932 392812 553084 392868
rect 553140 392812 553150 392868
rect 356514 392700 356524 392756
rect 356580 392700 490812 392756
rect 490868 392700 490878 392756
rect 360098 392588 360108 392644
rect 360164 392588 499772 392644
rect 499828 392588 499838 392644
rect 236226 392476 236236 392532
rect 236292 392476 290668 392532
rect 290724 392476 290734 392532
rect 361890 392476 361900 392532
rect 361956 392476 506940 392532
rect 506996 392476 507006 392532
rect 237906 392364 237916 392420
rect 237972 392364 295708 392420
rect 295764 392364 295774 392420
rect 318882 392364 318892 392420
rect 318948 392364 365372 392420
rect 365428 392364 365438 392420
rect 372642 392364 372652 392420
rect 372708 392364 539196 392420
rect 539252 392364 539262 392420
rect 236002 392252 236012 392308
rect 236068 392252 322588 392308
rect 322644 392252 322654 392308
rect 329634 392252 329644 392308
rect 329700 392252 360332 392308
rect 360388 392252 360398 392308
rect 364578 392252 364588 392308
rect 364644 392252 551964 392308
rect 552020 392252 552030 392308
rect 320674 392140 320684 392196
rect 320740 392140 383292 392196
rect 383348 392140 383358 392196
rect 229282 392028 229292 392084
rect 229348 392028 305452 392084
rect 305508 392028 305518 392084
rect 204082 391916 204092 391972
rect 204148 391916 314412 391972
rect 314468 391916 314478 391972
rect 120082 391804 120092 391860
rect 120148 391804 310828 391860
rect 310884 391804 310894 391860
rect 103282 391692 103292 391748
rect 103348 391692 307244 391748
rect 307300 391692 307310 391748
rect 100146 391580 100156 391636
rect 100212 391580 312620 391636
rect 312676 391580 312686 391636
rect 99922 391468 99932 391524
rect 99988 391468 313516 391524
rect 313572 391468 313582 391524
rect 399812 391132 409276 391188
rect 409332 391132 409342 391188
rect 419972 391132 420924 391188
rect 420980 391132 420990 391188
rect 399812 390964 399868 391132
rect 419972 391076 420028 391132
rect 371298 390908 371308 390964
rect 371364 390908 399868 390964
rect 405692 391020 420028 391076
rect 405692 390852 405748 391020
rect 409266 390908 409276 390964
rect 409332 390908 463932 390964
rect 463988 390908 463998 390964
rect 333218 390796 333228 390852
rect 333284 390796 405748 390852
rect 421586 390796 421596 390852
rect 421652 390796 552860 390852
rect 552916 390796 552926 390852
rect 177202 390684 177212 390740
rect 177268 390684 258860 390740
rect 258916 390684 258926 390740
rect 379810 390684 379820 390740
rect 379876 390684 552748 390740
rect 552804 390684 552814 390740
rect 33058 390572 33068 390628
rect 33124 390572 257964 390628
rect 258020 390572 258030 390628
rect 357410 390572 357420 390628
rect 357476 390572 556332 390628
rect 556388 390572 556398 390628
rect 245410 390460 245420 390516
rect 245476 390460 377132 390516
rect 377188 390460 377198 390516
rect 595560 390404 597000 390600
rect 242722 390348 242732 390404
rect 242788 390348 382172 390404
rect 382228 390348 382238 390404
rect 590146 390348 590156 390404
rect 590212 390376 597000 390404
rect 590212 390348 595672 390376
rect 240930 390236 240940 390292
rect 240996 390236 380492 390292
rect 380548 390236 380558 390292
rect 104962 390124 104972 390180
rect 105028 390124 311724 390180
rect 311780 390124 311790 390180
rect 100370 390012 100380 390068
rect 100436 390012 309932 390068
rect 309988 390012 309998 390068
rect 10882 389900 10892 389956
rect 10948 389900 270508 389956
rect 270564 389900 270574 389956
rect 272290 389900 272300 389956
rect 272356 389900 429212 389956
rect 429268 389900 429278 389956
rect -960 389620 480 389816
rect 240034 389788 240044 389844
rect 240100 389788 578732 389844
rect 578788 389788 578798 389844
rect 330530 389676 330540 389732
rect 330596 389676 333452 389732
rect 333508 389676 333518 389732
rect 366370 389676 366380 389732
rect 366436 389676 368732 389732
rect 368788 389676 368798 389732
rect -960 389592 4172 389620
rect 392 389564 4172 389592
rect 4228 389564 4238 389620
rect 371746 389340 371756 389396
rect 371812 389340 421596 389396
rect 421652 389340 421662 389396
rect 116722 389228 116732 389284
rect 116788 389228 301868 389284
rect 301924 389228 301934 389284
rect 326946 389228 326956 389284
rect 327012 389228 484876 389284
rect 484932 389228 484942 389284
rect 219202 389116 219212 389172
rect 219268 389116 300972 389172
rect 301028 389116 301038 389172
rect 347554 389116 347564 389172
rect 347620 389116 371308 389172
rect 371364 389116 371374 389172
rect 373538 389116 373548 389172
rect 373604 389116 556108 389172
rect 556164 389116 556174 389172
rect 325154 389004 325164 389060
rect 325220 389004 330876 389060
rect 330932 389004 330942 389060
rect 368162 389004 368172 389060
rect 368228 389004 554876 389060
rect 554932 389004 554942 389060
rect 217522 388892 217532 388948
rect 217588 388892 300076 388948
rect 300132 388892 300142 388948
rect 317090 388892 317100 388948
rect 317156 388892 326732 388948
rect 326788 388892 326798 388948
rect 334114 388892 334124 388948
rect 334180 388892 548492 388948
rect 548548 388892 548558 388948
rect 215842 388780 215852 388836
rect 215908 388780 299180 388836
rect 299236 388780 299246 388836
rect 210802 388668 210812 388724
rect 210868 388668 296492 388724
rect 296548 388668 296558 388724
rect 217746 388556 217756 388612
rect 217812 388556 308140 388612
rect 308196 388556 308206 388612
rect 205762 388444 205772 388500
rect 205828 388444 298284 388500
rect 298340 388444 298350 388500
rect 277666 388332 277676 388388
rect 277732 388332 377244 388388
rect 377300 388332 377310 388388
rect 126802 388220 126812 388276
rect 126868 388220 295596 388276
rect 295652 388220 295662 388276
rect 238214 388108 238252 388164
rect 238308 388108 238318 388164
rect 282118 388108 282156 388164
rect 282212 388108 282222 388164
rect 297350 388108 297388 388164
rect 297444 388108 297454 388164
rect 375330 388108 375340 388164
rect 375396 388108 379820 388164
rect 379876 388108 379886 388164
rect 234994 387324 235004 387380
rect 235060 387324 274092 387380
rect 274148 387324 274158 387380
rect 234770 387212 234780 387268
rect 234836 387212 590156 387268
rect 590212 387212 590222 387268
rect 243618 387100 243628 387156
rect 243684 387100 383852 387156
rect 383908 387100 383918 387156
rect 237346 386988 237356 387044
rect 237412 386988 424172 387044
rect 424228 386988 424238 387044
rect 99922 386876 99932 386932
rect 99988 386876 306348 386932
rect 306404 386876 306414 386932
rect 31042 386764 31052 386820
rect 31108 386764 268716 386820
rect 268772 386764 268782 386820
rect 278562 386764 278572 386820
rect 278628 386764 385532 386820
rect 385588 386764 385598 386820
rect 14242 386652 14252 386708
rect 14308 386652 266924 386708
rect 266980 386652 266990 386708
rect 283938 386652 283948 386708
rect 284004 386652 474572 386708
rect 474628 386652 474638 386708
rect 241826 386540 241836 386596
rect 241892 386540 521612 386596
rect 521668 386540 521678 386596
rect 239138 386428 239148 386484
rect 239204 386428 585452 386484
rect 585508 386428 585518 386484
rect 138562 386316 138572 386372
rect 138628 386316 263340 386372
rect 263396 386316 263406 386372
rect 280354 386316 280364 386372
rect 280420 386316 387212 386372
rect 387268 386316 387278 386372
rect 212482 386204 212492 386260
rect 212548 386204 264236 386260
rect 264292 386204 264302 386260
rect 279458 386204 279468 386260
rect 279524 386204 397292 386260
rect 397348 386204 397358 386260
rect 234546 386092 234556 386148
rect 234612 386092 302764 386148
rect 302820 386092 302830 386148
rect 318322 386092 318332 386148
rect 318388 386092 372316 386148
rect 372372 386092 372382 386148
rect 234322 385980 234332 386036
rect 234388 385980 302988 386036
rect 303044 385980 303054 386036
rect 308802 385980 308812 386036
rect 308868 385980 308878 386036
rect 313282 385980 313292 386036
rect 313348 385980 372428 386036
rect 372484 385980 372494 386036
rect 308812 385924 308868 385980
rect 237794 385868 237804 385924
rect 237860 385868 280588 385924
rect 280644 385868 280654 385924
rect 308812 385868 375564 385924
rect 375620 385868 375630 385924
rect 235106 385756 235116 385812
rect 235172 385756 243852 385812
rect 243908 385756 243918 385812
rect 244514 385756 244524 385812
rect 244580 385756 380604 385812
rect 380660 385756 380670 385812
rect 235666 385644 235676 385700
rect 235732 385644 274988 385700
rect 275044 385644 275054 385700
rect 284834 385644 284844 385700
rect 284900 385644 472892 385700
rect 472948 385644 472958 385700
rect 235778 385532 235788 385588
rect 235844 385532 276780 385588
rect 276836 385532 276846 385588
rect 286626 385532 286636 385588
rect 286692 385532 477932 385588
rect 477988 385532 477998 385588
rect 34402 385420 34412 385476
rect 34468 385420 265132 385476
rect 265188 385420 265198 385476
rect 267782 385420 267820 385476
rect 267876 385420 267886 385476
rect 273158 385420 273196 385476
rect 273252 385420 273262 385476
rect 285730 385420 285740 385476
rect 285796 385420 479612 385476
rect 479668 385420 479678 385476
rect 236086 385308 236124 385364
rect 236180 385308 236190 385364
rect 265990 385308 266028 385364
rect 266084 385308 266094 385364
rect 269574 385308 269612 385364
rect 269668 385308 269678 385364
rect 271366 385308 271404 385364
rect 271460 385308 271470 385364
rect 275846 385308 275884 385364
rect 275940 385308 275950 385364
rect 281222 385308 281260 385364
rect 281316 385308 281326 385364
rect 283014 385308 283052 385364
rect 283108 385308 283118 385364
rect 287494 385308 287532 385364
rect 287588 385308 287598 385364
rect 288390 385308 288428 385364
rect 288484 385308 288494 385364
rect 289286 385308 289324 385364
rect 289380 385308 289390 385364
rect 290182 385308 290220 385364
rect 290276 385308 290286 385364
rect 291078 385308 291116 385364
rect 291172 385308 291182 385364
rect 292870 385308 292908 385364
rect 292964 385308 292974 385364
rect 293766 385308 293804 385364
rect 293860 385308 293870 385364
rect 294662 385308 294700 385364
rect 294756 385308 294766 385364
rect 308998 385308 309036 385364
rect 309092 385308 309102 385364
rect 233426 384524 233436 384580
rect 233492 384524 250348 384580
rect 250404 384524 250414 384580
rect 281250 384524 281260 384580
rect 281316 384524 398972 384580
rect 399028 384524 399038 384580
rect 235666 384412 235676 384468
rect 235732 384412 275884 384468
rect 275940 384412 275950 384468
rect 283042 384412 283052 384468
rect 283108 384412 400652 384468
rect 400708 384412 400718 384468
rect 110002 384300 110012 384356
rect 110068 384300 309036 384356
rect 309092 384300 309102 384356
rect 207442 384188 207452 384244
rect 207508 384188 266028 384244
rect 266084 384188 266094 384244
rect 291106 384188 291116 384244
rect 291172 384188 517468 384244
rect 517524 384188 517534 384244
rect 41122 384076 41132 384132
rect 41188 384076 292908 384132
rect 292964 384076 292974 384132
rect 41010 383964 41020 384020
rect 41076 383964 293804 384020
rect 293860 383964 293870 384020
rect 40226 383852 40236 383908
rect 40292 383852 294700 383908
rect 294756 383852 294766 383908
rect 215954 383180 215964 383236
rect 216020 383180 519932 383236
rect 519988 383180 519998 383236
rect 62402 383068 62412 383124
rect 62468 383068 376348 383124
rect 376404 383068 376414 383124
rect 375928 382396 378924 382452
rect 378980 382396 378990 382452
rect 375928 381276 376348 381332
rect 376404 381276 376414 381332
rect 4162 380492 4172 380548
rect 4228 380492 209132 380548
rect 209188 380492 209198 380548
rect 375928 380156 414092 380212
rect 414148 380156 414158 380212
rect 375928 379036 415772 379092
rect 415828 379036 415838 379092
rect 375928 377916 467852 377972
rect 467908 377916 467918 377972
rect 199714 377468 199724 377524
rect 199780 377468 236040 377524
rect 595560 377188 597000 377384
rect 377122 377132 377132 377188
rect 377188 377160 597000 377188
rect 377188 377132 595672 377160
rect 375928 376796 417452 376852
rect 417508 376796 417518 376852
rect 199490 376348 199500 376404
rect 199556 376348 236040 376404
rect -960 375508 480 375704
rect 375928 375676 457772 375732
rect 457828 375676 457838 375732
rect -960 375480 236012 375508
rect 392 375452 236012 375480
rect 236068 375452 236078 375508
rect 199266 375228 199276 375284
rect 199332 375228 236040 375284
rect 375928 374556 459452 374612
rect 459508 374556 459518 374612
rect 199378 374108 199388 374164
rect 199444 374108 236040 374164
rect 375928 373436 461132 373492
rect 461188 373436 461198 373492
rect 199154 372988 199164 373044
rect 199220 372988 236040 373044
rect 375928 372316 462812 372372
rect 462868 372316 462878 372372
rect 199042 371868 199052 371924
rect 199108 371868 236040 371924
rect 375928 371196 560252 371252
rect 560308 371196 560318 371252
rect 214162 370748 214172 370804
rect 214228 370748 236040 370804
rect 375928 370076 378924 370132
rect 378980 370076 378990 370132
rect 233202 369628 233212 369684
rect 233268 369628 236040 369684
rect 375928 368956 573132 369012
rect 573188 368956 573198 369012
rect 202402 368732 202412 368788
rect 202468 368732 233212 368788
rect 233268 368732 233278 368788
rect 378914 368732 378924 368788
rect 378980 368732 571564 368788
rect 571620 368732 571630 368788
rect 223234 368508 223244 368564
rect 223300 368508 236040 368564
rect 375928 367836 574700 367892
rect 574756 367836 574766 367892
rect 226706 367388 226716 367444
rect 226772 367388 236040 367444
rect 375928 366716 568204 366772
rect 568260 366716 568270 366772
rect 233202 366268 233212 366324
rect 233268 366268 236040 366324
rect 375928 365596 573020 365652
rect 573076 365596 573086 365652
rect 225026 365148 225036 365204
rect 225092 365148 236040 365204
rect 375928 364476 379596 364532
rect 379652 364476 379662 364532
rect 223346 364028 223356 364084
rect 223412 364028 236040 364084
rect 595560 363972 597000 364168
rect 587122 363916 587132 363972
rect 587188 363944 597000 363972
rect 587188 363916 595672 363944
rect 375928 363356 571452 363412
rect 571508 363356 571518 363412
rect 195944 363020 199724 363076
rect 199780 363020 199790 363076
rect 228386 362908 228396 362964
rect 228452 362908 236040 362964
rect 375928 362236 572908 362292
rect 572964 362236 572974 362292
rect 379586 362012 379596 362068
rect 379652 362012 564956 362068
rect 565012 362012 565022 362068
rect 223122 361788 223132 361844
rect 223188 361788 236040 361844
rect -960 361396 480 361592
rect -960 361368 138572 361396
rect 392 361340 138572 361368
rect 138628 361340 138638 361396
rect 375928 361116 379596 361172
rect 379652 361116 379662 361172
rect 232642 360668 232652 360724
rect 232708 360668 236040 360724
rect 375928 359996 566524 360052
rect 566580 359996 566590 360052
rect 195944 359660 199500 359716
rect 199556 359660 199566 359716
rect 226482 359548 226492 359604
rect 226548 359548 236040 359604
rect 375928 358876 571340 358932
rect 571396 358876 571406 358932
rect 379586 358652 379596 358708
rect 379652 358652 569772 358708
rect 569828 358652 569838 358708
rect 228274 358428 228284 358484
rect 228340 358428 236040 358484
rect 375928 357756 571228 357812
rect 571284 357756 571294 357812
rect 226370 357308 226380 357364
rect 226436 357308 236040 357364
rect 375928 356636 569548 356692
rect 569604 356636 569614 356692
rect 195944 356300 199276 356356
rect 199332 356300 199342 356356
rect 236012 356020 236068 356216
rect 236002 355964 236012 356020
rect 236068 355964 236078 356020
rect 375928 355516 569660 355572
rect 569716 355516 569726 355572
rect 226594 355068 226604 355124
rect 226660 355068 236040 355124
rect 375928 354396 566412 354452
rect 566468 354396 566478 354452
rect 230066 353948 230076 354004
rect 230132 353948 236040 354004
rect 375928 353276 564844 353332
rect 564900 353276 564910 353332
rect 195944 352940 199388 352996
rect 199444 352940 199454 352996
rect 228162 352828 228172 352884
rect 228228 352828 236040 352884
rect 375928 352156 379596 352212
rect 379652 352156 379662 352212
rect 234882 351708 234892 351764
rect 234948 351708 236040 351764
rect 375928 351036 567980 351092
rect 568036 351036 568046 351092
rect 595560 350756 597000 350952
rect 590482 350700 590492 350756
rect 590548 350728 597000 350756
rect 590548 350700 595672 350728
rect 227826 350588 227836 350644
rect 227892 350588 236040 350644
rect 379586 350252 379596 350308
rect 379652 350252 568092 350308
rect 568148 350252 568158 350308
rect 375928 349916 566188 349972
rect 566244 349916 566254 349972
rect 195944 349580 199164 349636
rect 199220 349580 199230 349636
rect 228050 349468 228060 349524
rect 228116 349468 236040 349524
rect 375928 348796 564732 348852
rect 564788 348796 564798 348852
rect 229842 348348 229852 348404
rect 229908 348348 236040 348404
rect 375928 347676 566300 347732
rect 566356 347676 566366 347732
rect -960 347284 480 347480
rect -960 347256 4172 347284
rect 392 347228 4172 347256
rect 4228 347228 4238 347284
rect 231522 347228 231532 347284
rect 231588 347228 236040 347284
rect 195916 346892 196588 346948
rect 196644 346892 222572 346948
rect 222628 346892 222638 346948
rect 195916 346248 195972 346892
rect 375928 346556 564620 346612
rect 564676 346556 564686 346612
rect 236124 345940 236180 346136
rect 236114 345884 236124 345940
rect 236180 345884 236190 345940
rect 375928 345436 559580 345492
rect 559636 345436 559646 345492
rect 4162 345212 4172 345268
rect 4228 345212 138572 345268
rect 138628 345212 138638 345268
rect 226258 344988 226268 345044
rect 226324 344988 236040 345044
rect 375928 344316 389116 344372
rect 389172 344316 389182 344372
rect 519922 344316 519932 344372
rect 519988 344316 587132 344372
rect 587188 344316 587198 344372
rect 219986 343868 219996 343924
rect 220052 343868 236040 343924
rect 195916 343532 196700 343588
rect 196756 343532 215964 343588
rect 216020 343532 216030 343588
rect 195916 342888 195972 343532
rect 375928 343196 559468 343252
rect 559524 343196 559534 343252
rect 232754 342748 232764 342804
rect 232820 342748 236040 342804
rect 375928 342076 540092 342132
rect 540148 342076 540158 342132
rect 224914 341628 224924 341684
rect 224980 341628 236040 341684
rect 375928 340956 555212 341012
rect 555268 340956 555278 341012
rect 229730 340508 229740 340564
rect 229796 340508 236040 340564
rect 375928 339836 556892 339892
rect 556948 339836 556958 339892
rect 195804 339332 195860 339528
rect 229954 339500 229964 339556
rect 230020 339500 232652 339556
rect 232708 339500 232718 339556
rect 196140 339388 199220 339444
rect 223010 339388 223020 339444
rect 223076 339388 236040 339444
rect 196140 339332 196196 339388
rect 195804 339276 196196 339332
rect 199164 339220 199220 339388
rect 199154 339164 199164 339220
rect 199220 339164 211260 339220
rect 211316 339164 235900 339220
rect 235956 339164 235966 339220
rect 375928 338716 574588 338772
rect 574644 338716 574654 338772
rect 236236 337988 236292 338296
rect 236226 337932 236236 337988
rect 236292 337932 236302 337988
rect 375928 337596 425852 337652
rect 425908 337596 425918 337652
rect 595560 337540 597000 337736
rect 380594 337484 380604 337540
rect 380660 337512 597000 337540
rect 380660 337484 595672 337512
rect 231410 337148 231420 337204
rect 231476 337148 236040 337204
rect 195916 336812 198380 336868
rect 198436 336812 205884 336868
rect 205940 336812 205950 336868
rect 195916 336168 195972 336812
rect 375928 336476 567868 336532
rect 567924 336476 567934 336532
rect 231298 336028 231308 336084
rect 231364 336028 236040 336084
rect 375928 335356 564508 335412
rect 564564 335356 564574 335412
rect 234770 334908 234780 334964
rect 234836 334908 236040 334964
rect 375928 334236 393932 334292
rect 393988 334236 393998 334292
rect 223346 333788 223356 333844
rect 223412 333788 236040 333844
rect 195916 333452 199052 333508
rect 199108 333452 200508 333508
rect 200564 333452 200574 333508
rect -960 333172 480 333368
rect -960 333144 4172 333172
rect 392 333116 4172 333144
rect 4228 333116 4238 333172
rect 195916 332808 195972 333452
rect 375928 333116 390572 333172
rect 390628 333116 390638 333172
rect 219986 332668 219996 332724
rect 220052 332668 236040 332724
rect 375928 331996 388892 332052
rect 388948 331996 388958 332052
rect 233202 331772 233212 331828
rect 233268 331772 234444 331828
rect 234500 331772 234510 331828
rect 389106 331772 389116 331828
rect 389172 331772 563276 331828
rect 563332 331772 563342 331828
rect 200722 331548 200732 331604
rect 200788 331548 236040 331604
rect 375928 330876 380492 330932
rect 380548 330876 380558 330932
rect 234994 330428 235004 330484
rect 235060 330428 236040 330484
rect 375928 329756 387212 329812
rect 387268 329756 387278 329812
rect 195944 329420 198492 329476
rect 198548 329420 198558 329476
rect 234434 329308 234444 329364
rect 234500 329308 236040 329364
rect 375928 328636 385532 328692
rect 385588 328636 385598 328692
rect 226706 328188 226716 328244
rect 226772 328188 236040 328244
rect 375928 327516 451052 327572
rect 451108 327516 451118 327572
rect 229954 327068 229964 327124
rect 230020 327068 236040 327124
rect 375928 326396 382172 326452
rect 382228 326396 382238 326452
rect 195944 326060 199052 326116
rect 199108 326060 199118 326116
rect 227714 326060 227724 326116
rect 227780 326060 232764 326116
rect 232820 326060 232830 326116
rect 228386 325948 228396 326004
rect 228452 325948 236040 326004
rect 375928 325276 392252 325332
rect 392308 325276 392318 325332
rect 231410 324828 231420 324884
rect 231476 324828 236040 324884
rect 595560 324324 597000 324520
rect 520006 324268 520044 324324
rect 520100 324296 597000 324324
rect 520100 324268 595672 324296
rect 375928 324156 383852 324212
rect 383908 324156 383918 324212
rect 226594 323708 226604 323764
rect 226660 323708 236040 323764
rect 195468 323372 227612 323428
rect 227668 323372 227678 323428
rect 195468 322756 195524 323372
rect 375928 323036 456092 323092
rect 456148 323036 456158 323092
rect 195234 322700 195244 322756
rect 195300 322728 195524 322756
rect 195300 322700 195496 322728
rect 231298 322588 231308 322644
rect 231364 322588 236040 322644
rect 4162 322476 4172 322532
rect 4228 322476 173068 322532
rect 173012 322308 173068 322476
rect 203252 322476 231196 322532
rect 231252 322476 231868 322532
rect 231924 322476 231934 322532
rect 203252 322420 203308 322476
rect 199892 322364 203308 322420
rect 199892 322308 199948 322364
rect 173012 322252 199948 322308
rect 173012 321916 195244 321972
rect 195300 321916 195310 321972
rect 375928 321916 442652 321972
rect 442708 321916 442718 321972
rect 173012 321748 173068 321916
rect 113362 321692 113372 321748
rect 113428 321692 173068 321748
rect 229842 321468 229852 321524
rect 229908 321468 236040 321524
rect 231186 320348 231196 320404
rect 231252 320348 236040 320404
rect 375900 320068 375956 320824
rect 115042 320012 115052 320068
rect 115108 320012 199164 320068
rect 199220 320012 199230 320068
rect 375900 320012 378812 320068
rect 378868 320012 437612 320068
rect 437668 320012 437678 320068
rect 375666 319676 375676 319732
rect 375732 319676 434252 319732
rect 434308 319676 434318 319732
rect -960 319060 480 319256
rect 232418 319228 232428 319284
rect 232484 319228 236040 319284
rect -960 319032 212492 319060
rect 392 319004 212492 319032
rect 212548 319004 212558 319060
rect 375900 318388 375956 318584
rect 375900 318332 378700 318388
rect 378756 318332 432572 318388
rect 432628 318332 432638 318388
rect 233202 318108 233212 318164
rect 233268 318108 236040 318164
rect 375928 317436 376460 317492
rect 376516 317436 378812 317492
rect 378868 317436 378878 317492
rect 233314 316988 233324 317044
rect 233380 316988 236040 317044
rect 375900 316652 378476 316708
rect 378532 316652 427532 316708
rect 427588 316652 427598 316708
rect 375900 316344 375956 316652
rect 233090 315868 233100 315924
rect 233156 315868 236040 315924
rect 375928 315196 376572 315252
rect 376628 315196 376638 315252
rect 376572 315028 376628 315196
rect 378802 315084 378812 315140
rect 378868 315084 430892 315140
rect 430948 315084 430958 315140
rect 376572 314972 429212 315028
rect 429268 314972 429278 315028
rect 232642 314748 232652 314804
rect 232708 314748 236040 314804
rect 375928 314104 376348 314132
rect 375900 314076 376348 314104
rect 376404 314076 376414 314132
rect 232530 313628 232540 313684
rect 232596 313628 236040 313684
rect 375900 313348 375956 314076
rect 378578 313404 378588 313460
rect 378644 313404 425964 313460
rect 426020 313404 426030 313460
rect 181346 313292 181356 313348
rect 181412 313292 214172 313348
rect 214228 313292 214238 313348
rect 375900 313292 454412 313348
rect 454468 313292 454478 313348
rect 375928 312956 378588 313012
rect 378644 312956 378654 313012
rect 232866 312508 232876 312564
rect 232932 312508 236040 312564
rect 375928 311836 379036 311892
rect 379092 311836 379102 311892
rect 10994 311612 11004 311668
rect 11060 311612 215964 311668
rect 216020 311612 216030 311668
rect 232754 311388 232764 311444
rect 232820 311388 236040 311444
rect 595560 311108 597000 311304
rect 590594 311052 590604 311108
rect 590660 311080 597000 311108
rect 590660 311052 595672 311080
rect 375928 310716 378924 310772
rect 378980 310716 378990 310772
rect 232978 310268 232988 310324
rect 233044 310268 236040 310324
rect 375928 309596 383068 309652
rect 383124 309596 383134 309652
rect 233202 309148 233212 309204
rect 233268 309148 236040 309204
rect 375928 308476 384748 308532
rect 384804 308476 384814 308532
rect 233090 308028 233100 308084
rect 233156 308028 236040 308084
rect 375928 307356 378812 307412
rect 378868 307356 378878 307412
rect 227490 306908 227500 306964
rect 227556 306908 236040 306964
rect 375928 306236 379484 306292
rect 379540 306236 379550 306292
rect 4162 305788 4172 305844
rect 4228 305788 236040 305844
rect -960 304948 480 305144
rect 375928 305116 379372 305172
rect 379428 305116 379438 305172
rect -960 304920 228284 304948
rect 392 304892 228284 304920
rect 228340 304892 228350 304948
rect 4274 304668 4284 304724
rect 4340 304668 236040 304724
rect 227938 303996 227948 304052
rect 228004 303996 229628 304052
rect 229684 303996 229694 304052
rect 375928 303996 379260 304052
rect 379316 303996 379326 304052
rect 29362 303548 29372 303604
rect 29428 303548 236040 303604
rect 77410 303212 77420 303268
rect 77476 303212 227948 303268
rect 228004 303212 228014 303268
rect 375928 302876 379036 302932
rect 379092 302876 379102 302932
rect 32722 302540 32732 302596
rect 32788 302540 236068 302596
rect 236012 302456 236068 302540
rect 375928 301756 378924 301812
rect 378980 301756 378990 301812
rect 92418 301532 92428 301588
rect 92484 301532 229516 301588
rect 229572 301532 229582 301588
rect 27794 301308 27804 301364
rect 27860 301308 236040 301364
rect 229506 300748 229516 300804
rect 229572 300748 230972 300804
rect 231028 300748 231038 300804
rect 375928 300636 379148 300692
rect 379204 300636 379214 300692
rect 12562 300188 12572 300244
rect 12628 300188 236040 300244
rect 375928 299516 378812 299572
rect 378868 299516 378878 299572
rect 31892 299404 55468 299460
rect 31892 299348 31948 299404
rect 55412 299348 55468 299404
rect 10882 299292 10892 299348
rect 10948 299292 31948 299348
rect 47366 299292 47404 299348
rect 47460 299292 47470 299348
rect 55412 299292 236068 299348
rect 236012 299096 236068 299292
rect 375928 298396 376348 298452
rect 376404 298396 376414 298452
rect 228274 297948 228284 298004
rect 228340 297948 236040 298004
rect 595560 297892 597000 298088
rect 383842 297836 383852 297892
rect 383908 297864 597000 297892
rect 383908 297836 595672 297864
rect 4162 297500 4172 297556
rect 4228 297500 227612 297556
rect 227668 297500 227678 297556
rect 47394 297388 47404 297444
rect 47460 297388 48524 297444
rect 48580 297388 163772 297444
rect 163828 297388 163838 297444
rect 375928 297276 377132 297332
rect 377188 297276 377198 297332
rect 138562 296828 138572 296884
rect 138628 296828 236040 296884
rect 375928 296156 376572 296212
rect 376628 296156 376638 296212
rect 99960 296044 186508 296100
rect 186564 296044 187292 296100
rect 187348 296044 187358 296100
rect 209122 295708 209132 295764
rect 209188 295708 236040 295764
rect 375928 295036 379708 295092
rect 379764 295036 379774 295092
rect 140242 294588 140252 294644
rect 140308 294588 236040 294644
rect 375928 293916 376684 293972
rect 376740 293916 376750 293972
rect 141922 293468 141932 293524
rect 141988 293468 236040 293524
rect 375928 292796 378364 292852
rect 378420 292796 378430 292852
rect 145282 292348 145292 292404
rect 145348 292348 236040 292404
rect 375928 291676 378476 291732
rect 378532 291676 378542 291732
rect 146962 291228 146972 291284
rect 147028 291228 236040 291284
rect 392 291032 4172 291060
rect -960 291004 4172 291032
rect 4228 291004 4238 291060
rect -960 290808 480 291004
rect 163762 290556 163772 290612
rect 163828 290556 188076 290612
rect 188132 290556 188142 290612
rect 375928 290556 376796 290612
rect 376852 290556 376862 290612
rect 99960 290220 187404 290276
rect 187460 290220 187470 290276
rect 215954 290108 215964 290164
rect 216020 290108 236040 290164
rect 172834 289884 172844 289940
rect 172900 289884 202412 289940
rect 202468 289884 202478 289940
rect 375928 289436 411740 289492
rect 411796 289436 411806 289492
rect 173012 289100 196588 289156
rect 173012 289044 173068 289100
rect 196532 289044 196588 289100
rect 148642 288988 148652 289044
rect 148708 288988 173068 289044
rect 186610 288988 186620 289044
rect 186676 288988 187404 289044
rect 187460 288988 187470 289044
rect 188066 288988 188076 289044
rect 188132 288988 192332 289044
rect 192388 288988 192398 289044
rect 196532 288988 236040 289044
rect 375218 288316 375228 288372
rect 375284 288316 375294 288372
rect 143378 287868 143388 287924
rect 143444 287868 236040 287924
rect 375928 287196 378588 287252
rect 378644 287196 378654 287252
rect 192882 286748 192892 286804
rect 192948 286748 236040 286804
rect 167794 286636 167804 286692
rect 167860 286636 188300 286692
rect 188356 286636 188366 286692
rect 162530 286524 162540 286580
rect 162596 286524 188524 286580
rect 188580 286524 188590 286580
rect 103394 286412 103404 286468
rect 103460 286412 196700 286468
rect 196756 286412 196766 286468
rect 375218 286076 375228 286132
rect 375284 286076 375294 286132
rect 197474 285628 197484 285684
rect 197540 285628 236040 285684
rect 167906 285516 167916 285572
rect 167972 285516 188188 285572
rect 188244 285516 188254 285572
rect 166114 285404 166124 285460
rect 166180 285404 188412 285460
rect 188468 285404 188478 285460
rect 103506 285292 103516 285348
rect 103572 285292 196588 285348
rect 196644 285292 196654 285348
rect 375928 284956 378252 285012
rect 378308 284956 378318 285012
rect 197362 284732 197372 284788
rect 197428 284732 198380 284788
rect 198436 284732 198446 284788
rect 595560 284676 597000 284872
rect 520146 284620 520156 284676
rect 520212 284648 597000 284676
rect 520212 284620 595672 284648
rect 192994 284508 193004 284564
rect 193060 284508 236040 284564
rect 379026 284508 379036 284564
rect 379092 284508 379820 284564
rect 379876 284508 379886 284564
rect 99960 284396 111692 284452
rect 111748 284396 111758 284452
rect 166226 284172 166236 284228
rect 166292 284172 185892 284228
rect 185836 284004 185892 284172
rect 185836 283976 234668 284004
rect 185864 283948 234668 283976
rect 234724 283948 234734 284004
rect 379810 283948 379820 284004
rect 379876 283948 424172 284004
rect 424228 283948 424238 284004
rect 375666 283836 375676 283892
rect 375732 283836 375742 283892
rect 190642 283388 190652 283444
rect 190708 283388 236040 283444
rect 375928 282716 378028 282772
rect 378084 282716 378094 282772
rect 193106 282268 193116 282324
rect 193172 282268 236040 282324
rect 378914 282156 378924 282212
rect 378980 282156 379932 282212
rect 379988 282156 379998 282212
rect 185836 281428 185892 281960
rect 375928 281596 376460 281652
rect 376516 281596 376526 281652
rect 185836 281372 188188 281428
rect 188244 281372 234220 281428
rect 234276 281372 234286 281428
rect 233314 281148 233324 281204
rect 233380 281148 236040 281204
rect 379922 280588 379932 280644
rect 379988 280588 420812 280644
rect 420868 280588 420878 280644
rect 375928 280476 377020 280532
rect 377076 280476 377086 280532
rect 234882 280028 234892 280084
rect 234948 280028 236040 280084
rect 185864 279916 188972 279972
rect 189028 279916 189038 279972
rect 375928 279356 378700 279412
rect 378756 279356 378766 279412
rect 231522 278908 231532 278964
rect 231588 278908 236040 278964
rect 99960 278572 113372 278628
rect 113428 278572 113438 278628
rect 375928 278236 411628 278292
rect 411684 278236 411694 278292
rect 185836 278012 189532 278068
rect 189588 278012 231084 278068
rect 231140 278012 231150 278068
rect 185836 277928 185892 278012
rect 230066 277788 230076 277844
rect 230132 277788 236040 277844
rect 375928 277116 378924 277172
rect 378980 277116 378990 277172
rect -960 276724 480 276920
rect -960 276696 34412 276724
rect 392 276668 34412 276696
rect 34468 276668 34478 276724
rect 231746 276668 231756 276724
rect 231812 276668 236040 276724
rect 185836 276332 189420 276388
rect 189476 276332 231084 276388
rect 231140 276332 231150 276388
rect 185836 275912 185892 276332
rect 375928 275996 376348 276052
rect 376404 275996 376414 276052
rect 231634 275548 231644 275604
rect 231700 275548 236040 275604
rect 378802 275548 378812 275604
rect 378868 275548 380044 275604
rect 380100 275548 452732 275604
rect 452788 275548 452798 275604
rect 375928 274876 378140 274932
rect 378196 274876 378206 274932
rect 234770 274428 234780 274484
rect 234836 274428 236040 274484
rect 185864 273868 188636 273924
rect 188692 273868 189084 273924
rect 189140 273868 189150 273924
rect 379474 273868 379484 273924
rect 379540 273868 380268 273924
rect 380324 273868 440972 273924
rect 441028 273868 441038 273924
rect 375928 273756 376460 273812
rect 376516 273756 376526 273812
rect 235778 273308 235788 273364
rect 235844 273308 236040 273364
rect 99960 272748 103516 272804
rect 103572 272748 103582 272804
rect 375928 272636 411852 272692
rect 411908 272636 411918 272692
rect 231746 272188 231756 272244
rect 231812 272188 236040 272244
rect 185836 271348 185892 271880
rect 375778 271516 375788 271572
rect 375844 271516 375854 271572
rect 595560 271460 597000 271656
rect 590818 271404 590828 271460
rect 590884 271432 597000 271460
rect 590884 271404 595672 271432
rect 185836 271292 188524 271348
rect 188580 271292 231532 271348
rect 231588 271292 231598 271348
rect 235106 271068 235116 271124
rect 235172 271068 236040 271124
rect 379810 270508 379820 270564
rect 379876 270508 447692 270564
rect 447748 270508 447758 270564
rect 375890 270396 375900 270452
rect 375956 270396 375966 270452
rect 379250 270396 379260 270452
rect 379316 270396 380044 270452
rect 380100 270396 380110 270452
rect 235330 269948 235340 270004
rect 235396 269948 236040 270004
rect 185864 269836 187964 269892
rect 188020 269836 189532 269892
rect 189588 269836 189598 269892
rect 375928 269276 379036 269332
rect 379092 269276 379102 269332
rect 234658 268828 234668 268884
rect 234724 268828 236040 268884
rect 380034 268828 380044 268884
rect 380100 268828 446012 268884
rect 446068 268828 446078 268884
rect 379026 268716 379036 268772
rect 379092 268716 379932 268772
rect 379988 268716 379998 268772
rect 375928 268156 381388 268212
rect 381444 268156 381454 268212
rect 185836 267932 188412 267988
rect 188468 267932 235676 267988
rect 235732 267932 235742 267988
rect 185836 267848 185892 267932
rect 234882 267708 234892 267764
rect 234948 267708 236040 267764
rect 379922 267148 379932 267204
rect 379988 267148 444332 267204
rect 444388 267148 444398 267204
rect 375928 267036 378588 267092
rect 378644 267036 378654 267092
rect 99960 266924 103404 266980
rect 103460 266924 103470 266980
rect 234546 266588 234556 266644
rect 234612 266588 236040 266644
rect 185836 266252 188300 266308
rect 188356 266252 235900 266308
rect 235956 266252 235966 266308
rect 185836 265832 185892 266252
rect 375218 265916 375228 265972
rect 375284 265916 375294 265972
rect 234770 265468 234780 265524
rect 234836 265468 236040 265524
rect 378914 265468 378924 265524
rect 378980 265468 379708 265524
rect 379764 265468 449372 265524
rect 449428 265468 449438 265524
rect 375928 264796 378700 264852
rect 378756 264796 378766 264852
rect 185836 264572 186508 264628
rect 186564 264572 235564 264628
rect 235620 264572 235630 264628
rect 185836 263816 185892 264572
rect 233314 264348 233324 264404
rect 233380 264348 236040 264404
rect 379138 263788 379148 263844
rect 379204 263788 380156 263844
rect 380212 263788 419356 263844
rect 419412 263788 419422 263844
rect 375928 263676 378924 263732
rect 378980 263676 378990 263732
rect 392 262808 10892 262836
rect -960 262780 10892 262808
rect 10948 262780 10958 262836
rect -960 262584 480 262780
rect 375928 262556 378476 262612
rect 378532 262556 378542 262612
rect 185864 261772 186620 261828
rect 186676 261772 189196 261828
rect 189252 261772 189262 261828
rect 375928 261436 376124 261492
rect 376180 261436 376190 261492
rect 99960 261100 115052 261156
rect 115108 261100 115118 261156
rect 378802 260428 378812 260484
rect 378868 260428 422492 260484
rect 422548 260428 422558 260484
rect 375928 260316 376908 260372
rect 376964 260316 376974 260372
rect 375928 259196 376236 259252
rect 376292 259196 376302 259252
rect 595560 258244 597000 258440
rect 382162 258188 382172 258244
rect 382228 258216 597000 258244
rect 382228 258188 595672 258216
rect 237570 257404 237580 257460
rect 237636 257404 380044 257460
rect 380100 257404 380110 257460
rect 233090 257292 233100 257348
rect 233156 257292 269276 257348
rect 269332 257292 269342 257348
rect 348562 257292 348572 257348
rect 348628 257292 378476 257348
rect 378532 257292 378542 257348
rect 102498 257068 102508 257124
rect 102564 257068 196476 257124
rect 196532 257068 197372 257124
rect 197428 257068 197438 257124
rect 235778 256508 235788 256564
rect 235844 256508 590492 256564
rect 590548 256508 590558 256564
rect 234658 256396 234668 256452
rect 234724 256396 379820 256452
rect 379876 256396 379886 256452
rect 235890 256284 235900 256340
rect 235956 256284 379708 256340
rect 379764 256284 379774 256340
rect 232530 256172 232540 256228
rect 232596 256172 273868 256228
rect 273924 256172 273934 256228
rect 331772 256172 378588 256228
rect 378644 256172 378654 256228
rect 233202 256060 233212 256116
rect 233268 256060 267148 256116
rect 267092 255892 267148 256060
rect 331772 256004 331828 256172
rect 350476 256060 378364 256116
rect 378420 256060 378430 256116
rect 350476 256004 350532 256060
rect 331762 255948 331772 256004
rect 331828 255948 331838 256004
rect 350466 255948 350476 256004
rect 350532 255948 350542 256004
rect 362002 255948 362012 256004
rect 362068 255948 375788 256004
rect 375844 255948 375854 256004
rect 267092 255836 273868 255892
rect 273924 255836 273934 255892
rect 362114 255836 362124 255892
rect 362180 255836 375900 255892
rect 375956 255836 375966 255892
rect 235442 255724 235452 255780
rect 235508 255724 379932 255780
rect 379988 255724 379998 255780
rect 99960 255276 102508 255332
rect 102564 255276 102574 255332
rect 231746 255276 231756 255332
rect 231812 255276 590604 255332
rect 590660 255276 590670 255332
rect 235106 255164 235116 255220
rect 235172 255164 590828 255220
rect 590884 255164 590894 255220
rect 189186 255052 189196 255108
rect 189252 255052 378812 255108
rect 378868 255052 378878 255108
rect 231074 254940 231084 254996
rect 231140 254940 380044 254996
rect 380100 254940 380110 254996
rect 234210 254828 234220 254884
rect 234276 254828 379932 254884
rect 379988 254828 379998 254884
rect 235778 254716 235788 254772
rect 235844 254716 380156 254772
rect 380212 254716 380222 254772
rect 232642 254604 232652 254660
rect 232708 254604 273980 254660
rect 274036 254604 274046 254660
rect 330082 254604 330092 254660
rect 330148 254604 378252 254660
rect 378308 254604 378318 254660
rect 233314 254492 233324 254548
rect 233380 254492 326732 254548
rect 326788 254492 326798 254548
rect 328402 254492 328412 254548
rect 328468 254492 378140 254548
rect 378196 254492 378206 254548
rect 336802 254380 336812 254436
rect 336868 254380 378028 254436
rect 378084 254380 378094 254436
rect 192322 253596 192332 253652
rect 192388 253596 242732 253652
rect 242788 253596 242798 253652
rect 251878 253596 251916 253652
rect 251972 253596 251982 253652
rect 252550 253596 252588 253652
rect 252644 253596 252654 253652
rect 258822 253596 258860 253652
rect 258916 253596 258926 253652
rect 259718 253596 259756 253652
rect 259812 253596 259822 253652
rect 260614 253596 260652 253652
rect 260708 253596 260718 253652
rect 266018 253484 266028 253540
rect 266084 253484 275660 253540
rect 275716 253484 275726 253540
rect 290322 253372 290332 253428
rect 290388 253372 298284 253428
rect 298340 253372 298350 253428
rect 358642 253372 358652 253428
rect 358708 253372 376796 253428
rect 376852 253372 376862 253428
rect 264226 253260 264236 253316
rect 264292 253260 275548 253316
rect 275604 253260 275614 253316
rect 288306 253260 288316 253316
rect 288372 253260 296492 253316
rect 296548 253260 296558 253316
rect 355282 253260 355292 253316
rect 355348 253260 373772 253316
rect 373828 253260 373838 253316
rect 265122 253148 265132 253204
rect 265188 253148 279020 253204
rect 279076 253148 279086 253204
rect 284946 253148 284956 253204
rect 285012 253148 295596 253204
rect 295652 253148 295662 253204
rect 367266 253148 367276 253204
rect 367332 253148 412412 253204
rect 412468 253148 412478 253204
rect 263330 253036 263340 253092
rect 263396 253036 277228 253092
rect 277284 253036 277294 253092
rect 284722 253036 284732 253092
rect 284788 253036 300972 253092
rect 301028 253036 301038 253092
rect 364578 253036 364588 253092
rect 364644 253036 523292 253092
rect 523348 253036 523358 253092
rect 261538 252924 261548 252980
rect 261604 252924 277340 252980
rect 277396 252924 277406 252980
rect 283378 252924 283388 252980
rect 283444 252924 300076 252980
rect 300132 252924 300142 252980
rect 312610 252924 312620 252980
rect 312676 252924 320012 252980
rect 320068 252924 320078 252980
rect 369058 252924 369068 252980
rect 369124 252924 548492 252980
rect 548548 252924 548558 252980
rect 262434 252812 262444 252868
rect 262500 252812 278908 252868
rect 278964 252812 278974 252868
rect 281362 252812 281372 252868
rect 281428 252812 299180 252868
rect 299236 252812 299246 252868
rect 310818 252812 310828 252868
rect 310884 252812 321692 252868
rect 321748 252812 321758 252868
rect 360994 252812 361004 252868
rect 361060 252812 560252 252868
rect 560308 252812 560318 252868
rect 289762 252700 289772 252756
rect 289828 252700 294700 252756
rect 294756 252700 294766 252756
rect 283154 252476 283164 252532
rect 283220 252476 291116 252532
rect 291172 252476 291182 252532
rect 290612 252364 292012 252420
rect 292068 252364 292078 252420
rect 319778 252364 319788 252420
rect 319844 252364 323484 252420
rect 323540 252364 323550 252420
rect 290612 252308 290668 252364
rect 267810 252252 267820 252308
rect 267876 252252 277564 252308
rect 277620 252252 277630 252308
rect 289986 252252 289996 252308
rect 290052 252252 290668 252308
rect 290882 252252 290892 252308
rect 290948 252252 297388 252308
rect 297444 252252 297454 252308
rect 321570 252252 321580 252308
rect 321636 252252 325388 252308
rect 325444 252252 325454 252308
rect 366370 252252 366380 252308
rect 366436 252252 372988 252308
rect 268706 252140 268716 252196
rect 268772 252140 277452 252196
rect 277508 252140 277518 252196
rect 291106 252140 291116 252196
rect 291172 252140 293804 252196
rect 293860 252140 293870 252196
rect 301858 252140 301868 252196
rect 301924 252140 304892 252196
rect 304948 252140 304958 252196
rect 317090 252140 317100 252196
rect 317156 252140 320236 252196
rect 320292 252140 320302 252196
rect 325154 252140 325164 252196
rect 325220 252140 326844 252196
rect 326900 252140 326910 252196
rect 361890 252140 361900 252196
rect 361956 252140 370412 252196
rect 370468 252140 370478 252196
rect 372932 252084 372988 252252
rect 266914 252028 266924 252084
rect 266980 252028 269724 252084
rect 269780 252028 269790 252084
rect 272290 252028 272300 252084
rect 272356 252028 279132 252084
rect 279188 252028 279198 252084
rect 288082 252028 288092 252084
rect 288148 252028 289324 252084
rect 289380 252028 289390 252084
rect 291442 252028 291452 252084
rect 291508 252028 292908 252084
rect 292964 252028 292974 252084
rect 304546 252028 304556 252084
rect 304612 252028 310044 252084
rect 310100 252028 310110 252084
rect 313506 252028 313516 252084
rect 313572 252028 314972 252084
rect 315028 252028 315038 252084
rect 316194 252028 316204 252084
rect 316260 252028 318332 252084
rect 318388 252028 318398 252084
rect 318882 252028 318892 252084
rect 318948 252028 321916 252084
rect 321972 252028 321982 252084
rect 326050 252028 326060 252084
rect 326116 252028 331884 252084
rect 331940 252028 331950 252084
rect 332322 252028 332332 252084
rect 332388 252028 333452 252084
rect 333508 252028 333518 252084
rect 334114 252028 334124 252084
rect 334180 252028 335132 252084
rect 335188 252028 335198 252084
rect 343074 252028 343084 252084
rect 343140 252028 345212 252084
rect 345268 252028 345278 252084
rect 355618 252028 355628 252084
rect 355684 252028 356972 252084
rect 357028 252028 357038 252084
rect 363682 252028 363692 252084
rect 363748 252028 372092 252084
rect 372148 252028 372158 252084
rect 372932 252028 376012 252084
rect 376068 252028 376078 252084
rect 189074 251916 189084 251972
rect 189140 251916 380268 251972
rect 380324 251916 380334 251972
rect 358978 251804 358988 251860
rect 359044 251804 376348 251860
rect 376404 251804 376414 251860
rect 227602 251692 227612 251748
rect 227668 251692 236012 251748
rect 236068 251692 272188 251748
rect 272244 251692 272254 251748
rect 358754 251692 358764 251748
rect 358820 251692 377020 251748
rect 377076 251692 377086 251748
rect 234770 251580 234780 251636
rect 234836 251580 481628 251636
rect 481684 251580 481694 251636
rect 231298 251468 231308 251524
rect 231364 251468 482748 251524
rect 482804 251468 482814 251524
rect 227826 251356 227836 251412
rect 227892 251356 497308 251412
rect 497364 251356 497374 251412
rect 226482 251244 226492 251300
rect 226548 251244 506268 251300
rect 506324 251244 506334 251300
rect 223234 251132 223244 251188
rect 223300 251132 515228 251188
rect 515284 251132 515294 251188
rect 359202 251020 359212 251076
rect 359268 251020 376460 251076
rect 376516 251020 376526 251076
rect 231522 250236 231532 250292
rect 231588 250236 379820 250292
rect 379876 250236 379886 250292
rect 256162 250124 256172 250180
rect 256228 250124 270620 250180
rect 270676 250124 270686 250180
rect 230962 250012 230972 250068
rect 231028 250012 273980 250068
rect 274036 250012 274046 250068
rect 236226 249900 236236 249956
rect 236292 249900 484988 249956
rect 485044 249900 485054 249956
rect 229842 249788 229852 249844
rect 229908 249788 495068 249844
rect 495124 249788 495134 249844
rect 236002 249676 236012 249732
rect 236068 249676 502908 249732
rect 502964 249676 502974 249732
rect 196532 249564 199052 249620
rect 199108 249564 467964 249620
rect 468020 249564 468030 249620
rect 196532 249508 196588 249564
rect 99960 249452 196588 249508
rect 223122 249452 223132 249508
rect 223188 249452 508508 249508
rect 508564 249452 508574 249508
rect 253474 249340 253484 249396
rect 253540 249340 267148 249396
rect 267204 249340 267214 249396
rect -960 248500 480 248696
rect 360322 248556 360332 248612
rect 360388 248556 378700 248612
rect 378756 248556 378766 248612
rect -960 248472 4060 248500
rect 392 248444 4060 248472
rect 4116 248444 4126 248500
rect 355730 248444 355740 248500
rect 355796 248444 376684 248500
rect 376740 248444 376750 248500
rect 355506 248332 355516 248388
rect 355572 248332 378588 248388
rect 378644 248332 378654 248388
rect 236114 248220 236124 248276
rect 236180 248220 492828 248276
rect 492884 248220 492894 248276
rect 224914 248108 224924 248164
rect 224980 248108 488348 248164
rect 488404 248108 488414 248164
rect 234882 247996 234892 248052
rect 234948 247996 498428 248052
rect 498484 247996 498494 248052
rect 226370 247884 226380 247940
rect 226436 247884 504028 247940
rect 504084 247884 504094 247940
rect 225026 247772 225036 247828
rect 225092 247772 511868 247828
rect 511924 247772 511934 247828
rect 360546 247660 360556 247716
rect 360612 247660 378924 247716
rect 378980 247660 378990 247716
rect 231858 246876 231868 246932
rect 231924 246876 231962 246932
rect 519474 246876 519484 246932
rect 519540 246876 520156 246932
rect 520212 246876 520222 246932
rect 188962 246764 188972 246820
rect 189028 246764 383068 246820
rect 383124 246764 395612 246820
rect 395668 246764 395678 246820
rect 231074 246652 231084 246708
rect 231140 246652 384748 246708
rect 384804 246652 384814 246708
rect 255266 246540 255276 246596
rect 255332 246540 270844 246596
rect 270900 246540 270910 246596
rect 254370 246428 254380 246484
rect 254436 246428 271068 246484
rect 271124 246428 271134 246484
rect 384692 246372 384748 246652
rect 227490 246316 227500 246372
rect 227556 246316 267372 246372
rect 267428 246316 267438 246372
rect 384692 246316 404012 246372
rect 404068 246316 404078 246372
rect 229730 246204 229740 246260
rect 229796 246204 487228 246260
rect 487284 246204 487294 246260
rect 228386 246092 228396 246148
rect 228452 246092 509628 246148
rect 509684 246092 509694 246148
rect 257058 245980 257068 246036
rect 257124 245980 270956 246036
rect 271012 245980 271022 246036
rect 196466 245868 196476 245924
rect 196532 245868 519484 245924
rect 519540 245868 519550 245924
rect 268706 245308 268716 245364
rect 268772 245308 272972 245364
rect 273028 245308 273038 245364
rect 595560 245028 597000 245224
rect 587122 244972 587132 245028
rect 587188 245000 597000 245028
rect 587188 244972 595672 245000
rect 355394 244636 355404 244692
rect 355460 244636 381388 244692
rect 381444 244636 381454 244692
rect 231410 244524 231420 244580
rect 231476 244524 483868 244580
rect 483924 244524 483934 244580
rect 226258 244412 226268 244468
rect 226324 244412 491708 244468
rect 491764 244412 491774 244468
rect 99960 243628 198492 243684
rect 198548 243628 198558 243684
rect 257954 243292 257964 243348
rect 258020 243292 270732 243348
rect 270788 243292 270798 243348
rect 230178 243180 230188 243236
rect 230244 243180 231644 243236
rect 231700 243180 273420 243236
rect 273476 243180 273486 243236
rect 231522 243068 231532 243124
rect 231588 243068 493948 243124
rect 494004 243068 494014 243124
rect 228162 242956 228172 243012
rect 228228 242956 499548 243012
rect 499604 242956 499614 243012
rect 228274 242844 228284 242900
rect 228340 242844 505148 242900
rect 505204 242844 505214 242900
rect 226706 242732 226716 242788
rect 226772 242732 514108 242788
rect 514164 242732 514174 242788
rect 24658 242620 24668 242676
rect 24724 242620 273196 242676
rect 273252 242620 273262 242676
rect 46162 242508 46172 242564
rect 46228 242508 230188 242564
rect 230244 242508 230254 242564
rect 40898 241948 40908 242004
rect 40964 241948 41580 242004
rect 41636 241948 41646 242004
rect 223010 241500 223020 241556
rect 223076 241500 486108 241556
rect 486164 241500 486174 241556
rect 228050 241388 228060 241444
rect 228116 241388 496188 241444
rect 496244 241388 496254 241444
rect 226594 241276 226604 241332
rect 226660 241276 501788 241332
rect 501844 241276 501854 241332
rect 223346 241164 223356 241220
rect 223412 241164 510748 241220
rect 510804 241164 510814 241220
rect 234658 241052 234668 241108
rect 234724 241052 590828 241108
rect 590884 241052 590894 241108
rect 50754 240716 50764 240772
rect 50820 240716 126812 240772
rect 126868 240716 126878 240772
rect 41458 240492 41468 240548
rect 41524 240492 44156 240548
rect 44212 240492 44222 240548
rect 54786 240492 54796 240548
rect 54852 240492 212492 240548
rect 212548 240492 212558 240548
rect 58818 240380 58828 240436
rect 58884 240380 215852 240436
rect 215908 240380 215918 240436
rect 62850 240268 62860 240324
rect 62916 240268 219212 240324
rect 219268 240268 219278 240324
rect 52770 240156 52780 240212
rect 52836 240156 60676 240212
rect 60834 240156 60844 240212
rect 60900 240156 217532 240212
rect 217588 240156 217598 240212
rect 60620 240100 60676 240156
rect 56802 240044 56812 240100
rect 56868 240044 56878 240100
rect 60620 240044 210812 240100
rect 210868 240044 210878 240100
rect 56812 239988 56868 240044
rect 56812 239932 205772 239988
rect 205828 239932 205838 239988
rect 227714 239932 227724 239988
rect 227780 239932 489468 239988
rect 489524 239932 489534 239988
rect 78978 239820 78988 239876
rect 79044 239820 217756 239876
rect 217812 239820 217822 239876
rect 230066 239820 230076 239876
rect 230132 239820 500668 239876
rect 500724 239820 500734 239876
rect 64866 239708 64876 239764
rect 64932 239708 116732 239764
rect 116788 239708 116798 239764
rect 229954 239708 229964 239764
rect 230020 239708 507388 239764
rect 507444 239708 507454 239764
rect 234434 239596 234444 239652
rect 234500 239596 512988 239652
rect 513044 239596 513054 239652
rect 235554 239484 235564 239540
rect 235620 239484 590156 239540
rect 590212 239484 590222 239540
rect 234546 239372 234556 239428
rect 234612 239372 590604 239428
rect 590660 239372 590670 239428
rect 99810 238588 99820 238644
rect 99876 238588 100212 238644
rect 100156 238532 100212 238588
rect 41010 238476 41020 238532
rect 41076 238476 46732 238532
rect 46788 238476 46798 238532
rect 74918 238476 74956 238532
rect 75012 238476 75022 238532
rect 76934 238476 76972 238532
rect 77028 238476 77038 238532
rect 91074 238476 91084 238532
rect 91140 238476 99932 238532
rect 99988 238476 99998 238532
rect 100156 238476 204092 238532
rect 204148 238476 204158 238532
rect 93090 238364 93100 238420
rect 93156 238364 93166 238420
rect 95106 238364 95116 238420
rect 95172 238364 100100 238420
rect 93100 238308 93156 238364
rect 100044 238308 100100 238364
rect 40226 238252 40236 238308
rect 40292 238252 48748 238308
rect 48804 238252 48814 238308
rect 93100 238252 99820 238308
rect 99876 238252 99886 238308
rect 100044 238252 103292 238308
rect 103348 238252 103358 238308
rect 89058 238140 89068 238196
rect 89124 238140 95452 238196
rect 95508 238140 95518 238196
rect 97122 238140 97132 238196
rect 97188 238140 106652 238196
rect 106708 238140 106718 238196
rect 87042 238028 87052 238084
rect 87108 238028 104972 238084
rect 105028 238028 105038 238084
rect 85026 237916 85036 237972
rect 85092 237916 120092 237972
rect 120148 237916 120158 237972
rect 80994 237804 81004 237860
rect 81060 237804 110012 237860
rect 110068 237804 110078 237860
rect 95442 237692 95452 237748
rect 95508 237692 100156 237748
rect 100212 237692 100222 237748
rect 219986 237692 219996 237748
rect 220052 237692 490588 237748
rect 490644 237692 490654 237748
rect 83010 237580 83020 237636
rect 83076 237580 100380 237636
rect 100436 237580 100446 237636
rect 66882 236796 66892 236852
rect 66948 236796 234556 236852
rect 234612 236796 234622 236852
rect 343970 236796 343980 236852
rect 344036 236796 536172 236852
rect 536228 236796 536238 236852
rect 223346 236684 223356 236740
rect 223412 236684 519148 236740
rect 519204 236684 519214 236740
rect 70914 236572 70924 236628
rect 70980 236572 229404 236628
rect 229460 236572 229470 236628
rect 236114 236572 236124 236628
rect 236180 236572 565292 236628
rect 565348 236572 565358 236628
rect 234770 236460 234780 236516
rect 234836 236460 590492 236516
rect 590548 236460 590558 236516
rect 234882 236348 234892 236404
rect 234948 236348 590716 236404
rect 590772 236348 590782 236404
rect 38546 236012 38556 236068
rect 38612 236012 274988 236068
rect 275044 236012 275054 236068
rect 68898 235116 68908 235172
rect 68964 235116 234332 235172
rect 234388 235116 234398 235172
rect 422482 235116 422492 235172
rect 422548 235116 423276 235172
rect 423332 235116 423342 235172
rect 72930 235004 72940 235060
rect 72996 235004 229292 235060
rect 229348 235004 229358 235060
rect 478772 234668 516292 234724
rect 478772 234612 478828 234668
rect -960 234388 480 234584
rect 423266 234556 423276 234612
rect 423332 234556 478828 234612
rect 516236 234584 516292 234668
rect 32274 234444 32284 234500
rect 32340 234444 274092 234500
rect 274148 234444 274158 234500
rect 314962 234444 314972 234500
rect 315028 234444 388892 234500
rect 388948 234444 388958 234500
rect -960 234360 207452 234388
rect 392 234332 207452 234360
rect 207508 234332 207518 234388
rect 232754 234332 232764 234388
rect 232820 234332 270620 234388
rect 270676 234332 270686 234388
rect 322466 234332 322476 234388
rect 322532 234332 407372 234388
rect 407428 234332 407438 234388
rect 318322 232876 318332 232932
rect 318388 232876 394940 232932
rect 394996 232876 395006 232932
rect 37986 232764 37996 232820
rect 38052 232764 246316 232820
rect 246372 232764 246382 232820
rect 326834 232764 326844 232820
rect 326900 232764 415100 232820
rect 415156 232764 415166 232820
rect 41010 232652 41020 232708
rect 41076 232652 376124 232708
rect 376180 232652 376190 232708
rect 590146 231980 590156 232036
rect 590212 232008 595672 232036
rect 590212 231980 597000 232008
rect 516936 231868 517468 231924
rect 517524 231868 517534 231924
rect 595560 231784 597000 231980
rect 309026 231196 309036 231252
rect 309092 231196 375452 231252
rect 375508 231196 375518 231252
rect 51986 231084 51996 231140
rect 52052 231084 249004 231140
rect 249060 231084 249070 231140
rect 320226 231084 320236 231140
rect 320292 231084 396956 231140
rect 397012 231084 397022 231140
rect 41122 230972 41132 231028
rect 41188 230972 378476 231028
rect 378532 230972 378542 231028
rect 40226 229404 40236 229460
rect 40292 229404 250796 229460
rect 250852 229404 250862 229460
rect 323474 229404 323484 229460
rect 323540 229404 403004 229460
rect 403060 229404 403070 229460
rect 15138 229292 15148 229348
rect 15204 229292 376348 229348
rect 376404 229292 376414 229348
rect 516936 229180 517580 229236
rect 517636 229180 517646 229236
rect 38434 227724 38444 227780
rect 38500 227724 247212 227780
rect 247268 227724 247278 227780
rect 320674 227724 320684 227780
rect 320740 227724 399084 227780
rect 399140 227724 399150 227780
rect 17042 227612 17052 227668
rect 17108 227612 376572 227668
rect 376628 227612 376638 227668
rect 516936 226492 517468 226548
rect 517524 226492 519372 226548
rect 519428 226492 519438 226548
rect 22754 224364 22764 224420
rect 22820 224364 244524 224420
rect 244580 224364 244590 224420
rect 325378 224364 325388 224420
rect 325444 224364 407036 224420
rect 407092 224364 407102 224420
rect 34178 224252 34188 224308
rect 34244 224252 376908 224308
rect 376964 224252 376974 224308
rect 516936 223804 517692 223860
rect 517748 223804 519372 223860
rect 519428 223804 519438 223860
rect 13234 222684 13244 222740
rect 13300 222684 242956 222740
rect 243012 222684 243022 222740
rect 323362 222684 323372 222740
rect 323428 222684 411068 222740
rect 411124 222684 411134 222740
rect 18946 222572 18956 222628
rect 19012 222572 377132 222628
rect 377188 222572 377198 222628
rect 516908 221676 517804 221732
rect 517860 221676 519148 221732
rect 519204 221676 519214 221732
rect 516908 221144 516964 221676
rect -960 220276 480 220472
rect -960 220248 12572 220276
rect 392 220220 12572 220248
rect 12628 220220 12638 220276
rect 595560 218596 597000 218792
rect 521602 218540 521612 218596
rect 521668 218568 597000 218596
rect 521668 218540 595672 218568
rect 516936 218428 519372 218484
rect 519428 218428 519438 218484
rect 232866 217756 232876 217812
rect 232932 217756 269724 217812
rect 269780 217756 269790 217812
rect 306338 217756 306348 217812
rect 306404 217756 325052 217812
rect 325108 217756 325118 217812
rect 40114 217644 40124 217700
rect 40180 217644 248108 217700
rect 248164 217644 248174 217700
rect 324258 217644 324268 217700
rect 324324 217644 413084 217700
rect 413140 217644 413150 217700
rect 20850 217532 20860 217588
rect 20916 217532 379708 217588
rect 379764 217532 379774 217588
rect 233090 216524 233100 216580
rect 233156 216524 270732 216580
rect 270788 216524 270798 216580
rect 231746 216412 231756 216468
rect 231812 216412 269388 216468
rect 269444 216412 269454 216468
rect 233202 216300 233212 216356
rect 233268 216300 274204 216356
rect 274260 216300 274270 216356
rect 229618 216188 229628 216244
rect 229684 216188 273084 216244
rect 273140 216188 273150 216244
rect 234994 216076 235004 216132
rect 235060 216076 289884 216132
rect 289940 216076 289950 216132
rect 51874 215964 51884 216020
rect 51940 215964 249900 216020
rect 249956 215964 249966 216020
rect 199042 215852 199052 215908
rect 199108 215852 464492 215908
rect 464548 215852 464558 215908
rect 516936 215740 519596 215796
rect 519652 215740 519662 215796
rect 233314 214284 233324 214340
rect 233380 214284 269388 214340
rect 269444 214284 269454 214340
rect 154914 214172 154924 214228
rect 154980 214172 200732 214228
rect 200788 214172 200798 214228
rect 219986 214172 219996 214228
rect 220052 214172 457772 214228
rect 457828 214172 457838 214228
rect 235106 213276 235116 213332
rect 235172 213276 269276 213332
rect 269332 213276 269342 213332
rect 232978 213164 232988 213220
rect 233044 213164 274092 213220
rect 274148 213164 274158 213220
rect 233426 213052 233436 213108
rect 233492 213052 274876 213108
rect 274932 213052 274942 213108
rect 516936 213052 519260 213108
rect 519316 213052 519326 213108
rect 232418 212940 232428 212996
rect 232484 212940 275772 212996
rect 275828 212940 275838 212996
rect 235778 212828 235788 212884
rect 235844 212828 307468 212884
rect 307524 212828 307534 212884
rect 235666 212716 235676 212772
rect 235732 212716 314188 212772
rect 314244 212716 314254 212772
rect 235890 212604 235900 212660
rect 235956 212604 320908 212660
rect 320964 212604 320974 212660
rect 26562 212492 26572 212548
rect 26628 212492 376236 212548
rect 376292 212492 376302 212548
rect 237794 211484 237804 211540
rect 237860 211484 274652 211540
rect 274708 211484 274718 211540
rect 234994 211372 235004 211428
rect 235060 211372 269836 211428
rect 269892 211372 269902 211428
rect 231186 211260 231196 211316
rect 231252 211260 272412 211316
rect 272468 211260 272478 211316
rect 229842 211148 229852 211204
rect 229908 211148 269500 211204
rect 269556 211148 269566 211204
rect 226706 211036 226716 211092
rect 226772 211036 269836 211092
rect 269892 211036 269902 211092
rect 237682 210924 237692 210980
rect 237748 210924 286412 210980
rect 286468 210924 286478 210980
rect 30370 210812 30380 210868
rect 30436 210812 245420 210868
rect 245476 210812 245486 210868
rect 331874 210812 331884 210868
rect 331940 210812 417116 210868
rect 417172 210812 417182 210868
rect 516908 210812 519484 210868
rect 519540 210812 587132 210868
rect 587188 210812 587198 210868
rect 269490 210700 269500 210756
rect 269556 210700 272748 210756
rect 272804 210700 272814 210756
rect 516908 210392 516964 210812
rect 50306 210140 50316 210196
rect 50372 210140 272748 210196
rect 272804 210140 272814 210196
rect 49522 210028 49532 210084
rect 49588 210028 272524 210084
rect 272580 210028 272590 210084
rect 234434 209916 234444 209972
rect 234500 209916 269556 209972
rect 231298 209804 231308 209860
rect 231364 209804 269332 209860
rect 231410 209692 231420 209748
rect 231476 209692 269220 209748
rect 229954 209580 229964 209636
rect 230020 209580 269108 209636
rect 228386 209468 228396 209524
rect 228452 209468 268212 209524
rect 226594 209356 226604 209412
rect 226660 209356 267148 209412
rect 267092 209076 267148 209356
rect 268156 209188 268212 209468
rect 269052 209300 269108 209580
rect 269164 209524 269220 209692
rect 269276 209636 269332 209804
rect 269500 209748 269556 209916
rect 272374 209804 272412 209860
rect 272468 209804 272478 209860
rect 269490 209692 269500 209748
rect 269556 209692 269566 209748
rect 269276 209580 272916 209636
rect 272860 209524 272916 209580
rect 269164 209468 272692 209524
rect 272850 209468 272860 209524
rect 272916 209468 272926 209524
rect 272636 209412 272692 209468
rect 272626 209356 272636 209412
rect 272692 209356 272702 209412
rect 269052 209244 273196 209300
rect 273252 209244 273262 209300
rect 268156 209132 273084 209188
rect 273140 209132 273150 209188
rect 267092 209020 272524 209076
rect 272580 209020 272590 209076
rect 4162 208684 4172 208740
rect 4228 208684 272300 208740
rect 272356 208684 272366 208740
rect 269826 207900 269836 207956
rect 269892 207900 269902 207956
rect 269836 207032 269892 207900
rect 516936 207676 519148 207732
rect 519204 207676 519214 207732
rect 464482 206668 464492 206724
rect 464548 206668 465948 206724
rect 466004 206668 466014 206724
rect 392 206360 4172 206388
rect -960 206332 4172 206360
rect 4228 206332 4238 206388
rect -960 206136 480 206332
rect 321906 205772 321916 205828
rect 321972 205772 400988 205828
rect 401044 205772 401054 205828
rect 595560 205380 597000 205576
rect 519138 205324 519148 205380
rect 519204 205352 597000 205380
rect 519204 205324 595672 205352
rect 516936 204988 519148 205044
rect 519204 204988 519214 205044
rect 269490 204652 269500 204708
rect 269556 204652 269566 204708
rect 269500 204120 269556 204652
rect 314402 204092 314412 204148
rect 314468 204092 390908 204148
rect 390964 204092 390974 204148
rect 516236 201684 516292 202328
rect 516226 201628 516236 201684
rect 516292 201628 516302 201684
rect 269826 201516 269836 201572
rect 269892 201516 269902 201572
rect 269836 201208 269892 201516
rect 472994 200844 473004 200900
rect 473060 200844 517804 200900
rect 517860 200844 517870 200900
rect 356962 200620 356972 200676
rect 357028 200620 553644 200676
rect 553700 200620 553710 200676
rect 345202 200508 345212 200564
rect 345268 200508 534828 200564
rect 534884 200508 534894 200564
rect 467842 200396 467852 200452
rect 467908 200396 511644 200452
rect 511700 200396 511710 200452
rect 461122 200284 461132 200340
rect 461188 200284 505372 200340
rect 505428 200284 505438 200340
rect 507938 200284 507948 200340
rect 508004 200284 517580 200340
rect 517636 200284 517646 200340
rect 457762 200172 457772 200228
rect 457828 200172 508508 200228
rect 508564 200172 508574 200228
rect 383954 200060 383964 200116
rect 384020 200060 488124 200116
rect 488180 200060 488190 200116
rect 415762 199948 415772 200004
rect 415828 199948 512428 200004
rect 512484 199948 512494 200004
rect 414082 199836 414092 199892
rect 414148 199836 514892 199892
rect 514948 199836 514958 199892
rect 417442 199724 417452 199780
rect 417508 199724 510076 199780
rect 510132 199724 510142 199780
rect 514052 199724 519148 199780
rect 519204 199724 519214 199780
rect 514052 199668 514108 199724
rect 465938 199612 465948 199668
rect 466004 199612 466284 199668
rect 466340 199612 514108 199668
rect 467954 199500 467964 199556
rect 468020 199500 519484 199556
rect 519540 199500 519550 199556
rect 459442 199388 459452 199444
rect 459508 199388 506492 199444
rect 506548 199388 506940 199444
rect 506996 199388 507006 199444
rect 510290 199388 510300 199444
rect 510356 199388 516236 199444
rect 516292 199388 516302 199444
rect 474674 199276 474684 199332
rect 474740 199276 517692 199332
rect 517748 199276 517758 199332
rect 330530 199164 330540 199220
rect 330596 199164 513436 199220
rect 513492 199164 513502 199220
rect 344866 199052 344876 199108
rect 344932 199052 533372 199108
rect 533428 199052 533438 199108
rect 462802 198940 462812 198996
rect 462868 198940 503132 198996
rect 503188 198940 503804 198996
rect 503860 198940 503870 198996
rect 269864 198268 273196 198324
rect 273252 198268 273262 198324
rect 479602 198156 479612 198212
rect 479668 198156 494396 198212
rect 494452 198156 494462 198212
rect 497522 198156 497532 198212
rect 497588 198156 497644 198212
rect 497700 198156 497710 198212
rect 499062 198156 499100 198212
rect 499156 198156 499166 198212
rect 502198 198156 502236 198212
rect 502292 198156 502302 198212
rect 481282 198044 481292 198100
rect 481348 198044 500668 198100
rect 500724 198044 500734 198100
rect 477922 197932 477932 197988
rect 477988 197932 495964 197988
rect 496020 197932 496030 197988
rect 398962 197820 398972 197876
rect 399028 197820 486556 197876
rect 486612 197820 486622 197876
rect 397282 197708 397292 197764
rect 397348 197708 483420 197764
rect 483476 197708 483486 197764
rect 474562 197596 474572 197652
rect 474628 197596 491260 197652
rect 491316 197596 491326 197652
rect 472882 197484 472892 197540
rect 472948 197484 492828 197540
rect 492884 197484 492894 197540
rect 305442 197372 305452 197428
rect 305508 197372 370748 197428
rect 370804 197372 370814 197428
rect 400642 197372 400652 197428
rect 400708 197372 489692 197428
rect 489748 197372 489758 197428
rect 387202 197260 387212 197316
rect 387268 197260 484988 197316
rect 485044 197260 485054 197316
rect 385522 197148 385532 197204
rect 385588 197148 481852 197204
rect 481908 197148 481918 197204
rect 453506 195916 453516 195972
rect 453572 195916 482412 195972
rect 482468 195916 482478 195972
rect 471650 195804 471660 195860
rect 471716 195804 519372 195860
rect 519428 195804 519438 195860
rect 349346 195692 349356 195748
rect 349412 195692 544236 195748
rect 544292 195692 544302 195748
rect 269864 195356 273084 195412
rect 273140 195356 273150 195412
rect 326946 194124 326956 194180
rect 327012 194124 506828 194180
rect 506884 194124 506894 194180
rect 352930 194012 352940 194068
rect 352996 194012 549612 194068
rect 549668 194012 549678 194068
rect 269864 192444 272524 192500
rect 272580 192444 272590 192500
rect 335906 192444 335916 192500
rect 335972 192444 515004 192500
rect 515060 192444 515070 192500
rect 309922 192332 309932 192388
rect 309988 192332 331884 192388
rect 331940 192332 331950 192388
rect 353826 192332 353836 192388
rect 353892 192332 547148 192388
rect 547204 192332 547214 192388
rect 590818 192332 590828 192388
rect 590884 192360 595672 192388
rect 590884 192332 597000 192360
rect -960 192052 480 192248
rect 595560 192136 597000 192332
rect -960 192024 14252 192052
rect 392 191996 14252 192024
rect 14308 191996 14318 192052
rect 269864 189532 272412 189588
rect 272468 189532 272478 189588
rect 331426 188972 331436 189028
rect 331492 188972 517356 189028
rect 517412 188972 517422 189028
rect 339490 187404 339500 187460
rect 339556 187404 529452 187460
rect 529508 187404 529518 187460
rect 354722 187292 354732 187348
rect 354788 187292 552300 187348
rect 552356 187292 552366 187348
rect 269864 186620 272860 186676
rect 272916 186620 272926 186676
rect 341282 185612 341292 185668
rect 341348 185612 526652 185668
rect 526708 185612 526718 185668
rect 269864 183708 272748 183764
rect 272804 183708 272814 183764
rect 327842 182364 327852 182420
rect 327908 182364 511980 182420
rect 512036 182364 512046 182420
rect 359314 182252 359324 182308
rect 359380 182252 559468 182308
rect 559524 182252 559534 182308
rect 269864 180796 272412 180852
rect 272468 180796 272478 180852
rect 345762 180572 345772 180628
rect 345828 180572 538860 180628
rect 538916 180572 538926 180628
rect 335122 179004 335132 179060
rect 335188 179004 521388 179060
rect 521444 179004 521454 179060
rect 595560 178948 597000 179144
rect 380482 178892 380492 178948
rect 380548 178920 597000 178948
rect 380548 178892 595672 178920
rect -960 177940 480 178136
rect -960 177912 27804 177940
rect 392 177884 27804 177912
rect 27860 177884 27870 177940
rect 269864 177884 275772 177940
rect 275828 177884 275838 177940
rect 350242 177212 350252 177268
rect 350308 177212 545580 177268
rect 545636 177212 545646 177268
rect 376002 175644 376012 175700
rect 376068 175644 562828 175700
rect 562884 175644 562894 175700
rect 351138 175532 351148 175588
rect 351204 175532 541772 175588
rect 541828 175532 541838 175588
rect 269864 174972 274204 175028
rect 274260 174972 274270 175028
rect 352034 173852 352044 173908
rect 352100 173852 548268 173908
rect 548324 173852 548334 173908
rect 269378 172060 269388 172116
rect 269444 172060 269454 172116
rect 328738 170604 328748 170660
rect 328804 170604 513324 170660
rect 513380 170604 513390 170660
rect 370402 170492 370412 170548
rect 370468 170492 563164 170548
rect 563220 170492 563230 170548
rect 269864 169148 270732 169204
rect 270788 169148 270798 169204
rect 372082 168924 372092 168980
rect 372148 168924 562940 168980
rect 562996 168924 563006 168980
rect 342178 168812 342188 168868
rect 342244 168812 533484 168868
rect 533540 168812 533550 168868
rect 362786 167132 362796 167188
rect 362852 167132 566188 167188
rect 566244 167132 566254 167188
rect 269864 166236 273980 166292
rect 274036 166236 274046 166292
rect 595560 165704 597000 165928
rect 392 164024 4172 164052
rect -960 163996 4172 164024
rect 4228 163996 4238 164052
rect -960 163800 480 163996
rect 340386 163884 340396 163940
rect 340452 163884 530796 163940
rect 530852 163884 530862 163940
rect 357410 163772 357420 163828
rect 357476 163772 559580 163828
rect 559636 163772 559646 163828
rect 269864 163324 273868 163380
rect 273924 163324 273934 163380
rect 468962 162316 468972 162372
rect 469028 162316 519260 162372
rect 519316 162316 519326 162372
rect 333442 162204 333452 162260
rect 333508 162204 518700 162260
rect 518756 162204 518766 162260
rect 358306 162092 358316 162148
rect 358372 162092 559804 162148
rect 559860 162092 559870 162148
rect 475682 160972 475692 161028
rect 475748 160972 517468 161028
rect 517524 160972 517534 161028
rect 470306 160860 470316 160916
rect 470372 160860 519596 160916
rect 519652 160860 519662 160916
rect 310930 160748 310940 160804
rect 310996 160748 375564 160804
rect 375620 160748 494508 160804
rect 494564 160748 494574 160804
rect 307346 160636 307356 160692
rect 307412 160636 373100 160692
rect 373156 160636 493164 160692
rect 493220 160636 493230 160692
rect 356514 160524 356524 160580
rect 356580 160524 559692 160580
rect 559748 160524 559758 160580
rect 269714 160412 269724 160468
rect 269780 160412 269790 160468
rect 360098 160412 360108 160468
rect 360164 160412 564508 160468
rect 564564 160412 564574 160468
rect 329634 158956 329644 159012
rect 329700 158956 514668 159012
rect 514724 158956 514734 159012
rect 514882 158956 514892 159012
rect 514948 158956 561708 159012
rect 561764 158956 561774 159012
rect 333218 158844 333228 158900
rect 333284 158844 520044 158900
rect 520100 158844 520110 158900
rect 335010 158732 335020 158788
rect 335076 158732 522732 158788
rect 522788 158732 522798 158788
rect 269864 157500 270620 157556
rect 270676 157500 270686 157556
rect 346658 157276 346668 157332
rect 346724 157276 540204 157332
rect 540260 157276 540270 157332
rect 347554 157164 347564 157220
rect 347620 157164 541548 157220
rect 541604 157164 541614 157220
rect 348450 157052 348460 157108
rect 348516 157052 542892 157108
rect 542948 157052 542958 157108
rect 296482 156604 296492 156660
rect 296548 156604 491820 156660
rect 491876 156604 491886 156660
rect 283826 156492 283836 156548
rect 283892 156492 487788 156548
rect 487844 156492 487854 156548
rect 275314 156380 275324 156436
rect 275380 156380 479724 156436
rect 479780 156380 479790 156436
rect 274642 156268 274652 156324
rect 274708 156268 275436 156324
rect 275492 156268 483756 156324
rect 483812 156268 483822 156324
rect 336914 155708 336924 155764
rect 336980 155708 525420 155764
rect 525476 155708 525486 155764
rect 337698 155596 337708 155652
rect 337764 155596 526764 155652
rect 526820 155596 526830 155652
rect 338594 155484 338604 155540
rect 338660 155484 528108 155540
rect 528164 155484 528174 155540
rect 273298 155372 273308 155428
rect 273364 155372 273980 155428
rect 274036 155372 486444 155428
rect 486500 155372 486510 155428
rect 513202 155372 513212 155428
rect 513268 155372 561372 155428
rect 561428 155372 561438 155428
rect 295138 154700 295148 154756
rect 295204 154700 490476 154756
rect 490532 154700 490542 154756
rect 269864 154588 274092 154644
rect 274148 154588 274158 154644
rect 293916 154588 489132 154644
rect 489188 154588 489198 154644
rect 293916 154532 293972 154588
rect 273634 154476 273644 154532
rect 273700 154476 275436 154532
rect 275492 154476 275502 154532
rect 286402 154476 286412 154532
rect 286468 154476 293972 154532
rect 308242 154476 308252 154532
rect 308308 154476 310940 154532
rect 310996 154476 311006 154532
rect 367042 154476 367052 154532
rect 367108 154476 375900 154532
rect 375956 154476 506660 154532
rect 506818 154476 506828 154532
rect 506884 154476 510636 154532
rect 510692 154476 510702 154532
rect 513426 154476 513436 154532
rect 513492 154476 516012 154532
rect 516068 154476 516078 154532
rect 526642 154476 526652 154532
rect 526708 154476 532140 154532
rect 532196 154476 532206 154532
rect 533362 154476 533372 154532
rect 533428 154476 537516 154532
rect 537572 154476 537582 154532
rect 541762 154476 541772 154532
rect 541828 154476 546924 154532
rect 546980 154476 546990 154532
rect 547138 154476 547148 154532
rect 547204 154476 550956 154532
rect 551012 154476 551022 154532
rect 506604 154420 506660 154476
rect 272738 154364 272748 154420
rect 272804 154364 272814 154420
rect 273186 154364 273196 154420
rect 273252 154364 275324 154420
rect 275380 154364 275390 154420
rect 278852 154364 367052 154420
rect 367108 154364 367118 154420
rect 376114 154364 376124 154420
rect 376180 154364 502404 154420
rect 506604 154364 510076 154420
rect 510132 154364 510142 154420
rect 514994 154364 515004 154420
rect 515060 154364 524076 154420
rect 524132 154364 524142 154420
rect 272748 154308 272804 154364
rect 278852 154308 278908 154364
rect 502348 154308 502404 154364
rect 272748 154252 278908 154308
rect 291554 154252 291564 154308
rect 291620 154252 295148 154308
rect 295204 154252 295214 154308
rect 356962 154252 356972 154308
rect 357028 154252 375676 154308
rect 375732 154252 376236 154308
rect 376292 154252 376302 154308
rect 502348 154252 503860 154308
rect 503804 154196 503860 154252
rect 371298 154140 371308 154196
rect 371364 154140 372316 154196
rect 372372 154140 497196 154196
rect 497252 154140 497262 154196
rect 503804 154140 507948 154196
rect 508004 154140 508014 154196
rect 272178 154028 272188 154084
rect 272244 154028 273756 154084
rect 273812 154028 273822 154084
rect 361172 154028 372988 154084
rect 373044 154028 498540 154084
rect 498596 154028 498606 154084
rect 361172 153860 361228 154028
rect 367042 153916 367052 153972
rect 367108 153916 375452 153972
rect 375508 153916 503916 153972
rect 503972 153916 503982 153972
rect 323362 153804 323372 153860
rect 323428 153804 361228 153860
rect 376002 153804 376012 153860
rect 376068 153804 505260 153860
rect 505316 153804 505326 153860
rect 318322 153692 318332 153748
rect 318388 153692 371308 153748
rect 371364 153692 371374 153748
rect 376226 153692 376236 153748
rect 376292 153692 506604 153748
rect 506660 153692 506670 153748
rect 362002 153580 362012 153636
rect 362068 153580 376124 153636
rect 376180 153580 376190 153636
rect 272514 153468 272524 153524
rect 272580 153468 375564 153524
rect 375620 153468 376012 153524
rect 376068 153468 376078 153524
rect 273410 153132 273420 153188
rect 273476 153132 502572 153188
rect 502628 153132 502638 153188
rect 272962 153020 272972 153076
rect 273028 153020 499884 153076
rect 499940 153020 499950 153076
rect 282156 152908 283836 152964
rect 283892 152908 283902 152964
rect 303986 152908 303996 152964
rect 304052 152908 307356 152964
rect 307412 152908 307422 152964
rect 495814 152908 495852 152964
rect 495908 152908 495918 152964
rect 501302 152908 501340 152964
rect 501396 152908 501406 152964
rect 282156 152852 282212 152908
rect 274642 152796 274652 152852
rect 274708 152796 282212 152852
rect 590706 152684 590716 152740
rect 590772 152712 595672 152740
rect 590772 152684 597000 152712
rect 595560 152488 597000 152684
rect 523282 152348 523292 152404
rect 523348 152348 563052 152404
rect 563108 152348 563118 152404
rect 511634 152236 511644 152292
rect 511700 152236 561596 152292
rect 561652 152236 561662 152292
rect 276322 152124 276332 152180
rect 276388 152124 476252 152180
rect 476308 152124 476318 152180
rect 509842 152124 509852 152180
rect 509908 152124 561148 152180
rect 561204 152124 561214 152180
rect 393922 152012 393932 152068
rect 393988 152012 456988 152068
rect 457044 152012 457054 152068
rect 503122 152012 503132 152068
rect 503188 152012 566300 152068
rect 566356 152012 566366 152068
rect 456082 151900 456092 151956
rect 456148 151900 467852 151956
rect 467908 151900 467918 151956
rect 456306 151788 456316 151844
rect 456372 151788 475692 151844
rect 475748 151788 475758 151844
rect 269864 151676 273868 151732
rect 273924 151676 273934 151732
rect 451042 151676 451052 151732
rect 451108 151676 473004 151732
rect 473060 151676 473070 151732
rect 437602 151564 437612 151620
rect 437668 151564 474684 151620
rect 474740 151564 474750 151620
rect 357746 151452 357756 151508
rect 357812 151452 485100 151508
rect 485156 151452 485166 151508
rect 309922 151340 309932 151396
rect 309988 151340 480508 151396
rect 480564 151340 480574 151396
rect 459442 151228 459452 151284
rect 459508 151228 470316 151284
rect 470372 151228 470382 151284
rect 548482 150780 548492 150836
rect 548548 150780 563388 150836
rect 563444 150780 563454 150836
rect 506482 150668 506492 150724
rect 506548 150668 564732 150724
rect 564788 150668 564798 150724
rect 310034 150556 310044 150612
rect 310100 150556 368732 150612
rect 368788 150556 368798 150612
rect 412402 150556 412412 150612
rect 412468 150556 563276 150612
rect 563332 150556 563342 150612
rect 368162 150444 368172 150500
rect 368228 150444 559916 150500
rect 559972 150444 559982 150500
rect 293122 150332 293132 150388
rect 293188 150332 303996 150388
rect 304052 150332 304062 150388
rect 365474 150332 365484 150388
rect 365540 150332 564620 150388
rect 564676 150332 564686 150388
rect 392 149912 7532 149940
rect -960 149884 7532 149912
rect 7588 149884 7598 149940
rect -960 149688 480 149884
rect 468962 149660 468972 149716
rect 469028 149660 469038 149716
rect 449362 149436 449372 149492
rect 449428 149436 465500 149492
rect 465556 149436 465566 149492
rect 465714 149436 465724 149492
rect 465780 149436 465790 149492
rect 465724 149380 465780 149436
rect 459890 149324 459900 149380
rect 459956 149324 465780 149380
rect 468972 149268 469028 149660
rect 508834 149548 508844 149604
rect 508900 149548 508910 149604
rect 471874 149436 471884 149492
rect 471940 149436 471950 149492
rect 505474 149436 505484 149492
rect 505540 149436 505550 149492
rect 471884 149268 471940 149436
rect 452722 149212 452732 149268
rect 452788 149212 469028 149268
rect 471650 149212 471660 149268
rect 471716 149212 471940 149268
rect 471660 149156 471716 149212
rect 465490 149100 465500 149156
rect 465556 149100 471716 149156
rect 505484 149156 505540 149436
rect 508844 149268 508900 149548
rect 509730 149436 509740 149492
rect 509796 149436 561260 149492
rect 561316 149436 561326 149492
rect 508844 149212 561484 149268
rect 561540 149212 561550 149268
rect 505484 149100 509740 149156
rect 509796 149100 509806 149156
rect 269266 148764 269276 148820
rect 269332 148764 269342 148820
rect 454402 148652 454412 148708
rect 454468 148652 459900 148708
rect 459956 148652 459966 148708
rect 540082 148652 540092 148708
rect 540148 148652 563164 148708
rect 563220 148652 563230 148708
rect 456978 148540 456988 148596
rect 457044 148540 460068 148596
rect 460012 147896 460068 148540
rect 555202 148092 555212 148148
rect 555268 148092 563052 148148
rect 563108 148092 563118 148148
rect 556882 147980 556892 148036
rect 556948 147980 562940 148036
rect 562996 147980 563006 148036
rect 269836 145348 269892 145880
rect 269836 145292 271180 145348
rect 271236 145292 367052 145348
rect 367108 145292 367118 145348
rect 390562 145068 390572 145124
rect 390628 145068 459396 145124
rect 459340 145012 460040 145068
rect 269528 142968 362012 142996
rect 269500 142940 362012 142968
rect 362068 142940 362078 142996
rect 559944 142940 563164 142996
rect 563220 142940 563230 142996
rect 269500 142884 269556 142940
rect 269490 142828 269500 142884
rect 269556 142828 269566 142884
rect 388882 142156 388892 142212
rect 388948 142156 459396 142212
rect 459340 142100 460040 142156
rect 320002 141932 320012 141988
rect 320068 141932 386876 141988
rect 386932 141932 386942 141988
rect 559944 141372 561708 141428
rect 561764 141372 561774 141428
rect 278852 141036 356972 141092
rect 357028 141036 357038 141092
rect 278852 140756 278908 141036
rect 269836 140700 272300 140756
rect 272356 140700 278908 140756
rect 269836 140056 269892 140700
rect 559944 139804 561372 139860
rect 561428 139804 561438 139860
rect 595560 139300 597000 139496
rect 380482 139244 380492 139300
rect 380548 139244 459396 139300
rect 578722 139244 578732 139300
rect 578788 139272 597000 139300
rect 578788 139244 595672 139272
rect 459340 139188 460040 139244
rect 315298 138572 315308 138628
rect 315364 138572 392924 138628
rect 392980 138572 392990 138628
rect 559944 138236 561596 138292
rect 561652 138236 561662 138292
rect 269864 137116 272524 137172
rect 272580 137116 272590 137172
rect 559944 136668 561148 136724
rect 561204 136668 561214 136724
rect 387202 136332 387212 136388
rect 387268 136332 459396 136388
rect 459340 136276 460040 136332
rect 273718 136108 273756 136164
rect 273812 136108 273822 136164
rect -960 135604 480 135800
rect -960 135576 32732 135604
rect 392 135548 32732 135576
rect 32788 135548 32798 135604
rect 559944 135100 561484 135156
rect 561540 135100 561550 135156
rect 269864 134204 272748 134260
rect 272804 134204 272814 134260
rect 304882 133532 304892 133588
rect 304948 133532 362684 133588
rect 362740 133532 362750 133588
rect 559944 133532 564732 133588
rect 564788 133532 564798 133588
rect 385522 133420 385532 133476
rect 385588 133420 459396 133476
rect 459340 133364 460040 133420
rect 559944 131964 561260 132020
rect 561316 131964 561326 132020
rect 311714 131852 311724 131908
rect 311780 131852 384860 131908
rect 384916 131852 384926 131908
rect 269864 131292 273420 131348
rect 273476 131292 273486 131348
rect 451042 130508 451052 130564
rect 451108 130508 459396 130564
rect 459340 130452 460040 130508
rect 559944 130396 566300 130452
rect 566356 130396 566366 130452
rect 559944 128828 563388 128884
rect 563444 128828 563454 128884
rect 321682 128492 321692 128548
rect 321748 128492 382844 128548
rect 382900 128492 382910 128548
rect 395602 128492 395612 128548
rect 395668 128492 457884 128548
rect 457940 128492 457950 128548
rect 269864 128380 273756 128436
rect 273812 128380 273822 128436
rect 382162 127596 382172 127652
rect 382228 127596 459396 127652
rect 559906 127596 559916 127652
rect 559972 127596 559982 127652
rect 459340 127540 460040 127596
rect 559916 127288 559972 127596
rect 307234 126924 307244 126980
rect 307300 126924 374780 126980
rect 374836 126924 374846 126980
rect 308130 126812 308140 126868
rect 308196 126812 376796 126868
rect 376852 126812 376862 126868
rect 595560 126056 597000 126280
rect 559944 125692 563276 125748
rect 563332 125692 563342 125748
rect 269864 125468 272972 125524
rect 273028 125468 273038 125524
rect 302754 125356 302764 125412
rect 302820 125356 364700 125412
rect 364756 125356 364766 125412
rect 303650 125244 303660 125300
rect 303716 125244 366716 125300
rect 366772 125244 366782 125300
rect 317986 125132 317996 125188
rect 318052 125132 398972 125188
rect 399028 125132 399038 125188
rect 392242 124684 392252 124740
rect 392308 124684 459396 124740
rect 459340 124628 460040 124684
rect 407362 124236 407372 124292
rect 407428 124236 409052 124292
rect 409108 124236 409118 124292
rect 559944 124124 562828 124180
rect 562884 124124 562894 124180
rect 325042 123676 325052 123732
rect 325108 123676 372764 123732
rect 372820 123676 372830 123732
rect 331874 123564 331884 123620
rect 331940 123564 380828 123620
rect 380884 123564 380894 123620
rect 274642 123452 274652 123508
rect 274708 123452 379036 123508
rect 379092 123452 379102 123508
rect 375442 122668 375452 122724
rect 375508 122668 378812 122724
rect 378868 122668 378878 122724
rect 399074 122668 399084 122724
rect 399140 122668 405020 122724
rect 405076 122668 405086 122724
rect 269864 122556 323372 122612
rect 323428 122556 323438 122612
rect 559944 122556 564620 122612
rect 564676 122556 564686 122612
rect 560242 122444 560252 122500
rect 560308 122444 562828 122500
rect 562884 122444 562894 122500
rect 274866 121772 274876 121828
rect 274932 121772 378700 121828
rect 378756 121772 378766 121828
rect 383842 121772 383852 121828
rect 383908 121772 459396 121828
rect 459340 121716 460040 121772
rect 392 121688 4172 121716
rect -960 121660 4172 121688
rect 4228 121660 4238 121716
rect -960 121464 480 121660
rect 559944 120988 563052 121044
rect 563108 120988 563118 121044
rect 560242 120876 560252 120932
rect 560308 120876 562828 120932
rect 562884 120876 562894 120932
rect 357634 120204 357644 120260
rect 357700 120204 377244 120260
rect 377300 120204 377310 120260
rect 272962 120092 272972 120148
rect 273028 120092 378924 120148
rect 378980 120092 378990 120148
rect 404002 120092 404012 120148
rect 404068 120092 457996 120148
rect 458052 120092 458062 120148
rect 269864 119644 318332 119700
rect 318388 119644 318398 119700
rect 559944 119420 562940 119476
rect 562996 119420 563006 119476
rect 456082 118860 456092 118916
rect 456148 118860 459396 118916
rect 459340 118804 460040 118860
rect 559944 117852 566188 117908
rect 566244 117852 566254 117908
rect 269864 116732 313404 116788
rect 313460 116732 313470 116788
rect 559944 116284 562828 116340
rect 562884 116284 562894 116340
rect 419346 116060 419356 116116
rect 419412 116060 441084 116116
rect 441140 116060 441150 116116
rect 459340 115892 460040 115948
rect 442642 115836 442652 115892
rect 442708 115836 459396 115892
rect 559944 114716 564508 114772
rect 564564 114716 564574 114772
rect 269864 113820 308252 113876
rect 308308 113820 308318 113876
rect 559458 113708 559468 113764
rect 559524 113708 559534 113764
rect 559468 113176 559524 113708
rect 437602 113036 437612 113092
rect 437668 113036 459396 113092
rect 590594 113036 590604 113092
rect 590660 113064 595672 113092
rect 590660 113036 597000 113064
rect 459340 112980 460040 113036
rect 595560 112840 597000 113036
rect 559794 112140 559804 112196
rect 559860 112140 559870 112196
rect 559804 111608 559860 112140
rect 269864 110908 293132 110964
rect 293188 110908 293198 110964
rect 559570 110572 559580 110628
rect 559636 110572 559646 110628
rect 434242 110124 434252 110180
rect 434308 110124 459396 110180
rect 459340 110068 460040 110124
rect 559580 110040 559636 110572
rect 273074 109116 273084 109172
rect 273140 109116 337708 109172
rect 419944 109116 423276 109172
rect 423332 109116 427644 109172
rect 427700 109116 427710 109172
rect 559682 109116 559692 109172
rect 559748 109116 559758 109172
rect 337652 108948 337708 109116
rect 337652 108892 357756 108948
rect 357812 108892 360164 108948
rect 360108 108248 360164 108892
rect 559692 108472 559748 109116
rect 269864 107996 296492 108052
rect 296548 107996 296558 108052
rect -960 107380 480 107576
rect -960 107352 31052 107380
rect 392 107324 31052 107352
rect 31108 107324 31118 107380
rect 432562 107212 432572 107268
rect 432628 107212 459396 107268
rect 459340 107156 460040 107212
rect 559944 106876 562828 106932
rect 562884 106876 562894 106932
rect 559944 105308 571564 105364
rect 571620 105308 571630 105364
rect 269864 105084 291564 105140
rect 291620 105084 291630 105140
rect 430882 104300 430892 104356
rect 430948 104300 459396 104356
rect 459340 104244 460040 104300
rect 559944 103740 573132 103796
rect 573188 103740 573198 103796
rect 269864 102172 286412 102228
rect 286468 102172 286478 102228
rect 419916 101668 419972 102200
rect 559944 102172 574700 102228
rect 574756 102172 574766 102228
rect 419916 101612 456316 101668
rect 456372 101612 456382 101668
rect 419916 101556 419972 101612
rect 419916 101500 420028 101556
rect 420084 101500 420094 101556
rect 427522 101388 427532 101444
rect 427588 101388 459396 101444
rect 459340 101332 460040 101388
rect 559944 100604 568204 100660
rect 568260 100604 568270 100660
rect 585442 99820 585452 99876
rect 585508 99848 595672 99876
rect 585508 99820 597000 99848
rect 595560 99624 597000 99820
rect 269864 99260 274764 99316
rect 274820 99260 274830 99316
rect 559944 99036 573020 99092
rect 573076 99036 573086 99092
rect 429202 98476 429212 98532
rect 429268 98476 459396 98532
rect 459340 98420 460040 98476
rect 559944 97468 564956 97524
rect 565012 97468 565022 97524
rect 269864 96348 273308 96404
rect 273364 96348 273374 96404
rect 559944 95900 571452 95956
rect 571508 95900 571518 95956
rect 454402 95564 454412 95620
rect 454468 95564 459396 95620
rect 459340 95508 460040 95564
rect 419916 94948 419972 95256
rect 419916 94892 420140 94948
rect 420196 94892 437612 94948
rect 437668 94892 437678 94948
rect 559944 94332 572908 94388
rect 572964 94332 572974 94388
rect -960 93268 480 93464
rect 269864 93436 273084 93492
rect 273140 93436 273150 93492
rect -960 93240 29372 93268
rect 392 93212 29372 93240
rect 29428 93212 29438 93268
rect 559944 92764 569772 92820
rect 569828 92764 569838 92820
rect 425954 92652 425964 92708
rect 426020 92652 459396 92708
rect 459340 92596 460040 92652
rect 559944 91196 566524 91252
rect 566580 91196 566590 91252
rect 269864 90524 273644 90580
rect 273700 90524 273710 90580
rect 424162 89740 424172 89796
rect 424228 89740 459396 89796
rect 459340 89684 460040 89740
rect 559944 89628 571340 89684
rect 571396 89628 571406 89684
rect 419916 88228 419972 88312
rect 269378 88172 269388 88228
rect 269444 88172 269454 88228
rect 419916 88172 420252 88228
rect 420308 88172 451052 88228
rect 451108 88172 451118 88228
rect 269388 87640 269444 88172
rect 559944 88060 571228 88116
rect 571284 88060 571294 88116
rect 420802 86828 420812 86884
rect 420868 86828 459396 86884
rect 459340 86772 460040 86828
rect 559944 86492 569548 86548
rect 569604 86492 569614 86548
rect 595560 86408 597000 86632
rect 357634 84924 357644 84980
rect 357700 84924 360136 84980
rect 559944 84924 569660 84980
rect 569716 84924 569726 84980
rect 269864 84700 309932 84756
rect 309988 84700 309998 84756
rect 457874 83916 457884 83972
rect 457940 83916 459396 83972
rect 459340 83860 460040 83916
rect 559944 83356 566412 83412
rect 566468 83356 566478 83412
rect 269864 81788 273196 81844
rect 273252 81788 273262 81844
rect 559944 81788 564844 81844
rect 564900 81788 564910 81844
rect 419916 81452 421708 81508
rect 421764 81452 449372 81508
rect 449428 81452 449438 81508
rect 419916 81368 419972 81452
rect 457986 81004 457996 81060
rect 458052 81004 459396 81060
rect 459340 80948 460040 81004
rect 559944 80220 568092 80276
rect 568148 80220 568158 80276
rect -960 79156 480 79352
rect 269266 79212 269276 79268
rect 269332 79212 269342 79268
rect -960 79128 4172 79156
rect 392 79100 4172 79128
rect 4228 79100 4238 79156
rect 269276 78904 269332 79212
rect 559944 78652 567980 78708
rect 568036 78652 568046 78708
rect 452722 78092 452732 78148
rect 452788 78092 459396 78148
rect 459340 78036 460040 78092
rect 559944 77084 566188 77140
rect 566244 77084 566254 77140
rect 269864 75964 276332 76020
rect 276388 75964 276398 76020
rect 559944 75516 564732 75572
rect 564788 75516 564798 75572
rect 440962 75180 440972 75236
rect 441028 75180 459396 75236
rect 459340 75124 460040 75180
rect 419916 74732 421820 74788
rect 421876 74732 459452 74788
rect 459508 74732 459518 74788
rect 419916 74424 419972 74732
rect 559944 73948 566300 74004
rect 566356 73948 566366 74004
rect 590482 73388 590492 73444
rect 590548 73416 595672 73444
rect 590548 73388 597000 73416
rect 595560 73192 597000 73388
rect 269864 73052 273084 73108
rect 273140 73052 273150 73108
rect 559944 72380 564620 72436
rect 564676 72380 564686 72436
rect 459340 72212 460040 72268
rect 447682 72156 447692 72212
rect 447748 72156 459396 72212
rect 559570 70812 559580 70868
rect 559636 70812 559646 70868
rect 269864 70140 273308 70196
rect 273364 70140 273374 70196
rect 446002 69356 446012 69412
rect 446068 69356 459396 69412
rect 459340 69300 460040 69356
rect 559944 69244 563276 69300
rect 563332 69244 563342 69300
rect 419916 68012 421932 68068
rect 421988 68012 452732 68068
rect 452788 68012 452798 68068
rect 419916 67480 419972 68012
rect 559458 67676 559468 67732
rect 559524 67676 559534 67732
rect 269864 67228 273196 67284
rect 273252 67228 273262 67284
rect 444322 66444 444332 66500
rect 444388 66444 459396 66500
rect 459340 66388 460040 66444
rect 559944 66108 563164 66164
rect 563220 66108 563230 66164
rect -960 65044 480 65240
rect -960 65016 27692 65044
rect 392 64988 27692 65016
rect 27748 64988 27758 65044
rect 559944 64540 563052 64596
rect 563108 64540 563118 64596
rect 269864 64316 290108 64372
rect 290164 64316 290174 64372
rect 449362 63532 449372 63588
rect 449428 63532 459396 63588
rect 459340 63476 460040 63532
rect 559944 62972 562940 63028
rect 562996 62972 563006 63028
rect 357746 61628 357756 61684
rect 357812 61628 360136 61684
rect 269864 61404 278012 61460
rect 278068 61404 278078 61460
rect 559944 61404 574588 61460
rect 574644 61404 574654 61460
rect 419972 61292 422044 61348
rect 422100 61292 456092 61348
rect 456148 61292 456158 61348
rect 419972 61236 420028 61292
rect 419916 61180 420028 61236
rect 419916 60536 419972 61180
rect 441074 60620 441084 60676
rect 441140 60620 459396 60676
rect 459340 60564 460040 60620
rect 595560 60004 597000 60200
rect 577042 59948 577052 60004
rect 577108 59976 597000 60004
rect 577108 59948 595672 59976
rect 559944 59836 562828 59892
rect 562884 59836 562894 59892
rect 427634 59612 427644 59668
rect 427700 59612 457660 59668
rect 457716 59612 457726 59668
rect 564396 58828 567868 58884
rect 567924 58828 567934 58884
rect 269864 58492 276332 58548
rect 276388 58492 276398 58548
rect 564396 58324 564452 58828
rect 559944 58268 564452 58324
rect 457650 57708 457660 57764
rect 457716 57708 459396 57764
rect 459340 57652 460040 57708
rect 559944 56700 564396 56756
rect 564452 56700 564462 56756
rect 269864 55580 287980 55636
rect 288036 55580 288046 55636
rect 457762 54796 457772 54852
rect 457828 54796 459396 54852
rect 459340 54740 460040 54796
rect 419356 52948 419412 53592
rect 419234 52892 419244 52948
rect 419300 52892 454412 52948
rect 454468 52892 454478 52948
rect 273074 52780 273084 52836
rect 273140 52780 420028 52836
rect 420084 52780 420094 52836
rect 269836 52612 269892 52696
rect 273298 52668 273308 52724
rect 273364 52668 420140 52724
rect 420196 52668 420206 52724
rect 269836 52556 290668 52612
rect 290612 52052 290668 52556
rect 290612 51996 419244 52052
rect 419300 51996 419310 52052
rect 356178 51884 356188 51940
rect 356244 51884 357756 51940
rect 357812 51884 459396 51940
rect 459340 51828 460040 51884
rect 290098 51772 290108 51828
rect 290164 51772 421708 51828
rect 421764 51772 421774 51828
rect 392 51128 4284 51156
rect -960 51100 4284 51128
rect 4340 51100 4350 51156
rect -960 50904 480 51100
rect 273186 50652 273196 50708
rect 273252 50652 420252 50708
rect 420308 50652 420318 50708
rect 276322 50540 276332 50596
rect 276388 50540 421932 50596
rect 421988 50540 421998 50596
rect 287970 50428 287980 50484
rect 288036 50428 422044 50484
rect 422100 50428 422110 50484
rect 4162 50316 4172 50372
rect 4228 50316 269500 50372
rect 269556 50316 269566 50372
rect 278002 50316 278012 50372
rect 278068 50316 421820 50372
rect 421876 50316 421886 50372
rect 425842 50316 425852 50372
rect 425908 50316 562828 50372
rect 562884 50316 562894 50372
rect 307430 50204 307468 50260
rect 307524 50204 307534 50260
rect 314178 50204 314188 50260
rect 314244 50204 314282 50260
rect 320898 50204 320908 50260
rect 320964 50204 321356 50260
rect 321412 50204 321422 50260
rect 293570 50092 293580 50148
rect 293636 50092 356188 50148
rect 356244 50092 356254 50148
rect 180786 49868 180796 49924
rect 180852 49868 288316 49924
rect 288372 49868 288382 49924
rect 167458 49756 167468 49812
rect 167524 49756 275660 49812
rect 275716 49756 275726 49812
rect 4386 49644 4396 49700
rect 4452 49644 271180 49700
rect 271236 49644 271246 49700
rect 91298 49532 91308 49588
rect 91364 49532 362124 49588
rect 362180 49532 362190 49588
rect 47842 48636 47852 48692
rect 47908 48636 48524 48692
rect 48580 48636 97356 48692
rect 97412 48636 293580 48692
rect 293636 48636 293646 48692
rect 212258 48524 212268 48580
rect 212324 48524 267260 48580
rect 267316 48524 267326 48580
rect 289874 48524 289884 48580
rect 289940 48524 300748 48580
rect 300804 48524 300814 48580
rect 197922 48300 197932 48356
rect 197988 48300 281372 48356
rect 281428 48300 281438 48356
rect 178882 48188 178892 48244
rect 178948 48188 277564 48244
rect 277620 48188 277630 48244
rect 127474 48076 127484 48132
rect 127540 48076 275660 48132
rect 275716 48076 275726 48132
rect 93202 47964 93212 48020
rect 93268 47964 271068 48020
rect 271124 47964 271134 48020
rect 87490 47852 87500 47908
rect 87556 47852 267148 47908
rect 267204 47852 267214 47908
rect 595560 46760 597000 46984
rect 184594 46172 184604 46228
rect 184660 46172 277452 46228
rect 277508 46172 277518 46228
rect 207442 45164 207452 45220
rect 207508 45164 279132 45220
rect 279188 45164 279198 45220
rect 138898 45052 138908 45108
rect 138964 45052 277340 45108
rect 277396 45052 277406 45108
rect 110338 44940 110348 44996
rect 110404 44940 270956 44996
rect 271012 44940 271022 44996
rect 104626 44828 104636 44884
rect 104692 44828 270620 44884
rect 270676 44828 270686 44884
rect 98914 44716 98924 44772
rect 98980 44716 270844 44772
rect 270900 44716 270910 44772
rect 148418 44604 148428 44660
rect 148484 44604 359212 44660
rect 359268 44604 359278 44660
rect 142818 44492 142828 44548
rect 142884 44492 358764 44548
rect 358820 44492 358830 44548
rect 156034 42924 156044 42980
rect 156100 42924 275548 42980
rect 275604 42924 275614 42980
rect 188402 42812 188412 42868
rect 188468 42812 411740 42868
rect 411796 42812 411806 42868
rect 203634 41692 203644 41748
rect 203700 41692 283388 41748
rect 283444 41692 283454 41748
rect 175074 41580 175084 41636
rect 175140 41580 284956 41636
rect 285012 41580 285022 41636
rect 116050 41468 116060 41524
rect 116116 41468 270732 41524
rect 270788 41468 270798 41524
rect 159842 41356 159852 41412
rect 159908 41356 358988 41412
rect 359044 41356 359054 41412
rect 97010 41244 97020 41300
rect 97076 41244 362012 41300
rect 362068 41244 362078 41300
rect 68450 41132 68460 41188
rect 68516 41132 358652 41188
rect 358708 41132 358718 41188
rect 161746 39452 161756 39508
rect 161812 39452 279020 39508
rect 279076 39452 279086 39508
rect 192210 38332 192220 38388
rect 192276 38332 290332 38388
rect 290388 38332 290398 38388
rect 182690 38220 182700 38276
rect 182756 38220 355292 38276
rect 355348 38220 355358 38276
rect 171378 38108 171388 38164
rect 171444 38108 358764 38164
rect 358820 38108 358830 38164
rect 119858 37996 119868 38052
rect 119924 37996 358988 38052
rect 359044 37996 359054 38052
rect 108434 37884 108444 37940
rect 108500 37884 359212 37940
rect 359268 37884 359278 37940
rect 57138 37772 57148 37828
rect 57204 37772 360556 37828
rect 360612 37772 360622 37828
rect -960 36932 480 37016
rect -960 36876 4396 36932
rect 4452 36876 4462 36932
rect -960 36792 480 36876
rect 209346 36204 209356 36260
rect 209412 36204 284732 36260
rect 284788 36204 284798 36260
rect 76066 36092 76076 36148
rect 76132 36092 270508 36148
rect 270564 36092 270574 36148
rect 211250 34972 211260 35028
rect 211316 34972 355740 35028
rect 355796 34972 355806 35028
rect 121762 34860 121772 34916
rect 121828 34860 275548 34916
rect 275604 34860 275614 34916
rect 194114 34748 194124 34804
rect 194180 34748 358652 34804
rect 358708 34748 358718 34804
rect 81778 34636 81788 34692
rect 81844 34636 269612 34692
rect 269668 34636 269678 34692
rect 74162 34524 74172 34580
rect 74228 34524 355516 34580
rect 355572 34524 355582 34580
rect 62738 34412 62748 34468
rect 62804 34412 360332 34468
rect 360388 34412 360398 34468
rect 595560 33684 597000 33768
rect 326722 33628 326732 33684
rect 326788 33628 597000 33684
rect 595560 33544 597000 33628
rect 133186 32956 133196 33012
rect 133252 32956 269500 33012
rect 269556 32956 269566 33012
rect 89394 32844 89404 32900
rect 89460 32844 282156 32900
rect 282212 32844 282222 32900
rect 102722 32732 102732 32788
rect 102788 32732 411852 32788
rect 411908 32732 411918 32788
rect 144610 31276 144620 31332
rect 144676 31276 278908 31332
rect 278964 31276 278974 31332
rect 152226 31164 152236 31220
rect 152292 31164 289996 31220
rect 290052 31164 290062 31220
rect 79874 31052 79884 31108
rect 79940 31052 355404 31108
rect 355460 31052 355470 31108
rect 169362 29484 169372 29540
rect 169428 29484 289772 29540
rect 289828 29484 289838 29540
rect 83682 29372 83692 29428
rect 83748 29372 281260 29428
rect 281316 29372 281326 29428
rect 173170 26124 173180 26180
rect 173236 26124 269724 26180
rect 269780 26124 269790 26180
rect 146514 26012 146524 26068
rect 146580 26012 283164 26068
rect 283220 26012 283230 26068
rect 196018 24556 196028 24612
rect 196084 24556 270508 24612
rect 270564 24556 270574 24612
rect 135090 24444 135100 24500
rect 135156 24444 288092 24500
rect 288148 24444 288158 24500
rect 72258 24332 72268 24388
rect 72324 24332 279468 24388
rect 279524 24332 279534 24388
rect 392 22904 10892 22932
rect -960 22876 10892 22904
rect 10948 22876 10958 22932
rect -960 22680 480 22876
rect 186498 20972 186508 21028
rect 186564 20972 290892 21028
rect 290948 20972 290958 21028
rect 595560 20356 597000 20552
rect 424162 20300 424172 20356
rect 424228 20328 597000 20356
rect 424228 20300 595672 20328
rect 95106 19404 95116 19460
rect 95172 19404 283052 19460
rect 283108 19404 283118 19460
rect 60834 19292 60844 19348
rect 60900 19292 277676 19348
rect 277732 19292 277742 19348
rect 123666 17724 123676 17780
rect 123732 17724 287532 17780
rect 287588 17724 287598 17780
rect 55122 17612 55132 17668
rect 55188 17612 276780 17668
rect 276836 17612 276846 17668
rect 129378 16044 129388 16100
rect 129444 16044 288428 16100
rect 288484 16044 288494 16100
rect 47506 15932 47516 15988
rect 47572 15932 275884 15988
rect 275940 15932 275950 15988
rect 201730 14476 201740 14532
rect 201796 14476 271404 14532
rect 271460 14476 271470 14532
rect 140802 14364 140812 14420
rect 140868 14364 290220 14420
rect 290276 14364 290286 14420
rect 77970 14252 77980 14308
rect 78036 14252 280364 14308
rect 280420 14252 280430 14308
rect 163650 12572 163660 12628
rect 163716 12572 291116 12628
rect 291172 12572 291182 12628
rect 150546 10892 150556 10948
rect 150612 10892 277228 10948
rect 277284 10892 277294 10948
rect 68898 9324 68908 9380
rect 68964 9324 278572 9380
rect 278628 9324 278638 9380
rect 131506 9212 131516 9268
rect 131572 9212 411628 9268
rect 411684 9212 411694 9268
rect 392 8792 4172 8820
rect -960 8764 4172 8792
rect 4228 8764 4238 8820
rect -960 8568 480 8764
rect 118178 7756 118188 7812
rect 118244 7756 286636 7812
rect 286692 7756 286702 7812
rect 112466 7644 112476 7700
rect 112532 7644 285740 7700
rect 285796 7644 285806 7700
rect 106754 7532 106764 7588
rect 106820 7532 284844 7588
rect 284900 7532 284910 7588
rect 595560 7140 597000 7336
rect 565282 7084 565292 7140
rect 565348 7112 597000 7140
rect 565348 7084 595672 7112
rect 190530 6076 190540 6132
rect 190596 6076 269612 6132
rect 269668 6076 269678 6132
rect 158162 5964 158172 6020
rect 158228 5964 291452 6020
rect 291508 5964 291518 6020
rect 11554 5852 11564 5908
rect 11620 5852 47852 5908
rect 47908 5852 47918 5908
rect 101042 5852 101052 5908
rect 101108 5852 283948 5908
rect 284004 5852 284014 5908
rect 205762 4956 205772 5012
rect 205828 4956 350476 5012
rect 350532 4956 350542 5012
rect 38434 4844 38444 4900
rect 38500 4844 45612 4900
rect 45668 4844 45678 4900
rect 125794 4844 125804 4900
rect 125860 4844 272972 4900
rect 273028 4844 273038 4900
rect 200050 4732 200060 4788
rect 200116 4732 348572 4788
rect 348628 4732 348638 4788
rect 66770 4620 66780 4676
rect 66836 4620 68908 4676
rect 68964 4620 68974 4676
rect 177202 4620 177212 4676
rect 177268 4620 331772 4676
rect 331828 4620 331838 4676
rect 51986 4508 51996 4564
rect 52052 4508 58940 4564
rect 58996 4508 59006 4564
rect 165778 4508 165788 4564
rect 165844 4508 330092 4564
rect 330148 4508 330158 4564
rect 41122 4396 41132 4452
rect 41188 4396 49420 4452
rect 49476 4396 49486 4452
rect 51874 4396 51884 4452
rect 51940 4396 64652 4452
rect 64708 4396 64718 4452
rect 154354 4396 154364 4452
rect 154420 4396 336812 4452
rect 336868 4396 336878 4452
rect 40114 4284 40124 4340
rect 40180 4284 53228 4340
rect 53284 4284 53294 4340
rect 85810 4284 85820 4340
rect 85876 4284 274652 4340
rect 274708 4284 274718 4340
rect 38546 4172 38556 4228
rect 38612 4172 39900 4228
rect 39956 4172 39966 4228
rect 40226 4172 40236 4228
rect 40292 4172 70364 4228
rect 70420 4172 70430 4228
rect 114370 4172 114380 4228
rect 114436 4172 328412 4228
rect 328468 4172 328478 4228
rect 429202 4172 429212 4228
rect 429268 4172 572908 4228
rect 579618 4172 579628 4228
rect 579684 4172 580636 4228
rect 580692 4172 580702 4228
rect 582978 4172 582988 4228
rect 583044 4172 584444 4228
rect 584500 4172 584510 4228
rect 572852 4116 572908 4172
rect 137218 4060 137228 4116
rect 137284 4060 274876 4116
rect 274932 4060 274942 4116
rect 572852 4060 582540 4116
rect 582596 4060 582606 4116
<< via3 >>
rect 190428 591276 190484 591332
rect 408268 591276 408324 591332
rect 474348 591276 474404 591332
rect 192780 591052 192836 591108
rect 193004 590828 193060 590884
rect 190540 590604 190596 590660
rect 546028 590604 546084 590660
rect 192668 590492 192724 590548
rect 545580 590492 545636 590548
rect 192892 590380 192948 590436
rect 590492 588588 590548 588644
rect 184716 565068 184772 565124
rect 4172 558908 4228 558964
rect 187852 557900 187908 557956
rect 186396 550732 186452 550788
rect 590604 548940 590660 548996
rect 7532 544796 7588 544852
rect 187516 543564 187572 543620
rect 186284 536396 186340 536452
rect 187740 529228 187796 529284
rect 187628 522060 187684 522116
rect 4284 516572 4340 516628
rect 186172 514892 186228 514948
rect 590716 509292 590772 509348
rect 187404 507724 187460 507780
rect 166236 506492 166292 506548
rect 187404 506492 187460 506548
rect 57932 502460 57988 502516
rect 167916 500556 167972 500612
rect 188972 493388 189028 493444
rect 189532 486220 189588 486276
rect 189420 479052 189476 479108
rect 4172 476252 4228 476308
rect 146972 476252 147028 476308
rect 141932 474236 141988 474292
rect 187964 471884 188020 471940
rect 590828 469644 590884 469700
rect 4284 469532 4340 469588
rect 145292 469532 145348 469588
rect 162540 464716 162596 464772
rect 187964 457548 188020 457604
rect 166124 450380 166180 450436
rect 167804 443212 167860 443268
rect 187292 436044 187348 436100
rect 140252 431900 140308 431956
rect 590940 430108 590996 430164
rect 187404 428876 187460 428932
rect 189308 421708 189364 421764
rect 188076 414540 188132 414596
rect 192668 409388 192724 409444
rect 192780 409276 192836 409332
rect 308028 409276 308084 409332
rect 546028 409164 546084 409220
rect 187628 408940 187684 408996
rect 376348 408940 376404 408996
rect 302652 408828 302708 408884
rect 261212 407932 261268 407988
rect 238140 407708 238196 407764
rect 477148 407708 477204 407764
rect 245196 407596 245252 407652
rect 250348 407596 250404 407652
rect 375452 407596 375508 407652
rect 475468 407596 475524 407652
rect 545580 407484 545636 407540
rect 286300 406924 286356 406980
rect 303996 406924 304052 406980
rect 250348 406812 250404 406868
rect 190540 406476 190596 406532
rect 230972 406476 231028 406532
rect 186284 405916 186340 405972
rect 378476 405916 378532 405972
rect 261212 404796 261268 404852
rect 187516 404236 187572 404292
rect 376460 404236 376516 404292
rect 190428 404012 190484 404068
rect 187852 402780 187908 402836
rect 375676 402780 375732 402836
rect 231532 402444 231588 402500
rect 590604 402444 590660 402500
rect 231644 402332 231700 402388
rect 590940 402332 590996 402388
rect 236012 400876 236068 400932
rect 186396 399308 186452 399364
rect 378700 399308 378756 399364
rect 234892 398972 234948 399028
rect 590492 398972 590548 399028
rect 184716 397852 184772 397908
rect 378812 397852 378868 397908
rect 230076 397292 230132 397348
rect 590716 397292 590772 397348
rect 189308 396396 189364 396452
rect 378924 396396 378980 396452
rect 187740 396284 187796 396340
rect 376572 396284 376628 396340
rect 186172 396172 186228 396228
rect 378588 396172 378644 396228
rect 372988 393148 373044 393204
rect 236236 392476 236292 392532
rect 237916 392364 237972 392420
rect 103292 391692 103348 391748
rect 590156 390348 590212 390404
rect 4172 389564 4228 389620
rect 238252 388108 238308 388164
rect 282156 388108 282212 388164
rect 297388 388108 297444 388164
rect 234780 387212 234836 387268
rect 590156 387212 590212 387268
rect 99932 386876 99988 386932
rect 372316 386092 372372 386148
rect 372428 385980 372484 386036
rect 237804 385868 237860 385924
rect 375564 385868 375620 385924
rect 267820 385420 267876 385476
rect 273196 385420 273252 385476
rect 236124 385308 236180 385364
rect 266028 385308 266084 385364
rect 269612 385308 269668 385364
rect 271404 385308 271460 385364
rect 275884 385308 275940 385364
rect 281260 385308 281316 385364
rect 283052 385308 283108 385364
rect 287532 385308 287588 385364
rect 288428 385308 288484 385364
rect 289324 385308 289380 385364
rect 290220 385308 290276 385364
rect 291116 385308 291172 385364
rect 292908 385308 292964 385364
rect 293804 385308 293860 385364
rect 294700 385308 294756 385364
rect 309036 385308 309092 385364
rect 250348 384524 250404 384580
rect 281260 384524 281316 384580
rect 275884 384412 275940 384468
rect 283052 384412 283108 384468
rect 309036 384300 309092 384356
rect 266028 384188 266084 384244
rect 291116 384188 291172 384244
rect 292908 384076 292964 384132
rect 293804 383964 293860 384020
rect 294700 383852 294756 383908
rect 378924 382396 378980 382452
rect 4172 380492 4228 380548
rect 209132 380492 209188 380548
rect 199724 377468 199780 377524
rect 199500 376348 199556 376404
rect 199276 375228 199332 375284
rect 199388 374108 199444 374164
rect 199164 372988 199220 373044
rect 199052 371868 199108 371924
rect 560252 371196 560308 371252
rect 378924 370076 378980 370132
rect 573132 368956 573188 369012
rect 378924 368732 378980 368788
rect 571564 368732 571620 368788
rect 574700 367836 574756 367892
rect 568204 366716 568260 366772
rect 573020 365596 573076 365652
rect 379596 364476 379652 364532
rect 571452 363356 571508 363412
rect 199724 363020 199780 363076
rect 572908 362236 572964 362292
rect 379596 362012 379652 362068
rect 564956 362012 565012 362068
rect 379596 361116 379652 361172
rect 566524 359996 566580 360052
rect 199500 359660 199556 359716
rect 571340 358876 571396 358932
rect 379596 358652 379652 358708
rect 569772 358652 569828 358708
rect 571228 357756 571284 357812
rect 569548 356636 569604 356692
rect 199276 356300 199332 356356
rect 569660 355516 569716 355572
rect 566412 354396 566468 354452
rect 564844 353276 564900 353332
rect 199388 352940 199444 352996
rect 379596 352156 379652 352212
rect 567980 351036 568036 351092
rect 590492 350700 590548 350756
rect 379596 350252 379652 350308
rect 568092 350252 568148 350308
rect 566188 349916 566244 349972
rect 199164 349580 199220 349636
rect 564732 348796 564788 348852
rect 566300 347676 566356 347732
rect 4172 347228 4228 347284
rect 564620 346556 564676 346612
rect 559580 345436 559636 345492
rect 4172 345212 4228 345268
rect 138572 345212 138628 345268
rect 389116 344316 389172 344372
rect 559468 343196 559524 343252
rect 540092 342076 540148 342132
rect 555212 340956 555268 341012
rect 556892 339836 556948 339892
rect 235900 339164 235956 339220
rect 574588 338716 574644 338772
rect 425852 337596 425908 337652
rect 567868 336476 567924 336532
rect 564508 335356 564564 335412
rect 393932 334236 393988 334292
rect 223356 333788 223412 333844
rect 390572 333116 390628 333172
rect 219996 332668 220052 332724
rect 388892 331996 388948 332052
rect 389116 331772 389172 331828
rect 563276 331772 563332 331828
rect 380492 330876 380548 330932
rect 235004 330428 235060 330484
rect 387212 329756 387268 329812
rect 234444 329308 234500 329364
rect 385532 328636 385588 328692
rect 226716 328188 226772 328244
rect 451052 327516 451108 327572
rect 229964 327068 230020 327124
rect 382172 326396 382228 326452
rect 199052 326060 199108 326116
rect 228396 325948 228452 326004
rect 392252 325276 392308 325332
rect 231420 324828 231476 324884
rect 520044 324268 520100 324324
rect 383852 324156 383908 324212
rect 226604 323708 226660 323764
rect 456092 323036 456148 323092
rect 195244 322700 195300 322756
rect 231308 322588 231364 322644
rect 195244 321916 195300 321972
rect 442652 321916 442708 321972
rect 229852 321468 229908 321524
rect 231196 320348 231252 320404
rect 378812 320012 378868 320068
rect 437612 320012 437668 320068
rect 375676 319676 375732 319732
rect 434252 319676 434308 319732
rect 232428 319228 232484 319284
rect 378700 318332 378756 318388
rect 432572 318332 432628 318388
rect 233212 318108 233268 318164
rect 376460 317436 376516 317492
rect 378812 317436 378868 317492
rect 233324 316988 233380 317044
rect 378476 316652 378532 316708
rect 427532 316652 427588 316708
rect 233100 315868 233156 315924
rect 376572 315196 376628 315252
rect 378812 315084 378868 315140
rect 430892 315084 430948 315140
rect 429212 314972 429268 315028
rect 232652 314748 232708 314804
rect 376348 314076 376404 314132
rect 232540 313628 232596 313684
rect 378588 313404 378644 313460
rect 425964 313404 426020 313460
rect 454412 313292 454468 313348
rect 378588 312956 378644 313012
rect 232876 312508 232932 312564
rect 232764 311388 232820 311444
rect 590604 311052 590660 311108
rect 232988 310268 233044 310324
rect 383068 309596 383124 309652
rect 384748 308476 384804 308532
rect 379484 306236 379540 306292
rect 4172 305788 4228 305844
rect 379372 305116 379428 305172
rect 228284 304892 228340 304948
rect 4284 304668 4340 304724
rect 379260 303996 379316 304052
rect 29372 303548 29428 303604
rect 379036 302876 379092 302932
rect 32732 302540 32788 302596
rect 378924 301756 378980 301812
rect 27804 301308 27860 301364
rect 379148 300636 379204 300692
rect 12572 300188 12628 300244
rect 378812 299516 378868 299572
rect 10892 299292 10948 299348
rect 47404 299292 47460 299348
rect 376348 298396 376404 298452
rect 228284 297948 228340 298004
rect 47404 297388 47460 297444
rect 48524 297388 48580 297444
rect 138572 296828 138628 296884
rect 186508 296044 186564 296100
rect 187292 296044 187348 296100
rect 209132 295708 209188 295764
rect 140252 294588 140308 294644
rect 141932 293468 141988 293524
rect 145292 292348 145348 292404
rect 146972 291228 147028 291284
rect 188076 290556 188132 290612
rect 187404 290220 187460 290276
rect 411740 289436 411796 289492
rect 186620 288988 186676 289044
rect 187404 288988 187460 289044
rect 188076 288988 188132 289044
rect 375228 288316 375284 288372
rect 192892 286748 192948 286804
rect 167804 286636 167860 286692
rect 188300 286636 188356 286692
rect 162540 286524 162596 286580
rect 188524 286524 188580 286580
rect 375228 286076 375284 286132
rect 167916 285516 167972 285572
rect 188188 285516 188244 285572
rect 166124 285404 166180 285460
rect 188412 285404 188468 285460
rect 193004 284508 193060 284564
rect 166236 284172 166292 284228
rect 424172 283948 424228 284004
rect 375676 283836 375732 283892
rect 190652 283388 190708 283444
rect 193116 282268 193172 282324
rect 376460 281596 376516 281652
rect 188188 281372 188244 281428
rect 420812 280588 420868 280644
rect 234892 280028 234948 280084
rect 188972 279916 189028 279972
rect 231532 278908 231588 278964
rect 411628 278236 411684 278292
rect 189532 278012 189588 278068
rect 231084 278012 231140 278068
rect 230076 277788 230132 277844
rect 231756 276668 231812 276724
rect 189420 276332 189476 276388
rect 231644 275548 231700 275604
rect 452732 275548 452788 275604
rect 234780 274428 234836 274484
rect 188636 273868 188692 273924
rect 189084 273868 189140 273924
rect 379484 273868 379540 273924
rect 380268 273868 380324 273924
rect 440972 273868 441028 273924
rect 235788 273308 235844 273364
rect 411852 272636 411908 272692
rect 231756 272188 231812 272244
rect 375788 271516 375844 271572
rect 590828 271404 590884 271460
rect 188524 271292 188580 271348
rect 231532 271292 231588 271348
rect 235116 271068 235172 271124
rect 379820 270508 379876 270564
rect 447692 270508 447748 270564
rect 375900 270396 375956 270452
rect 379260 270396 379316 270452
rect 380044 270396 380100 270452
rect 235340 269948 235396 270004
rect 187964 269836 188020 269892
rect 189532 269836 189588 269892
rect 234668 268828 234724 268884
rect 380044 268828 380100 268884
rect 446012 268828 446068 268884
rect 379036 268716 379092 268772
rect 379932 268716 379988 268772
rect 188412 267932 188468 267988
rect 235676 267932 235732 267988
rect 234892 267708 234948 267764
rect 379932 267148 379988 267204
rect 444332 267148 444388 267204
rect 378588 267036 378644 267092
rect 234556 266588 234612 266644
rect 188300 266252 188356 266308
rect 235900 266252 235956 266308
rect 375228 265916 375284 265972
rect 234780 265468 234836 265524
rect 378924 265468 378980 265524
rect 379708 265468 379764 265524
rect 449372 265468 449428 265524
rect 378700 264796 378756 264852
rect 186508 264572 186564 264628
rect 235564 264572 235620 264628
rect 379148 263788 379204 263844
rect 380156 263788 380212 263844
rect 419356 263788 419412 263844
rect 378924 263676 378980 263732
rect 10892 262780 10948 262836
rect 378476 262556 378532 262612
rect 186620 261772 186676 261828
rect 189196 261772 189252 261828
rect 376124 261436 376180 261492
rect 378812 260428 378868 260484
rect 422492 260428 422548 260484
rect 376236 259196 376292 259252
rect 237580 257404 237636 257460
rect 380044 257404 380100 257460
rect 269276 257292 269332 257348
rect 348572 257292 348628 257348
rect 235788 256508 235844 256564
rect 590492 256508 590548 256564
rect 235900 256284 235956 256340
rect 379708 256284 379764 256340
rect 232540 256172 232596 256228
rect 273868 256172 273924 256228
rect 362012 255948 362068 256004
rect 375788 255948 375844 256004
rect 362124 255836 362180 255892
rect 375900 255836 375956 255892
rect 235452 255724 235508 255780
rect 379932 255724 379988 255780
rect 231756 255276 231812 255332
rect 590604 255276 590660 255332
rect 235116 255164 235172 255220
rect 590828 255164 590884 255220
rect 189196 255052 189252 255108
rect 378812 255052 378868 255108
rect 235788 254716 235844 254772
rect 380156 254716 380212 254772
rect 232652 254604 232708 254660
rect 273980 254604 274036 254660
rect 251916 253596 251972 253652
rect 252588 253596 252644 253652
rect 258860 253596 258916 253652
rect 259756 253596 259812 253652
rect 260652 253596 260708 253652
rect 373772 253260 373828 253316
rect 291452 252028 291508 252084
rect 189084 251916 189140 251972
rect 380268 251916 380324 251972
rect 236012 251692 236068 251748
rect 231532 250236 231588 250292
rect 379820 250236 379876 250292
rect 267148 249340 267204 249396
rect 378700 248556 378756 248612
rect 4060 248444 4116 248500
rect 378588 248332 378644 248388
rect 378924 247660 378980 247716
rect 231868 246876 231924 246932
rect 188972 246764 189028 246820
rect 383068 246764 383124 246820
rect 395612 246764 395668 246820
rect 231084 246652 231140 246708
rect 384748 246652 384804 246708
rect 267372 246316 267428 246372
rect 404012 246316 404068 246372
rect 268716 245308 268772 245364
rect 46172 242508 46228 242564
rect 234668 241052 234724 241108
rect 590828 241052 590884 241108
rect 212492 240492 212548 240548
rect 235564 239484 235620 239540
rect 590156 239484 590212 239540
rect 234556 239372 234612 239428
rect 590604 239372 590660 239428
rect 74956 238476 75012 238532
rect 76972 238476 77028 238532
rect 95452 238140 95508 238196
rect 95452 237692 95508 237748
rect 223356 236684 223412 236740
rect 519148 236684 519204 236740
rect 236124 236572 236180 236628
rect 234780 236460 234836 236516
rect 590492 236460 590548 236516
rect 234892 236348 234948 236404
rect 590716 236348 590772 236404
rect 422492 235116 422548 235172
rect 423276 235116 423332 235172
rect 423276 234556 423332 234612
rect 232764 234332 232820 234388
rect 270620 234332 270676 234388
rect 376124 232652 376180 232708
rect 590156 231980 590212 232036
rect 51996 231084 52052 231140
rect 378476 230972 378532 231028
rect 376348 229292 376404 229348
rect 12572 220220 12628 220276
rect 232876 217756 232932 217812
rect 269724 217756 269780 217812
rect 233100 216524 233156 216580
rect 270732 216524 270788 216580
rect 233212 216300 233268 216356
rect 274204 216300 274260 216356
rect 51884 215964 51940 216020
rect 233324 214284 233380 214340
rect 269388 214284 269444 214340
rect 219996 214172 220052 214228
rect 457772 214172 457828 214228
rect 232988 213164 233044 213220
rect 274092 213164 274148 213220
rect 232428 212940 232484 212996
rect 275772 212940 275828 212996
rect 307468 212828 307524 212884
rect 314188 212716 314244 212772
rect 320908 212604 320964 212660
rect 376236 212492 376292 212548
rect 237804 211484 237860 211540
rect 235004 211372 235060 211428
rect 231196 211260 231252 211316
rect 272412 211260 272468 211316
rect 229852 211148 229908 211204
rect 226716 211036 226772 211092
rect 269836 211036 269892 211092
rect 237692 210924 237748 210980
rect 272748 210700 272804 210756
rect 50316 210140 50372 210196
rect 49532 210028 49588 210084
rect 234444 209916 234500 209972
rect 231308 209804 231364 209860
rect 231420 209692 231476 209748
rect 229964 209580 230020 209636
rect 228396 209468 228452 209524
rect 226604 209356 226660 209412
rect 272412 209804 272468 209860
rect 272860 209468 272916 209524
rect 272636 209356 272692 209412
rect 273196 209244 273252 209300
rect 273084 209132 273140 209188
rect 272524 209020 272580 209076
rect 4172 206332 4228 206388
rect 519148 204988 519204 205044
rect 516236 201628 516292 201684
rect 269836 201516 269892 201572
rect 383964 200060 384020 200116
rect 516236 199388 516292 199444
rect 273196 198268 273252 198324
rect 497644 198156 497700 198212
rect 499100 198156 499156 198212
rect 502236 198156 502292 198212
rect 481292 198044 481348 198100
rect 273084 195356 273140 195412
rect 272524 192444 272580 192500
rect 590828 192332 590884 192388
rect 272412 189532 272468 189588
rect 272860 186620 272916 186676
rect 272748 183708 272804 183764
rect 27804 177884 27860 177940
rect 275772 177884 275828 177940
rect 274204 174972 274260 175028
rect 269388 172060 269444 172116
rect 270732 169148 270788 169204
rect 273980 166236 274036 166292
rect 4172 163996 4228 164052
rect 273868 163324 273924 163380
rect 375564 160748 375620 160804
rect 373100 160636 373156 160692
rect 269724 160412 269780 160468
rect 270620 157500 270676 157556
rect 296492 156604 296548 156660
rect 274652 156268 274708 156324
rect 274092 154588 274148 154644
rect 367052 154364 367108 154420
rect 291564 154252 291620 154308
rect 371308 154140 371364 154196
rect 372316 154140 372372 154196
rect 273756 154028 273812 154084
rect 372988 154028 373044 154084
rect 367052 153916 367108 153972
rect 375452 153916 375508 153972
rect 371308 153692 371364 153748
rect 495852 152908 495908 152964
rect 501340 152908 501396 152964
rect 590716 152684 590772 152740
rect 393932 152012 393988 152068
rect 456988 152012 457044 152068
rect 7532 149884 7588 149940
rect 465500 149436 465556 149492
rect 465500 149100 465556 149156
rect 509740 149436 509796 149492
rect 509740 149100 509796 149156
rect 269276 148764 269332 148820
rect 540092 148652 540148 148708
rect 563164 148652 563220 148708
rect 456988 148540 457044 148596
rect 555212 148092 555268 148148
rect 563052 148092 563108 148148
rect 556892 147980 556948 148036
rect 562940 147980 562996 148036
rect 390572 145068 390628 145124
rect 388892 142156 388948 142212
rect 380492 139244 380548 139300
rect 387212 136332 387268 136388
rect 273756 136108 273812 136164
rect 32732 135548 32788 135604
rect 385532 133420 385588 133476
rect 451052 130508 451108 130564
rect 395612 128492 395668 128548
rect 457884 128492 457940 128548
rect 382172 127596 382228 127652
rect 392252 124684 392308 124740
rect 383852 121772 383908 121828
rect 560252 120876 560308 120932
rect 562828 120876 562884 120932
rect 404012 120092 404068 120148
rect 457996 120092 458052 120148
rect 456092 118860 456148 118916
rect 313404 116732 313460 116788
rect 419356 116060 419412 116116
rect 441084 116060 441140 116116
rect 442652 115836 442708 115892
rect 437612 113036 437668 113092
rect 590604 113036 590660 113092
rect 434252 110124 434308 110180
rect 423276 109116 423332 109172
rect 427644 109116 427700 109172
rect 296492 107996 296548 108052
rect 432572 107212 432628 107268
rect 562828 106876 562884 106932
rect 571564 105308 571620 105364
rect 291564 105084 291620 105140
rect 430892 104300 430948 104356
rect 573132 103740 573188 103796
rect 574700 102172 574756 102228
rect 427532 101388 427588 101444
rect 568204 100604 568260 100660
rect 573020 99036 573076 99092
rect 429212 98476 429268 98532
rect 564956 97468 565012 97524
rect 571452 95900 571508 95956
rect 454412 95564 454468 95620
rect 572908 94332 572964 94388
rect 29372 93212 29428 93268
rect 569772 92764 569828 92820
rect 425964 92652 426020 92708
rect 566524 91196 566580 91252
rect 424172 89740 424228 89796
rect 571340 89628 571396 89684
rect 571228 88060 571284 88116
rect 420812 86828 420868 86884
rect 569548 86492 569604 86548
rect 569660 84924 569716 84980
rect 457884 83916 457940 83972
rect 566412 83356 566468 83412
rect 564844 81788 564900 81844
rect 457996 81004 458052 81060
rect 568092 80220 568148 80276
rect 567980 78652 568036 78708
rect 452732 78092 452788 78148
rect 566188 77084 566244 77140
rect 564732 75516 564788 75572
rect 440972 75180 441028 75236
rect 566300 73948 566356 74004
rect 590492 73388 590548 73444
rect 564620 72380 564676 72436
rect 447692 72156 447748 72212
rect 559580 70812 559636 70868
rect 446012 69356 446068 69412
rect 563276 69244 563332 69300
rect 559468 67676 559524 67732
rect 444332 66444 444388 66500
rect 563164 66108 563220 66164
rect 27692 64988 27748 65044
rect 563052 64540 563108 64596
rect 449372 63532 449428 63588
rect 562940 62972 562996 63028
rect 574588 61404 574644 61460
rect 441084 60620 441140 60676
rect 577052 59948 577108 60004
rect 562828 59836 562884 59892
rect 427644 59612 427700 59668
rect 457660 59612 457716 59668
rect 567868 58828 567924 58884
rect 457660 57708 457716 57764
rect 564396 56700 564452 56756
rect 457772 54796 457828 54852
rect 419244 52892 419300 52948
rect 419244 51996 419300 52052
rect 4284 51100 4340 51156
rect 425852 50316 425908 50372
rect 562828 50316 562884 50372
rect 307468 50204 307524 50260
rect 314188 50204 314244 50260
rect 320908 50204 320964 50260
rect 362124 49532 362180 49588
rect 48524 48636 48580 48692
rect 267260 48524 267316 48580
rect 275660 48076 275716 48132
rect 267148 47852 267204 47908
rect 359212 44604 359268 44660
rect 411740 42812 411796 42868
rect 358988 41356 359044 41412
rect 362012 41244 362068 41300
rect 358652 41132 358708 41188
rect 358764 38108 358820 38164
rect 270508 36092 270564 36148
rect 275548 34860 275604 34916
rect 269612 34636 269668 34692
rect 269500 32956 269556 33012
rect 411852 32732 411908 32788
rect 411628 9212 411684 9268
rect 4172 8764 4228 8820
rect 291452 5964 291508 6020
rect 348572 4732 348628 4788
rect 51996 4508 52052 4564
rect 51884 4396 51940 4452
rect 579628 4172 579684 4228
rect 582988 4172 583044 4228
<< metal4 >>
rect -1916 598172 -1296 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 -1296 598172
rect -1916 598048 -1296 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 -1296 598048
rect -1916 597924 -1296 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 -1296 597924
rect -1916 597800 -1296 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 -1296 597800
rect -1916 586350 -1296 597744
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 -1296 586350
rect -1916 586226 -1296 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 -1296 586226
rect -1916 586102 -1296 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 -1296 586102
rect -1916 585978 -1296 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 -1296 585978
rect -1916 568350 -1296 585922
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 -1296 568350
rect -1916 568226 -1296 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 -1296 568226
rect -1916 568102 -1296 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 -1296 568102
rect -1916 567978 -1296 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 -1296 567978
rect -1916 550350 -1296 567922
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 -1296 550350
rect -1916 550226 -1296 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 -1296 550226
rect -1916 550102 -1296 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 -1296 550102
rect -1916 549978 -1296 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 -1296 549978
rect -1916 532350 -1296 549922
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 -1296 532350
rect -1916 532226 -1296 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 -1296 532226
rect -1916 532102 -1296 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 -1296 532102
rect -1916 531978 -1296 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 -1296 531978
rect -1916 514350 -1296 531922
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 -1296 514350
rect -1916 514226 -1296 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 -1296 514226
rect -1916 514102 -1296 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 -1296 514102
rect -1916 513978 -1296 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 -1296 513978
rect -1916 496350 -1296 513922
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 -1296 496350
rect -1916 496226 -1296 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 -1296 496226
rect -1916 496102 -1296 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 -1296 496102
rect -1916 495978 -1296 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 -1296 495978
rect -1916 478350 -1296 495922
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 -1296 478350
rect -1916 478226 -1296 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 -1296 478226
rect -1916 478102 -1296 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 -1296 478102
rect -1916 477978 -1296 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 -1296 477978
rect -1916 460350 -1296 477922
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 -1296 460350
rect -1916 460226 -1296 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 -1296 460226
rect -1916 460102 -1296 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 -1296 460102
rect -1916 459978 -1296 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 -1296 459978
rect -1916 442350 -1296 459922
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 -1296 442350
rect -1916 442226 -1296 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 -1296 442226
rect -1916 442102 -1296 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 -1296 442102
rect -1916 441978 -1296 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 -1296 441978
rect -1916 424350 -1296 441922
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 -1296 424350
rect -1916 424226 -1296 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 -1296 424226
rect -1916 424102 -1296 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 -1296 424102
rect -1916 423978 -1296 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 -1296 423978
rect -1916 406350 -1296 423922
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 -1296 406350
rect -1916 406226 -1296 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 -1296 406226
rect -1916 406102 -1296 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 -1296 406102
rect -1916 405978 -1296 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 -1296 405978
rect -1916 388350 -1296 405922
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 -1296 388350
rect -1916 388226 -1296 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 -1296 388226
rect -1916 388102 -1296 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 -1296 388102
rect -1916 387978 -1296 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 -1296 387978
rect -1916 370350 -1296 387922
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 -1296 370350
rect -1916 370226 -1296 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 -1296 370226
rect -1916 370102 -1296 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 -1296 370102
rect -1916 369978 -1296 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 -1296 369978
rect -1916 352350 -1296 369922
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 -1296 352350
rect -1916 352226 -1296 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 -1296 352226
rect -1916 352102 -1296 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 -1296 352102
rect -1916 351978 -1296 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 -1296 351978
rect -1916 334350 -1296 351922
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 -1296 334350
rect -1916 334226 -1296 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 -1296 334226
rect -1916 334102 -1296 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 -1296 334102
rect -1916 333978 -1296 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 -1296 333978
rect -1916 316350 -1296 333922
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 -1296 316350
rect -1916 316226 -1296 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 -1296 316226
rect -1916 316102 -1296 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 -1296 316102
rect -1916 315978 -1296 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 -1296 315978
rect -1916 298350 -1296 315922
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 -1296 298350
rect -1916 298226 -1296 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 -1296 298226
rect -1916 298102 -1296 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 -1296 298102
rect -1916 297978 -1296 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 -1296 297978
rect -1916 280350 -1296 297922
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 -1296 280350
rect -1916 280226 -1296 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 -1296 280226
rect -1916 280102 -1296 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 -1296 280102
rect -1916 279978 -1296 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 -1296 279978
rect -1916 262350 -1296 279922
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 -1296 262350
rect -1916 262226 -1296 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 -1296 262226
rect -1916 262102 -1296 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 -1296 262102
rect -1916 261978 -1296 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 -1296 261978
rect -1916 244350 -1296 261922
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 -1296 244350
rect -1916 244226 -1296 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 -1296 244226
rect -1916 244102 -1296 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 -1296 244102
rect -1916 243978 -1296 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 -1296 243978
rect -1916 226350 -1296 243922
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 -1296 226350
rect -1916 226226 -1296 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 -1296 226226
rect -1916 226102 -1296 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 -1296 226102
rect -1916 225978 -1296 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 -1296 225978
rect -1916 208350 -1296 225922
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 -1296 208350
rect -1916 208226 -1296 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 -1296 208226
rect -1916 208102 -1296 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 -1296 208102
rect -1916 207978 -1296 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 -1296 207978
rect -1916 190350 -1296 207922
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 -1296 190350
rect -1916 190226 -1296 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 -1296 190226
rect -1916 190102 -1296 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 -1296 190102
rect -1916 189978 -1296 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 -1296 189978
rect -1916 172350 -1296 189922
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 -1296 172350
rect -1916 172226 -1296 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 -1296 172226
rect -1916 172102 -1296 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 -1296 172102
rect -1916 171978 -1296 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 -1296 171978
rect -1916 154350 -1296 171922
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 -1296 154350
rect -1916 154226 -1296 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 -1296 154226
rect -1916 154102 -1296 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 -1296 154102
rect -1916 153978 -1296 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 -1296 153978
rect -1916 136350 -1296 153922
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 -1296 136350
rect -1916 136226 -1296 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 -1296 136226
rect -1916 136102 -1296 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 -1296 136102
rect -1916 135978 -1296 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 -1296 135978
rect -1916 118350 -1296 135922
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 -1296 118350
rect -1916 118226 -1296 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 -1296 118226
rect -1916 118102 -1296 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 -1296 118102
rect -1916 117978 -1296 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 -1296 117978
rect -1916 100350 -1296 117922
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 -1296 100350
rect -1916 100226 -1296 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 -1296 100226
rect -1916 100102 -1296 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 -1296 100102
rect -1916 99978 -1296 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 -1296 99978
rect -1916 82350 -1296 99922
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 -1296 82350
rect -1916 82226 -1296 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 -1296 82226
rect -1916 82102 -1296 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 -1296 82102
rect -1916 81978 -1296 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 -1296 81978
rect -1916 64350 -1296 81922
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 -1296 64350
rect -1916 64226 -1296 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 -1296 64226
rect -1916 64102 -1296 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 -1296 64102
rect -1916 63978 -1296 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 -1296 63978
rect -1916 46350 -1296 63922
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 -1296 46350
rect -1916 46226 -1296 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 -1296 46226
rect -1916 46102 -1296 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 -1296 46102
rect -1916 45978 -1296 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 -1296 45978
rect -1916 28350 -1296 45922
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 -1296 28350
rect -1916 28226 -1296 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 -1296 28226
rect -1916 28102 -1296 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 -1296 28102
rect -1916 27978 -1296 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 -1296 27978
rect -1916 10350 -1296 27922
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 -1296 10350
rect -1916 10226 -1296 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 -1296 10226
rect -1916 10102 -1296 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 -1296 10102
rect -1916 9978 -1296 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 -1296 9978
rect -1916 -1120 -1296 9922
rect -956 597212 -336 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 -336 597212
rect -956 597088 -336 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 -336 597088
rect -956 596964 -336 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 -336 596964
rect -956 596840 -336 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 -336 596840
rect -956 580350 -336 596784
rect -956 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 -336 580350
rect -956 580226 -336 580294
rect -956 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 -336 580226
rect -956 580102 -336 580170
rect -956 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 -336 580102
rect -956 579978 -336 580046
rect -956 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 -336 579978
rect -956 562350 -336 579922
rect -956 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 -336 562350
rect -956 562226 -336 562294
rect -956 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 -336 562226
rect -956 562102 -336 562170
rect -956 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 -336 562102
rect -956 561978 -336 562046
rect -956 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 -336 561978
rect -956 544350 -336 561922
rect 5418 597212 6038 598268
rect 5418 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 6038 597212
rect 5418 597088 6038 597156
rect 5418 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 6038 597088
rect 5418 596964 6038 597032
rect 5418 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 6038 596964
rect 5418 596840 6038 596908
rect 5418 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 6038 596840
rect 5418 580350 6038 596784
rect 5418 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 6038 580350
rect 5418 580226 6038 580294
rect 5418 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 6038 580226
rect 5418 580102 6038 580170
rect 5418 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 6038 580102
rect 5418 579978 6038 580046
rect 5418 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 6038 579978
rect 5418 562350 6038 579922
rect 5418 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 6038 562350
rect 5418 562226 6038 562294
rect 5418 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 6038 562226
rect 5418 562102 6038 562170
rect 5418 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 6038 562102
rect 5418 561978 6038 562046
rect 5418 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 6038 561978
rect -956 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 -336 544350
rect -956 544226 -336 544294
rect -956 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 -336 544226
rect -956 544102 -336 544170
rect -956 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 -336 544102
rect -956 543978 -336 544046
rect -956 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 -336 543978
rect -956 526350 -336 543922
rect -956 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 -336 526350
rect -956 526226 -336 526294
rect -956 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 -336 526226
rect -956 526102 -336 526170
rect -956 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 -336 526102
rect -956 525978 -336 526046
rect -956 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 -336 525978
rect -956 508350 -336 525922
rect -956 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 -336 508350
rect -956 508226 -336 508294
rect -956 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 -336 508226
rect -956 508102 -336 508170
rect -956 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 -336 508102
rect -956 507978 -336 508046
rect -956 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 -336 507978
rect -956 490350 -336 507922
rect -956 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 -336 490350
rect -956 490226 -336 490294
rect -956 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 -336 490226
rect -956 490102 -336 490170
rect -956 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 -336 490102
rect -956 489978 -336 490046
rect -956 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 -336 489978
rect -956 472350 -336 489922
rect 4172 558964 4228 558974
rect 4172 476308 4228 558908
rect 5418 544350 6038 561922
rect 9138 598172 9758 598268
rect 9138 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 9758 598172
rect 9138 598048 9758 598116
rect 9138 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 9758 598048
rect 9138 597924 9758 597992
rect 9138 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 9758 597924
rect 9138 597800 9758 597868
rect 9138 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 9758 597800
rect 9138 586350 9758 597744
rect 9138 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 9758 586350
rect 9138 586226 9758 586294
rect 9138 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 9758 586226
rect 9138 586102 9758 586170
rect 9138 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 9758 586102
rect 9138 585978 9758 586046
rect 9138 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 9758 585978
rect 9138 568350 9758 585922
rect 9138 568294 9234 568350
rect 9290 568294 9358 568350
rect 9414 568294 9482 568350
rect 9538 568294 9606 568350
rect 9662 568294 9758 568350
rect 9138 568226 9758 568294
rect 9138 568170 9234 568226
rect 9290 568170 9358 568226
rect 9414 568170 9482 568226
rect 9538 568170 9606 568226
rect 9662 568170 9758 568226
rect 9138 568102 9758 568170
rect 9138 568046 9234 568102
rect 9290 568046 9358 568102
rect 9414 568046 9482 568102
rect 9538 568046 9606 568102
rect 9662 568046 9758 568102
rect 9138 567978 9758 568046
rect 9138 567922 9234 567978
rect 9290 567922 9358 567978
rect 9414 567922 9482 567978
rect 9538 567922 9606 567978
rect 9662 567922 9758 567978
rect 9138 550350 9758 567922
rect 9138 550294 9234 550350
rect 9290 550294 9358 550350
rect 9414 550294 9482 550350
rect 9538 550294 9606 550350
rect 9662 550294 9758 550350
rect 9138 550226 9758 550294
rect 9138 550170 9234 550226
rect 9290 550170 9358 550226
rect 9414 550170 9482 550226
rect 9538 550170 9606 550226
rect 9662 550170 9758 550226
rect 9138 550102 9758 550170
rect 9138 550046 9234 550102
rect 9290 550046 9358 550102
rect 9414 550046 9482 550102
rect 9538 550046 9606 550102
rect 9662 550046 9758 550102
rect 9138 549978 9758 550046
rect 9138 549922 9234 549978
rect 9290 549922 9358 549978
rect 9414 549922 9482 549978
rect 9538 549922 9606 549978
rect 9662 549922 9758 549978
rect 5418 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 6038 544350
rect 5418 544226 6038 544294
rect 5418 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 6038 544226
rect 5418 544102 6038 544170
rect 5418 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 6038 544102
rect 5418 543978 6038 544046
rect 5418 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 6038 543978
rect 5418 526350 6038 543922
rect 5418 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 6038 526350
rect 5418 526226 6038 526294
rect 5418 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 6038 526226
rect 5418 526102 6038 526170
rect 5418 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 6038 526102
rect 5418 525978 6038 526046
rect 5418 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 6038 525978
rect 4172 476242 4228 476252
rect 4284 516628 4340 516638
rect -956 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 -336 472350
rect -956 472226 -336 472294
rect -956 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 -336 472226
rect -956 472102 -336 472170
rect -956 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 -336 472102
rect -956 471978 -336 472046
rect -956 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 -336 471978
rect -956 454350 -336 471922
rect 4284 469588 4340 516572
rect 4284 469522 4340 469532
rect 5418 508350 6038 525922
rect 5418 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 6038 508350
rect 5418 508226 6038 508294
rect 5418 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 6038 508226
rect 5418 508102 6038 508170
rect 5418 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 6038 508102
rect 5418 507978 6038 508046
rect 5418 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 6038 507978
rect 5418 490350 6038 507922
rect 5418 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 6038 490350
rect 5418 490226 6038 490294
rect 5418 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 6038 490226
rect 5418 490102 6038 490170
rect 5418 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 6038 490102
rect 5418 489978 6038 490046
rect 5418 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 6038 489978
rect 5418 472350 6038 489922
rect 5418 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 6038 472350
rect 5418 472226 6038 472294
rect 5418 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 6038 472226
rect 5418 472102 6038 472170
rect 5418 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 6038 472102
rect 5418 471978 6038 472046
rect 5418 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 6038 471978
rect -956 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 -336 454350
rect -956 454226 -336 454294
rect -956 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 -336 454226
rect -956 454102 -336 454170
rect -956 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 -336 454102
rect -956 453978 -336 454046
rect -956 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 -336 453978
rect -956 436350 -336 453922
rect -956 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 -336 436350
rect -956 436226 -336 436294
rect -956 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 -336 436226
rect -956 436102 -336 436170
rect -956 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 -336 436102
rect -956 435978 -336 436046
rect -956 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 -336 435978
rect -956 418350 -336 435922
rect -956 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 -336 418350
rect -956 418226 -336 418294
rect -956 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 -336 418226
rect -956 418102 -336 418170
rect -956 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 -336 418102
rect -956 417978 -336 418046
rect -956 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 -336 417978
rect -956 400350 -336 417922
rect -956 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 -336 400350
rect -956 400226 -336 400294
rect -956 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 -336 400226
rect -956 400102 -336 400170
rect -956 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 -336 400102
rect -956 399978 -336 400046
rect -956 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 -336 399978
rect -956 382350 -336 399922
rect 5418 454350 6038 471922
rect 5418 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 6038 454350
rect 5418 454226 6038 454294
rect 5418 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 6038 454226
rect 5418 454102 6038 454170
rect 5418 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 6038 454102
rect 5418 453978 6038 454046
rect 5418 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 6038 453978
rect 5418 436350 6038 453922
rect 5418 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 6038 436350
rect 5418 436226 6038 436294
rect 5418 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 6038 436226
rect 5418 436102 6038 436170
rect 5418 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 6038 436102
rect 5418 435978 6038 436046
rect 5418 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 6038 435978
rect 5418 418350 6038 435922
rect 5418 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 6038 418350
rect 5418 418226 6038 418294
rect 5418 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 6038 418226
rect 5418 418102 6038 418170
rect 5418 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 6038 418102
rect 5418 417978 6038 418046
rect 5418 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 6038 417978
rect 5418 400350 6038 417922
rect 7532 544852 7588 544862
rect 7532 409078 7588 544796
rect 7532 409012 7588 409022
rect 9138 532350 9758 549922
rect 9138 532294 9234 532350
rect 9290 532294 9358 532350
rect 9414 532294 9482 532350
rect 9538 532294 9606 532350
rect 9662 532294 9758 532350
rect 9138 532226 9758 532294
rect 9138 532170 9234 532226
rect 9290 532170 9358 532226
rect 9414 532170 9482 532226
rect 9538 532170 9606 532226
rect 9662 532170 9758 532226
rect 9138 532102 9758 532170
rect 9138 532046 9234 532102
rect 9290 532046 9358 532102
rect 9414 532046 9482 532102
rect 9538 532046 9606 532102
rect 9662 532046 9758 532102
rect 9138 531978 9758 532046
rect 9138 531922 9234 531978
rect 9290 531922 9358 531978
rect 9414 531922 9482 531978
rect 9538 531922 9606 531978
rect 9662 531922 9758 531978
rect 9138 514350 9758 531922
rect 9138 514294 9234 514350
rect 9290 514294 9358 514350
rect 9414 514294 9482 514350
rect 9538 514294 9606 514350
rect 9662 514294 9758 514350
rect 9138 514226 9758 514294
rect 9138 514170 9234 514226
rect 9290 514170 9358 514226
rect 9414 514170 9482 514226
rect 9538 514170 9606 514226
rect 9662 514170 9758 514226
rect 9138 514102 9758 514170
rect 9138 514046 9234 514102
rect 9290 514046 9358 514102
rect 9414 514046 9482 514102
rect 9538 514046 9606 514102
rect 9662 514046 9758 514102
rect 9138 513978 9758 514046
rect 9138 513922 9234 513978
rect 9290 513922 9358 513978
rect 9414 513922 9482 513978
rect 9538 513922 9606 513978
rect 9662 513922 9758 513978
rect 9138 496350 9758 513922
rect 9138 496294 9234 496350
rect 9290 496294 9358 496350
rect 9414 496294 9482 496350
rect 9538 496294 9606 496350
rect 9662 496294 9758 496350
rect 9138 496226 9758 496294
rect 9138 496170 9234 496226
rect 9290 496170 9358 496226
rect 9414 496170 9482 496226
rect 9538 496170 9606 496226
rect 9662 496170 9758 496226
rect 9138 496102 9758 496170
rect 9138 496046 9234 496102
rect 9290 496046 9358 496102
rect 9414 496046 9482 496102
rect 9538 496046 9606 496102
rect 9662 496046 9758 496102
rect 9138 495978 9758 496046
rect 9138 495922 9234 495978
rect 9290 495922 9358 495978
rect 9414 495922 9482 495978
rect 9538 495922 9606 495978
rect 9662 495922 9758 495978
rect 9138 478350 9758 495922
rect 9138 478294 9234 478350
rect 9290 478294 9358 478350
rect 9414 478294 9482 478350
rect 9538 478294 9606 478350
rect 9662 478294 9758 478350
rect 9138 478226 9758 478294
rect 9138 478170 9234 478226
rect 9290 478170 9358 478226
rect 9414 478170 9482 478226
rect 9538 478170 9606 478226
rect 9662 478170 9758 478226
rect 9138 478102 9758 478170
rect 9138 478046 9234 478102
rect 9290 478046 9358 478102
rect 9414 478046 9482 478102
rect 9538 478046 9606 478102
rect 9662 478046 9758 478102
rect 9138 477978 9758 478046
rect 9138 477922 9234 477978
rect 9290 477922 9358 477978
rect 9414 477922 9482 477978
rect 9538 477922 9606 477978
rect 9662 477922 9758 477978
rect 9138 460350 9758 477922
rect 9138 460294 9234 460350
rect 9290 460294 9358 460350
rect 9414 460294 9482 460350
rect 9538 460294 9606 460350
rect 9662 460294 9758 460350
rect 9138 460226 9758 460294
rect 9138 460170 9234 460226
rect 9290 460170 9358 460226
rect 9414 460170 9482 460226
rect 9538 460170 9606 460226
rect 9662 460170 9758 460226
rect 9138 460102 9758 460170
rect 9138 460046 9234 460102
rect 9290 460046 9358 460102
rect 9414 460046 9482 460102
rect 9538 460046 9606 460102
rect 9662 460046 9758 460102
rect 9138 459978 9758 460046
rect 9138 459922 9234 459978
rect 9290 459922 9358 459978
rect 9414 459922 9482 459978
rect 9538 459922 9606 459978
rect 9662 459922 9758 459978
rect 9138 442350 9758 459922
rect 9138 442294 9234 442350
rect 9290 442294 9358 442350
rect 9414 442294 9482 442350
rect 9538 442294 9606 442350
rect 9662 442294 9758 442350
rect 9138 442226 9758 442294
rect 9138 442170 9234 442226
rect 9290 442170 9358 442226
rect 9414 442170 9482 442226
rect 9538 442170 9606 442226
rect 9662 442170 9758 442226
rect 9138 442102 9758 442170
rect 9138 442046 9234 442102
rect 9290 442046 9358 442102
rect 9414 442046 9482 442102
rect 9538 442046 9606 442102
rect 9662 442046 9758 442102
rect 9138 441978 9758 442046
rect 9138 441922 9234 441978
rect 9290 441922 9358 441978
rect 9414 441922 9482 441978
rect 9538 441922 9606 441978
rect 9662 441922 9758 441978
rect 9138 424350 9758 441922
rect 9138 424294 9234 424350
rect 9290 424294 9358 424350
rect 9414 424294 9482 424350
rect 9538 424294 9606 424350
rect 9662 424294 9758 424350
rect 9138 424226 9758 424294
rect 9138 424170 9234 424226
rect 9290 424170 9358 424226
rect 9414 424170 9482 424226
rect 9538 424170 9606 424226
rect 9662 424170 9758 424226
rect 9138 424102 9758 424170
rect 9138 424046 9234 424102
rect 9290 424046 9358 424102
rect 9414 424046 9482 424102
rect 9538 424046 9606 424102
rect 9662 424046 9758 424102
rect 9138 423978 9758 424046
rect 9138 423922 9234 423978
rect 9290 423922 9358 423978
rect 9414 423922 9482 423978
rect 9538 423922 9606 423978
rect 9662 423922 9758 423978
rect 5418 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 6038 400350
rect 5418 400226 6038 400294
rect 5418 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 6038 400226
rect 5418 400102 6038 400170
rect 5418 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 6038 400102
rect 5418 399978 6038 400046
rect 5418 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 6038 399978
rect -956 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 -336 382350
rect -956 382226 -336 382294
rect -956 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 -336 382226
rect -956 382102 -336 382170
rect -956 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 -336 382102
rect -956 381978 -336 382046
rect -956 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 -336 381978
rect -956 364350 -336 381922
rect 4172 389620 4228 389630
rect 4172 380548 4228 389564
rect 4172 380482 4228 380492
rect 5418 382350 6038 399922
rect 9138 406350 9758 423922
rect 9138 406294 9234 406350
rect 9290 406294 9358 406350
rect 9414 406294 9482 406350
rect 9538 406294 9606 406350
rect 9662 406294 9758 406350
rect 9138 406226 9758 406294
rect 9138 406170 9234 406226
rect 9290 406170 9358 406226
rect 9414 406170 9482 406226
rect 9538 406170 9606 406226
rect 9662 406170 9758 406226
rect 9138 406102 9758 406170
rect 9138 406046 9234 406102
rect 9290 406046 9358 406102
rect 9414 406046 9482 406102
rect 9538 406046 9606 406102
rect 9662 406046 9758 406102
rect 9138 405978 9758 406046
rect 9138 405922 9234 405978
rect 9290 405922 9358 405978
rect 9414 405922 9482 405978
rect 9538 405922 9606 405978
rect 9662 405922 9758 405978
rect 9138 388350 9758 405922
rect 9138 388294 9234 388350
rect 9290 388294 9358 388350
rect 9414 388294 9482 388350
rect 9538 388294 9606 388350
rect 9662 388294 9758 388350
rect 9138 388226 9758 388294
rect 9138 388170 9234 388226
rect 9290 388170 9358 388226
rect 9414 388170 9482 388226
rect 9538 388170 9606 388226
rect 9662 388170 9758 388226
rect 9138 388102 9758 388170
rect 9138 388046 9234 388102
rect 9290 388046 9358 388102
rect 9414 388046 9482 388102
rect 9538 388046 9606 388102
rect 9662 388046 9758 388102
rect 9138 387978 9758 388046
rect 9138 387922 9234 387978
rect 9290 387922 9358 387978
rect 9414 387922 9482 387978
rect 9538 387922 9606 387978
rect 9662 387922 9758 387978
rect 5418 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 6038 382350
rect 5418 382226 6038 382294
rect 5418 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 6038 382226
rect 5418 382102 6038 382170
rect 5418 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 6038 382102
rect 5418 381978 6038 382046
rect 5418 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 6038 381978
rect -956 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 -336 364350
rect -956 364226 -336 364294
rect -956 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 -336 364226
rect -956 364102 -336 364170
rect -956 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 -336 364102
rect -956 363978 -336 364046
rect -956 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 -336 363978
rect -956 346350 -336 363922
rect 5418 364350 6038 381922
rect 5418 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 6038 364350
rect 5418 364226 6038 364294
rect 5418 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 6038 364226
rect 5418 364102 6038 364170
rect 5418 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 6038 364102
rect 5418 363978 6038 364046
rect 5418 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 6038 363978
rect -956 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 -336 346350
rect -956 346226 -336 346294
rect -956 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 -336 346226
rect -956 346102 -336 346170
rect -956 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 -336 346102
rect -956 345978 -336 346046
rect -956 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 -336 345978
rect -956 328350 -336 345922
rect 4172 347284 4228 347294
rect 4172 345268 4228 347228
rect 4172 345202 4228 345212
rect 5418 346350 6038 363922
rect 5418 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 6038 346350
rect 5418 346226 6038 346294
rect 5418 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 6038 346226
rect 5418 346102 6038 346170
rect 5418 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 6038 346102
rect 5418 345978 6038 346046
rect 5418 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 6038 345978
rect -956 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 -336 328350
rect -956 328226 -336 328294
rect -956 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 -336 328226
rect -956 328102 -336 328170
rect -956 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 -336 328102
rect -956 327978 -336 328046
rect -956 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 -336 327978
rect -956 310350 -336 327922
rect -956 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 -336 310350
rect -956 310226 -336 310294
rect -956 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 -336 310226
rect -956 310102 -336 310170
rect -956 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 -336 310102
rect -956 309978 -336 310046
rect -956 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 -336 309978
rect -956 292350 -336 309922
rect 5418 328350 6038 345922
rect 5418 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 6038 328350
rect 5418 328226 6038 328294
rect 5418 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 6038 328226
rect 5418 328102 6038 328170
rect 5418 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 6038 328102
rect 5418 327978 6038 328046
rect 5418 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 6038 327978
rect 5418 310350 6038 327922
rect 5418 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 6038 310350
rect 5418 310226 6038 310294
rect 5418 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 6038 310226
rect 5418 310102 6038 310170
rect 5418 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 6038 310102
rect 5418 309978 6038 310046
rect 5418 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 6038 309978
rect -956 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 -336 292350
rect -956 292226 -336 292294
rect -956 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 -336 292226
rect -956 292102 -336 292170
rect -956 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 -336 292102
rect -956 291978 -336 292046
rect -956 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 -336 291978
rect -956 274350 -336 291922
rect -956 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 -336 274350
rect -956 274226 -336 274294
rect -956 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 -336 274226
rect -956 274102 -336 274170
rect -956 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 -336 274102
rect -956 273978 -336 274046
rect -956 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 -336 273978
rect -956 256350 -336 273922
rect -956 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 -336 256350
rect -956 256226 -336 256294
rect -956 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 -336 256226
rect -956 256102 -336 256170
rect -956 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 -336 256102
rect -956 255978 -336 256046
rect -956 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 -336 255978
rect -956 238350 -336 255922
rect 4172 305844 4228 305854
rect 4060 248500 4116 248510
rect 4060 247078 4116 248444
rect 4060 247012 4116 247022
rect -956 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 -336 238350
rect -956 238226 -336 238294
rect -956 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 -336 238226
rect -956 238102 -336 238170
rect -956 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 -336 238102
rect -956 237978 -336 238046
rect -956 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 -336 237978
rect -956 220350 -336 237922
rect -956 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 -336 220350
rect -956 220226 -336 220294
rect -956 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 -336 220226
rect -956 220102 -336 220170
rect -956 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 -336 220102
rect -956 219978 -336 220046
rect -956 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 -336 219978
rect -956 202350 -336 219922
rect 4172 208348 4228 305788
rect -956 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 -336 202350
rect -956 202226 -336 202294
rect -956 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 -336 202226
rect -956 202102 -336 202170
rect -956 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 -336 202102
rect -956 201978 -336 202046
rect -956 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 -336 201978
rect -956 184350 -336 201922
rect 4060 208292 4228 208348
rect 4284 304724 4340 304734
rect 4060 196588 4116 208292
rect 4172 206578 4228 206588
rect 4172 206388 4228 206522
rect 4172 206322 4228 206332
rect 4060 196532 4228 196588
rect -956 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 -336 184350
rect -956 184226 -336 184294
rect -956 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 -336 184226
rect -956 184102 -336 184170
rect -956 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 -336 184102
rect -956 183978 -336 184046
rect -956 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 -336 183978
rect -956 166350 -336 183922
rect 4172 173068 4228 196532
rect -956 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 -336 166350
rect -956 166226 -336 166294
rect -956 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 -336 166226
rect -956 166102 -336 166170
rect -956 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 -336 166102
rect -956 165978 -336 166046
rect -956 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 -336 165978
rect -956 148350 -336 165922
rect 4060 173012 4228 173068
rect 4060 161308 4116 173012
rect 4172 164638 4228 164648
rect 4172 164052 4228 164582
rect 4172 163986 4228 163996
rect 4060 161252 4228 161308
rect -956 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 -336 148350
rect -956 148226 -336 148294
rect -956 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 -336 148226
rect -956 148102 -336 148170
rect -956 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 -336 148102
rect -956 147978 -336 148046
rect -956 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 -336 147978
rect -956 130350 -336 147922
rect -956 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 -336 130350
rect -956 130226 -336 130294
rect -956 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 -336 130226
rect -956 130102 -336 130170
rect -956 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 -336 130102
rect -956 129978 -336 130046
rect -956 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 -336 129978
rect -956 112350 -336 129922
rect -956 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 -336 112350
rect -956 112226 -336 112294
rect -956 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 -336 112226
rect -956 112102 -336 112170
rect -956 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 -336 112102
rect -956 111978 -336 112046
rect -956 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 -336 111978
rect -956 94350 -336 111922
rect -956 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 -336 94350
rect -956 94226 -336 94294
rect -956 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 -336 94226
rect -956 94102 -336 94170
rect -956 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 -336 94102
rect -956 93978 -336 94046
rect -956 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 -336 93978
rect -956 76350 -336 93922
rect -956 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 -336 76350
rect -956 76226 -336 76294
rect -956 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 -336 76226
rect -956 76102 -336 76170
rect -956 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 -336 76102
rect -956 75978 -336 76046
rect -956 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 -336 75978
rect -956 58350 -336 75922
rect -956 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 -336 58350
rect -956 58226 -336 58294
rect -956 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 -336 58226
rect -956 58102 -336 58170
rect -956 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 -336 58102
rect -956 57978 -336 58046
rect -956 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 -336 57978
rect -956 40350 -336 57922
rect -956 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 -336 40350
rect -956 40226 -336 40294
rect -956 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 -336 40226
rect -956 40102 -336 40170
rect -956 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 -336 40102
rect -956 39978 -336 40046
rect -956 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 -336 39978
rect -956 22350 -336 39922
rect -956 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 -336 22350
rect -956 22226 -336 22294
rect -956 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 -336 22226
rect -956 22102 -336 22170
rect -956 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 -336 22102
rect -956 21978 -336 22046
rect -956 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 -336 21978
rect -956 4350 -336 21922
rect 4172 8820 4228 161252
rect 4284 51156 4340 304668
rect 4284 51090 4340 51100
rect 5418 292350 6038 309922
rect 5418 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 6038 292350
rect 5418 292226 6038 292294
rect 5418 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 6038 292226
rect 5418 292102 6038 292170
rect 5418 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 6038 292102
rect 5418 291978 6038 292046
rect 5418 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 6038 291978
rect 5418 274350 6038 291922
rect 5418 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 6038 274350
rect 5418 274226 6038 274294
rect 5418 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 6038 274226
rect 5418 274102 6038 274170
rect 5418 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 6038 274102
rect 5418 273978 6038 274046
rect 5418 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 6038 273978
rect 5418 256350 6038 273922
rect 5418 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 6038 256350
rect 5418 256226 6038 256294
rect 5418 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 6038 256226
rect 5418 256102 6038 256170
rect 5418 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 6038 256102
rect 5418 255978 6038 256046
rect 5418 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 6038 255978
rect 5418 238350 6038 255922
rect 5418 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 6038 238350
rect 5418 238226 6038 238294
rect 5418 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 6038 238226
rect 5418 238102 6038 238170
rect 5418 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 6038 238102
rect 5418 237978 6038 238046
rect 5418 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 6038 237978
rect 5418 220350 6038 237922
rect 5418 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 6038 220350
rect 5418 220226 6038 220294
rect 5418 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 6038 220226
rect 5418 220102 6038 220170
rect 5418 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 6038 220102
rect 5418 219978 6038 220046
rect 5418 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 6038 219978
rect 5418 202350 6038 219922
rect 5418 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 6038 202350
rect 5418 202226 6038 202294
rect 5418 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 6038 202226
rect 5418 202102 6038 202170
rect 5418 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 6038 202102
rect 5418 201978 6038 202046
rect 5418 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 6038 201978
rect 5418 184350 6038 201922
rect 5418 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 6038 184350
rect 5418 184226 6038 184294
rect 5418 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 6038 184226
rect 5418 184102 6038 184170
rect 5418 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 6038 184102
rect 5418 183978 6038 184046
rect 5418 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 6038 183978
rect 5418 166350 6038 183922
rect 5418 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 6038 166350
rect 5418 166226 6038 166294
rect 5418 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 6038 166226
rect 5418 166102 6038 166170
rect 5418 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 6038 166102
rect 5418 165978 6038 166046
rect 5418 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 6038 165978
rect 5418 148350 6038 165922
rect 7532 385498 7588 385508
rect 7532 149940 7588 385442
rect 7532 149874 7588 149884
rect 9138 370350 9758 387922
rect 36138 597212 36758 598268
rect 36138 597156 36234 597212
rect 36290 597156 36358 597212
rect 36414 597156 36482 597212
rect 36538 597156 36606 597212
rect 36662 597156 36758 597212
rect 36138 597088 36758 597156
rect 36138 597032 36234 597088
rect 36290 597032 36358 597088
rect 36414 597032 36482 597088
rect 36538 597032 36606 597088
rect 36662 597032 36758 597088
rect 36138 596964 36758 597032
rect 36138 596908 36234 596964
rect 36290 596908 36358 596964
rect 36414 596908 36482 596964
rect 36538 596908 36606 596964
rect 36662 596908 36758 596964
rect 36138 596840 36758 596908
rect 36138 596784 36234 596840
rect 36290 596784 36358 596840
rect 36414 596784 36482 596840
rect 36538 596784 36606 596840
rect 36662 596784 36758 596840
rect 36138 580350 36758 596784
rect 36138 580294 36234 580350
rect 36290 580294 36358 580350
rect 36414 580294 36482 580350
rect 36538 580294 36606 580350
rect 36662 580294 36758 580350
rect 36138 580226 36758 580294
rect 36138 580170 36234 580226
rect 36290 580170 36358 580226
rect 36414 580170 36482 580226
rect 36538 580170 36606 580226
rect 36662 580170 36758 580226
rect 36138 580102 36758 580170
rect 36138 580046 36234 580102
rect 36290 580046 36358 580102
rect 36414 580046 36482 580102
rect 36538 580046 36606 580102
rect 36662 580046 36758 580102
rect 36138 579978 36758 580046
rect 36138 579922 36234 579978
rect 36290 579922 36358 579978
rect 36414 579922 36482 579978
rect 36538 579922 36606 579978
rect 36662 579922 36758 579978
rect 36138 562350 36758 579922
rect 36138 562294 36234 562350
rect 36290 562294 36358 562350
rect 36414 562294 36482 562350
rect 36538 562294 36606 562350
rect 36662 562294 36758 562350
rect 36138 562226 36758 562294
rect 36138 562170 36234 562226
rect 36290 562170 36358 562226
rect 36414 562170 36482 562226
rect 36538 562170 36606 562226
rect 36662 562170 36758 562226
rect 36138 562102 36758 562170
rect 36138 562046 36234 562102
rect 36290 562046 36358 562102
rect 36414 562046 36482 562102
rect 36538 562046 36606 562102
rect 36662 562046 36758 562102
rect 36138 561978 36758 562046
rect 36138 561922 36234 561978
rect 36290 561922 36358 561978
rect 36414 561922 36482 561978
rect 36538 561922 36606 561978
rect 36662 561922 36758 561978
rect 36138 544350 36758 561922
rect 36138 544294 36234 544350
rect 36290 544294 36358 544350
rect 36414 544294 36482 544350
rect 36538 544294 36606 544350
rect 36662 544294 36758 544350
rect 36138 544226 36758 544294
rect 36138 544170 36234 544226
rect 36290 544170 36358 544226
rect 36414 544170 36482 544226
rect 36538 544170 36606 544226
rect 36662 544170 36758 544226
rect 36138 544102 36758 544170
rect 36138 544046 36234 544102
rect 36290 544046 36358 544102
rect 36414 544046 36482 544102
rect 36538 544046 36606 544102
rect 36662 544046 36758 544102
rect 36138 543978 36758 544046
rect 36138 543922 36234 543978
rect 36290 543922 36358 543978
rect 36414 543922 36482 543978
rect 36538 543922 36606 543978
rect 36662 543922 36758 543978
rect 36138 526350 36758 543922
rect 36138 526294 36234 526350
rect 36290 526294 36358 526350
rect 36414 526294 36482 526350
rect 36538 526294 36606 526350
rect 36662 526294 36758 526350
rect 36138 526226 36758 526294
rect 36138 526170 36234 526226
rect 36290 526170 36358 526226
rect 36414 526170 36482 526226
rect 36538 526170 36606 526226
rect 36662 526170 36758 526226
rect 36138 526102 36758 526170
rect 36138 526046 36234 526102
rect 36290 526046 36358 526102
rect 36414 526046 36482 526102
rect 36538 526046 36606 526102
rect 36662 526046 36758 526102
rect 36138 525978 36758 526046
rect 36138 525922 36234 525978
rect 36290 525922 36358 525978
rect 36414 525922 36482 525978
rect 36538 525922 36606 525978
rect 36662 525922 36758 525978
rect 36138 508350 36758 525922
rect 36138 508294 36234 508350
rect 36290 508294 36358 508350
rect 36414 508294 36482 508350
rect 36538 508294 36606 508350
rect 36662 508294 36758 508350
rect 36138 508226 36758 508294
rect 36138 508170 36234 508226
rect 36290 508170 36358 508226
rect 36414 508170 36482 508226
rect 36538 508170 36606 508226
rect 36662 508170 36758 508226
rect 36138 508102 36758 508170
rect 36138 508046 36234 508102
rect 36290 508046 36358 508102
rect 36414 508046 36482 508102
rect 36538 508046 36606 508102
rect 36662 508046 36758 508102
rect 36138 507978 36758 508046
rect 36138 507922 36234 507978
rect 36290 507922 36358 507978
rect 36414 507922 36482 507978
rect 36538 507922 36606 507978
rect 36662 507922 36758 507978
rect 36138 490350 36758 507922
rect 36138 490294 36234 490350
rect 36290 490294 36358 490350
rect 36414 490294 36482 490350
rect 36538 490294 36606 490350
rect 36662 490294 36758 490350
rect 36138 490226 36758 490294
rect 36138 490170 36234 490226
rect 36290 490170 36358 490226
rect 36414 490170 36482 490226
rect 36538 490170 36606 490226
rect 36662 490170 36758 490226
rect 36138 490102 36758 490170
rect 36138 490046 36234 490102
rect 36290 490046 36358 490102
rect 36414 490046 36482 490102
rect 36538 490046 36606 490102
rect 36662 490046 36758 490102
rect 36138 489978 36758 490046
rect 36138 489922 36234 489978
rect 36290 489922 36358 489978
rect 36414 489922 36482 489978
rect 36538 489922 36606 489978
rect 36662 489922 36758 489978
rect 36138 472350 36758 489922
rect 36138 472294 36234 472350
rect 36290 472294 36358 472350
rect 36414 472294 36482 472350
rect 36538 472294 36606 472350
rect 36662 472294 36758 472350
rect 36138 472226 36758 472294
rect 36138 472170 36234 472226
rect 36290 472170 36358 472226
rect 36414 472170 36482 472226
rect 36538 472170 36606 472226
rect 36662 472170 36758 472226
rect 36138 472102 36758 472170
rect 36138 472046 36234 472102
rect 36290 472046 36358 472102
rect 36414 472046 36482 472102
rect 36538 472046 36606 472102
rect 36662 472046 36758 472102
rect 36138 471978 36758 472046
rect 36138 471922 36234 471978
rect 36290 471922 36358 471978
rect 36414 471922 36482 471978
rect 36538 471922 36606 471978
rect 36662 471922 36758 471978
rect 36138 454350 36758 471922
rect 36138 454294 36234 454350
rect 36290 454294 36358 454350
rect 36414 454294 36482 454350
rect 36538 454294 36606 454350
rect 36662 454294 36758 454350
rect 36138 454226 36758 454294
rect 36138 454170 36234 454226
rect 36290 454170 36358 454226
rect 36414 454170 36482 454226
rect 36538 454170 36606 454226
rect 36662 454170 36758 454226
rect 36138 454102 36758 454170
rect 36138 454046 36234 454102
rect 36290 454046 36358 454102
rect 36414 454046 36482 454102
rect 36538 454046 36606 454102
rect 36662 454046 36758 454102
rect 36138 453978 36758 454046
rect 36138 453922 36234 453978
rect 36290 453922 36358 453978
rect 36414 453922 36482 453978
rect 36538 453922 36606 453978
rect 36662 453922 36758 453978
rect 36138 436350 36758 453922
rect 36138 436294 36234 436350
rect 36290 436294 36358 436350
rect 36414 436294 36482 436350
rect 36538 436294 36606 436350
rect 36662 436294 36758 436350
rect 36138 436226 36758 436294
rect 36138 436170 36234 436226
rect 36290 436170 36358 436226
rect 36414 436170 36482 436226
rect 36538 436170 36606 436226
rect 36662 436170 36758 436226
rect 36138 436102 36758 436170
rect 36138 436046 36234 436102
rect 36290 436046 36358 436102
rect 36414 436046 36482 436102
rect 36538 436046 36606 436102
rect 36662 436046 36758 436102
rect 36138 435978 36758 436046
rect 36138 435922 36234 435978
rect 36290 435922 36358 435978
rect 36414 435922 36482 435978
rect 36538 435922 36606 435978
rect 36662 435922 36758 435978
rect 36138 418350 36758 435922
rect 36138 418294 36234 418350
rect 36290 418294 36358 418350
rect 36414 418294 36482 418350
rect 36538 418294 36606 418350
rect 36662 418294 36758 418350
rect 36138 418226 36758 418294
rect 36138 418170 36234 418226
rect 36290 418170 36358 418226
rect 36414 418170 36482 418226
rect 36538 418170 36606 418226
rect 36662 418170 36758 418226
rect 36138 418102 36758 418170
rect 36138 418046 36234 418102
rect 36290 418046 36358 418102
rect 36414 418046 36482 418102
rect 36538 418046 36606 418102
rect 36662 418046 36758 418102
rect 36138 417978 36758 418046
rect 36138 417922 36234 417978
rect 36290 417922 36358 417978
rect 36414 417922 36482 417978
rect 36538 417922 36606 417978
rect 36662 417922 36758 417978
rect 36138 400350 36758 417922
rect 36138 400294 36234 400350
rect 36290 400294 36358 400350
rect 36414 400294 36482 400350
rect 36538 400294 36606 400350
rect 36662 400294 36758 400350
rect 36138 400226 36758 400294
rect 36138 400170 36234 400226
rect 36290 400170 36358 400226
rect 36414 400170 36482 400226
rect 36538 400170 36606 400226
rect 36662 400170 36758 400226
rect 36138 400102 36758 400170
rect 36138 400046 36234 400102
rect 36290 400046 36358 400102
rect 36414 400046 36482 400102
rect 36538 400046 36606 400102
rect 36662 400046 36758 400102
rect 36138 399978 36758 400046
rect 36138 399922 36234 399978
rect 36290 399922 36358 399978
rect 36414 399922 36482 399978
rect 36538 399922 36606 399978
rect 36662 399922 36758 399978
rect 9138 370294 9234 370350
rect 9290 370294 9358 370350
rect 9414 370294 9482 370350
rect 9538 370294 9606 370350
rect 9662 370294 9758 370350
rect 9138 370226 9758 370294
rect 9138 370170 9234 370226
rect 9290 370170 9358 370226
rect 9414 370170 9482 370226
rect 9538 370170 9606 370226
rect 9662 370170 9758 370226
rect 9138 370102 9758 370170
rect 9138 370046 9234 370102
rect 9290 370046 9358 370102
rect 9414 370046 9482 370102
rect 9538 370046 9606 370102
rect 9662 370046 9758 370102
rect 9138 369978 9758 370046
rect 9138 369922 9234 369978
rect 9290 369922 9358 369978
rect 9414 369922 9482 369978
rect 9538 369922 9606 369978
rect 9662 369922 9758 369978
rect 9138 352350 9758 369922
rect 9138 352294 9234 352350
rect 9290 352294 9358 352350
rect 9414 352294 9482 352350
rect 9538 352294 9606 352350
rect 9662 352294 9758 352350
rect 9138 352226 9758 352294
rect 9138 352170 9234 352226
rect 9290 352170 9358 352226
rect 9414 352170 9482 352226
rect 9538 352170 9606 352226
rect 9662 352170 9758 352226
rect 9138 352102 9758 352170
rect 9138 352046 9234 352102
rect 9290 352046 9358 352102
rect 9414 352046 9482 352102
rect 9538 352046 9606 352102
rect 9662 352046 9758 352102
rect 9138 351978 9758 352046
rect 9138 351922 9234 351978
rect 9290 351922 9358 351978
rect 9414 351922 9482 351978
rect 9538 351922 9606 351978
rect 9662 351922 9758 351978
rect 9138 334350 9758 351922
rect 9138 334294 9234 334350
rect 9290 334294 9358 334350
rect 9414 334294 9482 334350
rect 9538 334294 9606 334350
rect 9662 334294 9758 334350
rect 9138 334226 9758 334294
rect 9138 334170 9234 334226
rect 9290 334170 9358 334226
rect 9414 334170 9482 334226
rect 9538 334170 9606 334226
rect 9662 334170 9758 334226
rect 9138 334102 9758 334170
rect 9138 334046 9234 334102
rect 9290 334046 9358 334102
rect 9414 334046 9482 334102
rect 9538 334046 9606 334102
rect 9662 334046 9758 334102
rect 9138 333978 9758 334046
rect 9138 333922 9234 333978
rect 9290 333922 9358 333978
rect 9414 333922 9482 333978
rect 9538 333922 9606 333978
rect 9662 333922 9758 333978
rect 9138 316350 9758 333922
rect 9138 316294 9234 316350
rect 9290 316294 9358 316350
rect 9414 316294 9482 316350
rect 9538 316294 9606 316350
rect 9662 316294 9758 316350
rect 9138 316226 9758 316294
rect 9138 316170 9234 316226
rect 9290 316170 9358 316226
rect 9414 316170 9482 316226
rect 9538 316170 9606 316226
rect 9662 316170 9758 316226
rect 9138 316102 9758 316170
rect 9138 316046 9234 316102
rect 9290 316046 9358 316102
rect 9414 316046 9482 316102
rect 9538 316046 9606 316102
rect 9662 316046 9758 316102
rect 9138 315978 9758 316046
rect 9138 315922 9234 315978
rect 9290 315922 9358 315978
rect 9414 315922 9482 315978
rect 9538 315922 9606 315978
rect 9662 315922 9758 315978
rect 9138 298350 9758 315922
rect 27692 385318 27748 385328
rect 12572 300244 12628 300254
rect 9138 298294 9234 298350
rect 9290 298294 9358 298350
rect 9414 298294 9482 298350
rect 9538 298294 9606 298350
rect 9662 298294 9758 298350
rect 9138 298226 9758 298294
rect 9138 298170 9234 298226
rect 9290 298170 9358 298226
rect 9414 298170 9482 298226
rect 9538 298170 9606 298226
rect 9662 298170 9758 298226
rect 9138 298102 9758 298170
rect 9138 298046 9234 298102
rect 9290 298046 9358 298102
rect 9414 298046 9482 298102
rect 9538 298046 9606 298102
rect 9662 298046 9758 298102
rect 9138 297978 9758 298046
rect 9138 297922 9234 297978
rect 9290 297922 9358 297978
rect 9414 297922 9482 297978
rect 9538 297922 9606 297978
rect 9662 297922 9758 297978
rect 9138 280350 9758 297922
rect 9138 280294 9234 280350
rect 9290 280294 9358 280350
rect 9414 280294 9482 280350
rect 9538 280294 9606 280350
rect 9662 280294 9758 280350
rect 9138 280226 9758 280294
rect 9138 280170 9234 280226
rect 9290 280170 9358 280226
rect 9414 280170 9482 280226
rect 9538 280170 9606 280226
rect 9662 280170 9758 280226
rect 9138 280102 9758 280170
rect 9138 280046 9234 280102
rect 9290 280046 9358 280102
rect 9414 280046 9482 280102
rect 9538 280046 9606 280102
rect 9662 280046 9758 280102
rect 9138 279978 9758 280046
rect 9138 279922 9234 279978
rect 9290 279922 9358 279978
rect 9414 279922 9482 279978
rect 9538 279922 9606 279978
rect 9662 279922 9758 279978
rect 9138 262350 9758 279922
rect 10892 299348 10948 299358
rect 10892 262836 10948 299292
rect 10892 262770 10948 262780
rect 9138 262294 9234 262350
rect 9290 262294 9358 262350
rect 9414 262294 9482 262350
rect 9538 262294 9606 262350
rect 9662 262294 9758 262350
rect 9138 262226 9758 262294
rect 9138 262170 9234 262226
rect 9290 262170 9358 262226
rect 9414 262170 9482 262226
rect 9538 262170 9606 262226
rect 9662 262170 9758 262226
rect 9138 262102 9758 262170
rect 9138 262046 9234 262102
rect 9290 262046 9358 262102
rect 9414 262046 9482 262102
rect 9538 262046 9606 262102
rect 9662 262046 9758 262102
rect 9138 261978 9758 262046
rect 9138 261922 9234 261978
rect 9290 261922 9358 261978
rect 9414 261922 9482 261978
rect 9538 261922 9606 261978
rect 9662 261922 9758 261978
rect 9138 244350 9758 261922
rect 9138 244294 9234 244350
rect 9290 244294 9358 244350
rect 9414 244294 9482 244350
rect 9538 244294 9606 244350
rect 9662 244294 9758 244350
rect 9138 244226 9758 244294
rect 9138 244170 9234 244226
rect 9290 244170 9358 244226
rect 9414 244170 9482 244226
rect 9538 244170 9606 244226
rect 9662 244170 9758 244226
rect 9138 244102 9758 244170
rect 9138 244046 9234 244102
rect 9290 244046 9358 244102
rect 9414 244046 9482 244102
rect 9538 244046 9606 244102
rect 9662 244046 9758 244102
rect 9138 243978 9758 244046
rect 9138 243922 9234 243978
rect 9290 243922 9358 243978
rect 9414 243922 9482 243978
rect 9538 243922 9606 243978
rect 9662 243922 9758 243978
rect 9138 226350 9758 243922
rect 9138 226294 9234 226350
rect 9290 226294 9358 226350
rect 9414 226294 9482 226350
rect 9538 226294 9606 226350
rect 9662 226294 9758 226350
rect 9138 226226 9758 226294
rect 9138 226170 9234 226226
rect 9290 226170 9358 226226
rect 9414 226170 9482 226226
rect 9538 226170 9606 226226
rect 9662 226170 9758 226226
rect 9138 226102 9758 226170
rect 9138 226046 9234 226102
rect 9290 226046 9358 226102
rect 9414 226046 9482 226102
rect 9538 226046 9606 226102
rect 9662 226046 9758 226102
rect 9138 225978 9758 226046
rect 9138 225922 9234 225978
rect 9290 225922 9358 225978
rect 9414 225922 9482 225978
rect 9538 225922 9606 225978
rect 9662 225922 9758 225978
rect 9138 208350 9758 225922
rect 12572 220276 12628 300188
rect 12572 220210 12628 220220
rect 9138 208294 9234 208350
rect 9290 208294 9358 208350
rect 9414 208294 9482 208350
rect 9538 208294 9606 208350
rect 9662 208294 9758 208350
rect 9138 208226 9758 208294
rect 9138 208170 9234 208226
rect 9290 208170 9358 208226
rect 9414 208170 9482 208226
rect 9538 208170 9606 208226
rect 9662 208170 9758 208226
rect 9138 208102 9758 208170
rect 9138 208046 9234 208102
rect 9290 208046 9358 208102
rect 9414 208046 9482 208102
rect 9538 208046 9606 208102
rect 9662 208046 9758 208102
rect 9138 207978 9758 208046
rect 9138 207922 9234 207978
rect 9290 207922 9358 207978
rect 9414 207922 9482 207978
rect 9538 207922 9606 207978
rect 9662 207922 9758 207978
rect 9138 190350 9758 207922
rect 9138 190294 9234 190350
rect 9290 190294 9358 190350
rect 9414 190294 9482 190350
rect 9538 190294 9606 190350
rect 9662 190294 9758 190350
rect 9138 190226 9758 190294
rect 9138 190170 9234 190226
rect 9290 190170 9358 190226
rect 9414 190170 9482 190226
rect 9538 190170 9606 190226
rect 9662 190170 9758 190226
rect 9138 190102 9758 190170
rect 9138 190046 9234 190102
rect 9290 190046 9358 190102
rect 9414 190046 9482 190102
rect 9538 190046 9606 190102
rect 9662 190046 9758 190102
rect 9138 189978 9758 190046
rect 9138 189922 9234 189978
rect 9290 189922 9358 189978
rect 9414 189922 9482 189978
rect 9538 189922 9606 189978
rect 9662 189922 9758 189978
rect 9138 172350 9758 189922
rect 9138 172294 9234 172350
rect 9290 172294 9358 172350
rect 9414 172294 9482 172350
rect 9538 172294 9606 172350
rect 9662 172294 9758 172350
rect 9138 172226 9758 172294
rect 9138 172170 9234 172226
rect 9290 172170 9358 172226
rect 9414 172170 9482 172226
rect 9538 172170 9606 172226
rect 9662 172170 9758 172226
rect 9138 172102 9758 172170
rect 9138 172046 9234 172102
rect 9290 172046 9358 172102
rect 9414 172046 9482 172102
rect 9538 172046 9606 172102
rect 9662 172046 9758 172102
rect 9138 171978 9758 172046
rect 9138 171922 9234 171978
rect 9290 171922 9358 171978
rect 9414 171922 9482 171978
rect 9538 171922 9606 171978
rect 9662 171922 9758 171978
rect 9138 154350 9758 171922
rect 9138 154294 9234 154350
rect 9290 154294 9358 154350
rect 9414 154294 9482 154350
rect 9538 154294 9606 154350
rect 9662 154294 9758 154350
rect 9138 154226 9758 154294
rect 9138 154170 9234 154226
rect 9290 154170 9358 154226
rect 9414 154170 9482 154226
rect 9538 154170 9606 154226
rect 9662 154170 9758 154226
rect 9138 154102 9758 154170
rect 9138 154046 9234 154102
rect 9290 154046 9358 154102
rect 9414 154046 9482 154102
rect 9538 154046 9606 154102
rect 9662 154046 9758 154102
rect 9138 153978 9758 154046
rect 9138 153922 9234 153978
rect 9290 153922 9358 153978
rect 9414 153922 9482 153978
rect 9538 153922 9606 153978
rect 9662 153922 9758 153978
rect 5418 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 6038 148350
rect 5418 148226 6038 148294
rect 5418 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 6038 148226
rect 5418 148102 6038 148170
rect 5418 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 6038 148102
rect 5418 147978 6038 148046
rect 5418 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 6038 147978
rect 5418 130350 6038 147922
rect 5418 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 6038 130350
rect 5418 130226 6038 130294
rect 5418 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 6038 130226
rect 5418 130102 6038 130170
rect 5418 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 6038 130102
rect 5418 129978 6038 130046
rect 5418 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 6038 129978
rect 5418 112350 6038 129922
rect 5418 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 6038 112350
rect 5418 112226 6038 112294
rect 5418 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 6038 112226
rect 5418 112102 6038 112170
rect 5418 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 6038 112102
rect 5418 111978 6038 112046
rect 5418 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 6038 111978
rect 5418 94350 6038 111922
rect 5418 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 6038 94350
rect 5418 94226 6038 94294
rect 5418 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 6038 94226
rect 5418 94102 6038 94170
rect 5418 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 6038 94102
rect 5418 93978 6038 94046
rect 5418 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 6038 93978
rect 5418 76350 6038 93922
rect 5418 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 6038 76350
rect 5418 76226 6038 76294
rect 5418 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 6038 76226
rect 5418 76102 6038 76170
rect 5418 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 6038 76102
rect 5418 75978 6038 76046
rect 5418 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 6038 75978
rect 5418 58350 6038 75922
rect 5418 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 6038 58350
rect 5418 58226 6038 58294
rect 5418 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 6038 58226
rect 5418 58102 6038 58170
rect 5418 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 6038 58102
rect 5418 57978 6038 58046
rect 5418 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 6038 57978
rect 4172 8754 4228 8764
rect 5418 40350 6038 57922
rect 5418 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 6038 40350
rect 5418 40226 6038 40294
rect 5418 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 6038 40226
rect 5418 40102 6038 40170
rect 5418 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 6038 40102
rect 5418 39978 6038 40046
rect 5418 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 6038 39978
rect 5418 22350 6038 39922
rect 5418 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 6038 22350
rect 5418 22226 6038 22294
rect 5418 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 6038 22226
rect 5418 22102 6038 22170
rect 5418 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 6038 22102
rect 5418 21978 6038 22046
rect 5418 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 6038 21978
rect -956 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 -336 4350
rect -956 4226 -336 4294
rect -956 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 -336 4226
rect -956 4102 -336 4170
rect -956 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 -336 4102
rect -956 3978 -336 4046
rect -956 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 -336 3978
rect -956 -160 -336 3922
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 -336 -160
rect -956 -284 -336 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 -336 -284
rect -956 -408 -336 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 -336 -408
rect -956 -532 -336 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 -336 -532
rect -956 -684 -336 -588
rect 5418 4350 6038 21922
rect 5418 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 6038 4350
rect 5418 4226 6038 4294
rect 5418 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 6038 4226
rect 5418 4102 6038 4170
rect 5418 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 6038 4102
rect 5418 3978 6038 4046
rect 5418 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 6038 3978
rect 5418 -160 6038 3922
rect 5418 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 6038 -160
rect 5418 -284 6038 -216
rect 5418 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 6038 -284
rect 5418 -408 6038 -340
rect 5418 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 6038 -408
rect 5418 -532 6038 -464
rect 5418 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 6038 -532
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 -1296 -1120
rect -1916 -1244 -1296 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 -1296 -1244
rect -1916 -1368 -1296 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 -1296 -1368
rect -1916 -1492 -1296 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 -1296 -1492
rect -1916 -1644 -1296 -1548
rect 5418 -1644 6038 -588
rect 9138 136350 9758 153922
rect 9138 136294 9234 136350
rect 9290 136294 9358 136350
rect 9414 136294 9482 136350
rect 9538 136294 9606 136350
rect 9662 136294 9758 136350
rect 9138 136226 9758 136294
rect 9138 136170 9234 136226
rect 9290 136170 9358 136226
rect 9414 136170 9482 136226
rect 9538 136170 9606 136226
rect 9662 136170 9758 136226
rect 9138 136102 9758 136170
rect 9138 136046 9234 136102
rect 9290 136046 9358 136102
rect 9414 136046 9482 136102
rect 9538 136046 9606 136102
rect 9662 136046 9758 136102
rect 9138 135978 9758 136046
rect 9138 135922 9234 135978
rect 9290 135922 9358 135978
rect 9414 135922 9482 135978
rect 9538 135922 9606 135978
rect 9662 135922 9758 135978
rect 9138 118350 9758 135922
rect 9138 118294 9234 118350
rect 9290 118294 9358 118350
rect 9414 118294 9482 118350
rect 9538 118294 9606 118350
rect 9662 118294 9758 118350
rect 9138 118226 9758 118294
rect 9138 118170 9234 118226
rect 9290 118170 9358 118226
rect 9414 118170 9482 118226
rect 9538 118170 9606 118226
rect 9662 118170 9758 118226
rect 9138 118102 9758 118170
rect 9138 118046 9234 118102
rect 9290 118046 9358 118102
rect 9414 118046 9482 118102
rect 9538 118046 9606 118102
rect 9662 118046 9758 118102
rect 9138 117978 9758 118046
rect 9138 117922 9234 117978
rect 9290 117922 9358 117978
rect 9414 117922 9482 117978
rect 9538 117922 9606 117978
rect 9662 117922 9758 117978
rect 9138 100350 9758 117922
rect 9138 100294 9234 100350
rect 9290 100294 9358 100350
rect 9414 100294 9482 100350
rect 9538 100294 9606 100350
rect 9662 100294 9758 100350
rect 9138 100226 9758 100294
rect 9138 100170 9234 100226
rect 9290 100170 9358 100226
rect 9414 100170 9482 100226
rect 9538 100170 9606 100226
rect 9662 100170 9758 100226
rect 9138 100102 9758 100170
rect 9138 100046 9234 100102
rect 9290 100046 9358 100102
rect 9414 100046 9482 100102
rect 9538 100046 9606 100102
rect 9662 100046 9758 100102
rect 9138 99978 9758 100046
rect 9138 99922 9234 99978
rect 9290 99922 9358 99978
rect 9414 99922 9482 99978
rect 9538 99922 9606 99978
rect 9662 99922 9758 99978
rect 9138 82350 9758 99922
rect 9138 82294 9234 82350
rect 9290 82294 9358 82350
rect 9414 82294 9482 82350
rect 9538 82294 9606 82350
rect 9662 82294 9758 82350
rect 9138 82226 9758 82294
rect 9138 82170 9234 82226
rect 9290 82170 9358 82226
rect 9414 82170 9482 82226
rect 9538 82170 9606 82226
rect 9662 82170 9758 82226
rect 9138 82102 9758 82170
rect 9138 82046 9234 82102
rect 9290 82046 9358 82102
rect 9414 82046 9482 82102
rect 9538 82046 9606 82102
rect 9662 82046 9758 82102
rect 9138 81978 9758 82046
rect 9138 81922 9234 81978
rect 9290 81922 9358 81978
rect 9414 81922 9482 81978
rect 9538 81922 9606 81978
rect 9662 81922 9758 81978
rect 9138 64350 9758 81922
rect 27692 65044 27748 385262
rect 36138 382350 36758 399922
rect 36138 382294 36234 382350
rect 36290 382294 36358 382350
rect 36414 382294 36482 382350
rect 36538 382294 36606 382350
rect 36662 382294 36758 382350
rect 36138 382226 36758 382294
rect 36138 382170 36234 382226
rect 36290 382170 36358 382226
rect 36414 382170 36482 382226
rect 36538 382170 36606 382226
rect 36662 382170 36758 382226
rect 36138 382102 36758 382170
rect 36138 382046 36234 382102
rect 36290 382046 36358 382102
rect 36414 382046 36482 382102
rect 36538 382046 36606 382102
rect 36662 382046 36758 382102
rect 36138 381978 36758 382046
rect 36138 381922 36234 381978
rect 36290 381922 36358 381978
rect 36414 381922 36482 381978
rect 36538 381922 36606 381978
rect 36662 381922 36758 381978
rect 36138 364350 36758 381922
rect 36138 364294 36234 364350
rect 36290 364294 36358 364350
rect 36414 364294 36482 364350
rect 36538 364294 36606 364350
rect 36662 364294 36758 364350
rect 36138 364226 36758 364294
rect 36138 364170 36234 364226
rect 36290 364170 36358 364226
rect 36414 364170 36482 364226
rect 36538 364170 36606 364226
rect 36662 364170 36758 364226
rect 36138 364102 36758 364170
rect 36138 364046 36234 364102
rect 36290 364046 36358 364102
rect 36414 364046 36482 364102
rect 36538 364046 36606 364102
rect 36662 364046 36758 364102
rect 36138 363978 36758 364046
rect 36138 363922 36234 363978
rect 36290 363922 36358 363978
rect 36414 363922 36482 363978
rect 36538 363922 36606 363978
rect 36662 363922 36758 363978
rect 36138 346350 36758 363922
rect 36138 346294 36234 346350
rect 36290 346294 36358 346350
rect 36414 346294 36482 346350
rect 36538 346294 36606 346350
rect 36662 346294 36758 346350
rect 36138 346226 36758 346294
rect 36138 346170 36234 346226
rect 36290 346170 36358 346226
rect 36414 346170 36482 346226
rect 36538 346170 36606 346226
rect 36662 346170 36758 346226
rect 36138 346102 36758 346170
rect 36138 346046 36234 346102
rect 36290 346046 36358 346102
rect 36414 346046 36482 346102
rect 36538 346046 36606 346102
rect 36662 346046 36758 346102
rect 36138 345978 36758 346046
rect 36138 345922 36234 345978
rect 36290 345922 36358 345978
rect 36414 345922 36482 345978
rect 36538 345922 36606 345978
rect 36662 345922 36758 345978
rect 36138 328350 36758 345922
rect 36138 328294 36234 328350
rect 36290 328294 36358 328350
rect 36414 328294 36482 328350
rect 36538 328294 36606 328350
rect 36662 328294 36758 328350
rect 36138 328226 36758 328294
rect 36138 328170 36234 328226
rect 36290 328170 36358 328226
rect 36414 328170 36482 328226
rect 36538 328170 36606 328226
rect 36662 328170 36758 328226
rect 36138 328102 36758 328170
rect 36138 328046 36234 328102
rect 36290 328046 36358 328102
rect 36414 328046 36482 328102
rect 36538 328046 36606 328102
rect 36662 328046 36758 328102
rect 36138 327978 36758 328046
rect 36138 327922 36234 327978
rect 36290 327922 36358 327978
rect 36414 327922 36482 327978
rect 36538 327922 36606 327978
rect 36662 327922 36758 327978
rect 36138 310350 36758 327922
rect 36138 310294 36234 310350
rect 36290 310294 36358 310350
rect 36414 310294 36482 310350
rect 36538 310294 36606 310350
rect 36662 310294 36758 310350
rect 36138 310226 36758 310294
rect 36138 310170 36234 310226
rect 36290 310170 36358 310226
rect 36414 310170 36482 310226
rect 36538 310170 36606 310226
rect 36662 310170 36758 310226
rect 36138 310102 36758 310170
rect 36138 310046 36234 310102
rect 36290 310046 36358 310102
rect 36414 310046 36482 310102
rect 36538 310046 36606 310102
rect 36662 310046 36758 310102
rect 36138 309978 36758 310046
rect 36138 309922 36234 309978
rect 36290 309922 36358 309978
rect 36414 309922 36482 309978
rect 36538 309922 36606 309978
rect 36662 309922 36758 309978
rect 29372 303604 29428 303614
rect 27804 301364 27860 301374
rect 27804 177940 27860 301308
rect 27804 177874 27860 177884
rect 29372 93268 29428 303548
rect 32732 302596 32788 302606
rect 32732 135604 32788 302540
rect 32732 135538 32788 135548
rect 36138 292350 36758 309922
rect 36138 292294 36234 292350
rect 36290 292294 36358 292350
rect 36414 292294 36482 292350
rect 36538 292294 36606 292350
rect 36662 292294 36758 292350
rect 36138 292226 36758 292294
rect 36138 292170 36234 292226
rect 36290 292170 36358 292226
rect 36414 292170 36482 292226
rect 36538 292170 36606 292226
rect 36662 292170 36758 292226
rect 36138 292102 36758 292170
rect 36138 292046 36234 292102
rect 36290 292046 36358 292102
rect 36414 292046 36482 292102
rect 36538 292046 36606 292102
rect 36662 292046 36758 292102
rect 36138 291978 36758 292046
rect 36138 291922 36234 291978
rect 36290 291922 36358 291978
rect 36414 291922 36482 291978
rect 36538 291922 36606 291978
rect 36662 291922 36758 291978
rect 36138 274350 36758 291922
rect 36138 274294 36234 274350
rect 36290 274294 36358 274350
rect 36414 274294 36482 274350
rect 36538 274294 36606 274350
rect 36662 274294 36758 274350
rect 36138 274226 36758 274294
rect 36138 274170 36234 274226
rect 36290 274170 36358 274226
rect 36414 274170 36482 274226
rect 36538 274170 36606 274226
rect 36662 274170 36758 274226
rect 36138 274102 36758 274170
rect 36138 274046 36234 274102
rect 36290 274046 36358 274102
rect 36414 274046 36482 274102
rect 36538 274046 36606 274102
rect 36662 274046 36758 274102
rect 36138 273978 36758 274046
rect 36138 273922 36234 273978
rect 36290 273922 36358 273978
rect 36414 273922 36482 273978
rect 36538 273922 36606 273978
rect 36662 273922 36758 273978
rect 36138 256350 36758 273922
rect 36138 256294 36234 256350
rect 36290 256294 36358 256350
rect 36414 256294 36482 256350
rect 36538 256294 36606 256350
rect 36662 256294 36758 256350
rect 36138 256226 36758 256294
rect 36138 256170 36234 256226
rect 36290 256170 36358 256226
rect 36414 256170 36482 256226
rect 36538 256170 36606 256226
rect 36662 256170 36758 256226
rect 36138 256102 36758 256170
rect 36138 256046 36234 256102
rect 36290 256046 36358 256102
rect 36414 256046 36482 256102
rect 36538 256046 36606 256102
rect 36662 256046 36758 256102
rect 36138 255978 36758 256046
rect 36138 255922 36234 255978
rect 36290 255922 36358 255978
rect 36414 255922 36482 255978
rect 36538 255922 36606 255978
rect 36662 255922 36758 255978
rect 36138 238350 36758 255922
rect 36138 238294 36234 238350
rect 36290 238294 36358 238350
rect 36414 238294 36482 238350
rect 36538 238294 36606 238350
rect 36662 238294 36758 238350
rect 36138 238226 36758 238294
rect 36138 238170 36234 238226
rect 36290 238170 36358 238226
rect 36414 238170 36482 238226
rect 36538 238170 36606 238226
rect 36662 238170 36758 238226
rect 36138 238102 36758 238170
rect 36138 238046 36234 238102
rect 36290 238046 36358 238102
rect 36414 238046 36482 238102
rect 36538 238046 36606 238102
rect 36662 238046 36758 238102
rect 36138 237978 36758 238046
rect 36138 237922 36234 237978
rect 36290 237922 36358 237978
rect 36414 237922 36482 237978
rect 36538 237922 36606 237978
rect 36662 237922 36758 237978
rect 36138 220350 36758 237922
rect 36138 220294 36234 220350
rect 36290 220294 36358 220350
rect 36414 220294 36482 220350
rect 36538 220294 36606 220350
rect 36662 220294 36758 220350
rect 36138 220226 36758 220294
rect 36138 220170 36234 220226
rect 36290 220170 36358 220226
rect 36414 220170 36482 220226
rect 36538 220170 36606 220226
rect 36662 220170 36758 220226
rect 36138 220102 36758 220170
rect 36138 220046 36234 220102
rect 36290 220046 36358 220102
rect 36414 220046 36482 220102
rect 36538 220046 36606 220102
rect 36662 220046 36758 220102
rect 36138 219978 36758 220046
rect 36138 219922 36234 219978
rect 36290 219922 36358 219978
rect 36414 219922 36482 219978
rect 36538 219922 36606 219978
rect 36662 219922 36758 219978
rect 36138 202350 36758 219922
rect 36138 202294 36234 202350
rect 36290 202294 36358 202350
rect 36414 202294 36482 202350
rect 36538 202294 36606 202350
rect 36662 202294 36758 202350
rect 36138 202226 36758 202294
rect 36138 202170 36234 202226
rect 36290 202170 36358 202226
rect 36414 202170 36482 202226
rect 36538 202170 36606 202226
rect 36662 202170 36758 202226
rect 36138 202102 36758 202170
rect 36138 202046 36234 202102
rect 36290 202046 36358 202102
rect 36414 202046 36482 202102
rect 36538 202046 36606 202102
rect 36662 202046 36758 202102
rect 36138 201978 36758 202046
rect 36138 201922 36234 201978
rect 36290 201922 36358 201978
rect 36414 201922 36482 201978
rect 36538 201922 36606 201978
rect 36662 201922 36758 201978
rect 36138 184350 36758 201922
rect 36138 184294 36234 184350
rect 36290 184294 36358 184350
rect 36414 184294 36482 184350
rect 36538 184294 36606 184350
rect 36662 184294 36758 184350
rect 36138 184226 36758 184294
rect 36138 184170 36234 184226
rect 36290 184170 36358 184226
rect 36414 184170 36482 184226
rect 36538 184170 36606 184226
rect 36662 184170 36758 184226
rect 36138 184102 36758 184170
rect 36138 184046 36234 184102
rect 36290 184046 36358 184102
rect 36414 184046 36482 184102
rect 36538 184046 36606 184102
rect 36662 184046 36758 184102
rect 36138 183978 36758 184046
rect 36138 183922 36234 183978
rect 36290 183922 36358 183978
rect 36414 183922 36482 183978
rect 36538 183922 36606 183978
rect 36662 183922 36758 183978
rect 36138 166350 36758 183922
rect 36138 166294 36234 166350
rect 36290 166294 36358 166350
rect 36414 166294 36482 166350
rect 36538 166294 36606 166350
rect 36662 166294 36758 166350
rect 36138 166226 36758 166294
rect 36138 166170 36234 166226
rect 36290 166170 36358 166226
rect 36414 166170 36482 166226
rect 36538 166170 36606 166226
rect 36662 166170 36758 166226
rect 36138 166102 36758 166170
rect 36138 166046 36234 166102
rect 36290 166046 36358 166102
rect 36414 166046 36482 166102
rect 36538 166046 36606 166102
rect 36662 166046 36758 166102
rect 36138 165978 36758 166046
rect 36138 165922 36234 165978
rect 36290 165922 36358 165978
rect 36414 165922 36482 165978
rect 36538 165922 36606 165978
rect 36662 165922 36758 165978
rect 36138 148350 36758 165922
rect 36138 148294 36234 148350
rect 36290 148294 36358 148350
rect 36414 148294 36482 148350
rect 36538 148294 36606 148350
rect 36662 148294 36758 148350
rect 36138 148226 36758 148294
rect 36138 148170 36234 148226
rect 36290 148170 36358 148226
rect 36414 148170 36482 148226
rect 36538 148170 36606 148226
rect 36662 148170 36758 148226
rect 36138 148102 36758 148170
rect 36138 148046 36234 148102
rect 36290 148046 36358 148102
rect 36414 148046 36482 148102
rect 36538 148046 36606 148102
rect 36662 148046 36758 148102
rect 36138 147978 36758 148046
rect 36138 147922 36234 147978
rect 36290 147922 36358 147978
rect 36414 147922 36482 147978
rect 36538 147922 36606 147978
rect 36662 147922 36758 147978
rect 29372 93202 29428 93212
rect 36138 130350 36758 147922
rect 36138 130294 36234 130350
rect 36290 130294 36358 130350
rect 36414 130294 36482 130350
rect 36538 130294 36606 130350
rect 36662 130294 36758 130350
rect 36138 130226 36758 130294
rect 36138 130170 36234 130226
rect 36290 130170 36358 130226
rect 36414 130170 36482 130226
rect 36538 130170 36606 130226
rect 36662 130170 36758 130226
rect 36138 130102 36758 130170
rect 36138 130046 36234 130102
rect 36290 130046 36358 130102
rect 36414 130046 36482 130102
rect 36538 130046 36606 130102
rect 36662 130046 36758 130102
rect 36138 129978 36758 130046
rect 36138 129922 36234 129978
rect 36290 129922 36358 129978
rect 36414 129922 36482 129978
rect 36538 129922 36606 129978
rect 36662 129922 36758 129978
rect 36138 112350 36758 129922
rect 36138 112294 36234 112350
rect 36290 112294 36358 112350
rect 36414 112294 36482 112350
rect 36538 112294 36606 112350
rect 36662 112294 36758 112350
rect 36138 112226 36758 112294
rect 36138 112170 36234 112226
rect 36290 112170 36358 112226
rect 36414 112170 36482 112226
rect 36538 112170 36606 112226
rect 36662 112170 36758 112226
rect 36138 112102 36758 112170
rect 36138 112046 36234 112102
rect 36290 112046 36358 112102
rect 36414 112046 36482 112102
rect 36538 112046 36606 112102
rect 36662 112046 36758 112102
rect 36138 111978 36758 112046
rect 36138 111922 36234 111978
rect 36290 111922 36358 111978
rect 36414 111922 36482 111978
rect 36538 111922 36606 111978
rect 36662 111922 36758 111978
rect 36138 94350 36758 111922
rect 36138 94294 36234 94350
rect 36290 94294 36358 94350
rect 36414 94294 36482 94350
rect 36538 94294 36606 94350
rect 36662 94294 36758 94350
rect 36138 94226 36758 94294
rect 36138 94170 36234 94226
rect 36290 94170 36358 94226
rect 36414 94170 36482 94226
rect 36538 94170 36606 94226
rect 36662 94170 36758 94226
rect 36138 94102 36758 94170
rect 36138 94046 36234 94102
rect 36290 94046 36358 94102
rect 36414 94046 36482 94102
rect 36538 94046 36606 94102
rect 36662 94046 36758 94102
rect 36138 93978 36758 94046
rect 36138 93922 36234 93978
rect 36290 93922 36358 93978
rect 36414 93922 36482 93978
rect 36538 93922 36606 93978
rect 36662 93922 36758 93978
rect 27692 64978 27748 64988
rect 36138 76350 36758 93922
rect 36138 76294 36234 76350
rect 36290 76294 36358 76350
rect 36414 76294 36482 76350
rect 36538 76294 36606 76350
rect 36662 76294 36758 76350
rect 36138 76226 36758 76294
rect 36138 76170 36234 76226
rect 36290 76170 36358 76226
rect 36414 76170 36482 76226
rect 36538 76170 36606 76226
rect 36662 76170 36758 76226
rect 36138 76102 36758 76170
rect 36138 76046 36234 76102
rect 36290 76046 36358 76102
rect 36414 76046 36482 76102
rect 36538 76046 36606 76102
rect 36662 76046 36758 76102
rect 36138 75978 36758 76046
rect 36138 75922 36234 75978
rect 36290 75922 36358 75978
rect 36414 75922 36482 75978
rect 36538 75922 36606 75978
rect 36662 75922 36758 75978
rect 9138 64294 9234 64350
rect 9290 64294 9358 64350
rect 9414 64294 9482 64350
rect 9538 64294 9606 64350
rect 9662 64294 9758 64350
rect 9138 64226 9758 64294
rect 9138 64170 9234 64226
rect 9290 64170 9358 64226
rect 9414 64170 9482 64226
rect 9538 64170 9606 64226
rect 9662 64170 9758 64226
rect 9138 64102 9758 64170
rect 9138 64046 9234 64102
rect 9290 64046 9358 64102
rect 9414 64046 9482 64102
rect 9538 64046 9606 64102
rect 9662 64046 9758 64102
rect 9138 63978 9758 64046
rect 9138 63922 9234 63978
rect 9290 63922 9358 63978
rect 9414 63922 9482 63978
rect 9538 63922 9606 63978
rect 9662 63922 9758 63978
rect 9138 46350 9758 63922
rect 9138 46294 9234 46350
rect 9290 46294 9358 46350
rect 9414 46294 9482 46350
rect 9538 46294 9606 46350
rect 9662 46294 9758 46350
rect 9138 46226 9758 46294
rect 9138 46170 9234 46226
rect 9290 46170 9358 46226
rect 9414 46170 9482 46226
rect 9538 46170 9606 46226
rect 9662 46170 9758 46226
rect 9138 46102 9758 46170
rect 9138 46046 9234 46102
rect 9290 46046 9358 46102
rect 9414 46046 9482 46102
rect 9538 46046 9606 46102
rect 9662 46046 9758 46102
rect 9138 45978 9758 46046
rect 9138 45922 9234 45978
rect 9290 45922 9358 45978
rect 9414 45922 9482 45978
rect 9538 45922 9606 45978
rect 9662 45922 9758 45978
rect 9138 28350 9758 45922
rect 9138 28294 9234 28350
rect 9290 28294 9358 28350
rect 9414 28294 9482 28350
rect 9538 28294 9606 28350
rect 9662 28294 9758 28350
rect 9138 28226 9758 28294
rect 9138 28170 9234 28226
rect 9290 28170 9358 28226
rect 9414 28170 9482 28226
rect 9538 28170 9606 28226
rect 9662 28170 9758 28226
rect 9138 28102 9758 28170
rect 9138 28046 9234 28102
rect 9290 28046 9358 28102
rect 9414 28046 9482 28102
rect 9538 28046 9606 28102
rect 9662 28046 9758 28102
rect 9138 27978 9758 28046
rect 9138 27922 9234 27978
rect 9290 27922 9358 27978
rect 9414 27922 9482 27978
rect 9538 27922 9606 27978
rect 9662 27922 9758 27978
rect 9138 10350 9758 27922
rect 9138 10294 9234 10350
rect 9290 10294 9358 10350
rect 9414 10294 9482 10350
rect 9538 10294 9606 10350
rect 9662 10294 9758 10350
rect 9138 10226 9758 10294
rect 9138 10170 9234 10226
rect 9290 10170 9358 10226
rect 9414 10170 9482 10226
rect 9538 10170 9606 10226
rect 9662 10170 9758 10226
rect 9138 10102 9758 10170
rect 9138 10046 9234 10102
rect 9290 10046 9358 10102
rect 9414 10046 9482 10102
rect 9538 10046 9606 10102
rect 9662 10046 9758 10102
rect 9138 9978 9758 10046
rect 9138 9922 9234 9978
rect 9290 9922 9358 9978
rect 9414 9922 9482 9978
rect 9538 9922 9606 9978
rect 9662 9922 9758 9978
rect 9138 -1120 9758 9922
rect 9138 -1176 9234 -1120
rect 9290 -1176 9358 -1120
rect 9414 -1176 9482 -1120
rect 9538 -1176 9606 -1120
rect 9662 -1176 9758 -1120
rect 9138 -1244 9758 -1176
rect 9138 -1300 9234 -1244
rect 9290 -1300 9358 -1244
rect 9414 -1300 9482 -1244
rect 9538 -1300 9606 -1244
rect 9662 -1300 9758 -1244
rect 9138 -1368 9758 -1300
rect 9138 -1424 9234 -1368
rect 9290 -1424 9358 -1368
rect 9414 -1424 9482 -1368
rect 9538 -1424 9606 -1368
rect 9662 -1424 9758 -1368
rect 9138 -1492 9758 -1424
rect 9138 -1548 9234 -1492
rect 9290 -1548 9358 -1492
rect 9414 -1548 9482 -1492
rect 9538 -1548 9606 -1492
rect 9662 -1548 9758 -1492
rect 9138 -1644 9758 -1548
rect 36138 58350 36758 75922
rect 36138 58294 36234 58350
rect 36290 58294 36358 58350
rect 36414 58294 36482 58350
rect 36538 58294 36606 58350
rect 36662 58294 36758 58350
rect 36138 58226 36758 58294
rect 36138 58170 36234 58226
rect 36290 58170 36358 58226
rect 36414 58170 36482 58226
rect 36538 58170 36606 58226
rect 36662 58170 36758 58226
rect 36138 58102 36758 58170
rect 36138 58046 36234 58102
rect 36290 58046 36358 58102
rect 36414 58046 36482 58102
rect 36538 58046 36606 58102
rect 36662 58046 36758 58102
rect 36138 57978 36758 58046
rect 36138 57922 36234 57978
rect 36290 57922 36358 57978
rect 36414 57922 36482 57978
rect 36538 57922 36606 57978
rect 36662 57922 36758 57978
rect 36138 40350 36758 57922
rect 36138 40294 36234 40350
rect 36290 40294 36358 40350
rect 36414 40294 36482 40350
rect 36538 40294 36606 40350
rect 36662 40294 36758 40350
rect 36138 40226 36758 40294
rect 36138 40170 36234 40226
rect 36290 40170 36358 40226
rect 36414 40170 36482 40226
rect 36538 40170 36606 40226
rect 36662 40170 36758 40226
rect 36138 40102 36758 40170
rect 36138 40046 36234 40102
rect 36290 40046 36358 40102
rect 36414 40046 36482 40102
rect 36538 40046 36606 40102
rect 36662 40046 36758 40102
rect 36138 39978 36758 40046
rect 36138 39922 36234 39978
rect 36290 39922 36358 39978
rect 36414 39922 36482 39978
rect 36538 39922 36606 39978
rect 36662 39922 36758 39978
rect 36138 22350 36758 39922
rect 36138 22294 36234 22350
rect 36290 22294 36358 22350
rect 36414 22294 36482 22350
rect 36538 22294 36606 22350
rect 36662 22294 36758 22350
rect 36138 22226 36758 22294
rect 36138 22170 36234 22226
rect 36290 22170 36358 22226
rect 36414 22170 36482 22226
rect 36538 22170 36606 22226
rect 36662 22170 36758 22226
rect 36138 22102 36758 22170
rect 36138 22046 36234 22102
rect 36290 22046 36358 22102
rect 36414 22046 36482 22102
rect 36538 22046 36606 22102
rect 36662 22046 36758 22102
rect 36138 21978 36758 22046
rect 36138 21922 36234 21978
rect 36290 21922 36358 21978
rect 36414 21922 36482 21978
rect 36538 21922 36606 21978
rect 36662 21922 36758 21978
rect 36138 4350 36758 21922
rect 36138 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 36758 4350
rect 36138 4226 36758 4294
rect 36138 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 36758 4226
rect 36138 4102 36758 4170
rect 36138 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 36758 4102
rect 36138 3978 36758 4046
rect 36138 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 36758 3978
rect 36138 -160 36758 3922
rect 36138 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 36758 -160
rect 36138 -284 36758 -216
rect 36138 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 36758 -284
rect 36138 -408 36758 -340
rect 36138 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 36758 -408
rect 36138 -532 36758 -464
rect 36138 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 36758 -532
rect 36138 -1644 36758 -588
rect 39858 598172 40478 598268
rect 39858 598116 39954 598172
rect 40010 598116 40078 598172
rect 40134 598116 40202 598172
rect 40258 598116 40326 598172
rect 40382 598116 40478 598172
rect 39858 598048 40478 598116
rect 39858 597992 39954 598048
rect 40010 597992 40078 598048
rect 40134 597992 40202 598048
rect 40258 597992 40326 598048
rect 40382 597992 40478 598048
rect 39858 597924 40478 597992
rect 39858 597868 39954 597924
rect 40010 597868 40078 597924
rect 40134 597868 40202 597924
rect 40258 597868 40326 597924
rect 40382 597868 40478 597924
rect 39858 597800 40478 597868
rect 39858 597744 39954 597800
rect 40010 597744 40078 597800
rect 40134 597744 40202 597800
rect 40258 597744 40326 597800
rect 40382 597744 40478 597800
rect 39858 586350 40478 597744
rect 39858 586294 39954 586350
rect 40010 586294 40078 586350
rect 40134 586294 40202 586350
rect 40258 586294 40326 586350
rect 40382 586294 40478 586350
rect 39858 586226 40478 586294
rect 39858 586170 39954 586226
rect 40010 586170 40078 586226
rect 40134 586170 40202 586226
rect 40258 586170 40326 586226
rect 40382 586170 40478 586226
rect 39858 586102 40478 586170
rect 39858 586046 39954 586102
rect 40010 586046 40078 586102
rect 40134 586046 40202 586102
rect 40258 586046 40326 586102
rect 40382 586046 40478 586102
rect 39858 585978 40478 586046
rect 39858 585922 39954 585978
rect 40010 585922 40078 585978
rect 40134 585922 40202 585978
rect 40258 585922 40326 585978
rect 40382 585922 40478 585978
rect 39858 568350 40478 585922
rect 39858 568294 39954 568350
rect 40010 568294 40078 568350
rect 40134 568294 40202 568350
rect 40258 568294 40326 568350
rect 40382 568294 40478 568350
rect 39858 568226 40478 568294
rect 39858 568170 39954 568226
rect 40010 568170 40078 568226
rect 40134 568170 40202 568226
rect 40258 568170 40326 568226
rect 40382 568170 40478 568226
rect 39858 568102 40478 568170
rect 39858 568046 39954 568102
rect 40010 568046 40078 568102
rect 40134 568046 40202 568102
rect 40258 568046 40326 568102
rect 40382 568046 40478 568102
rect 39858 567978 40478 568046
rect 39858 567922 39954 567978
rect 40010 567922 40078 567978
rect 40134 567922 40202 567978
rect 40258 567922 40326 567978
rect 40382 567922 40478 567978
rect 39858 550350 40478 567922
rect 39858 550294 39954 550350
rect 40010 550294 40078 550350
rect 40134 550294 40202 550350
rect 40258 550294 40326 550350
rect 40382 550294 40478 550350
rect 39858 550226 40478 550294
rect 39858 550170 39954 550226
rect 40010 550170 40078 550226
rect 40134 550170 40202 550226
rect 40258 550170 40326 550226
rect 40382 550170 40478 550226
rect 39858 550102 40478 550170
rect 39858 550046 39954 550102
rect 40010 550046 40078 550102
rect 40134 550046 40202 550102
rect 40258 550046 40326 550102
rect 40382 550046 40478 550102
rect 39858 549978 40478 550046
rect 39858 549922 39954 549978
rect 40010 549922 40078 549978
rect 40134 549922 40202 549978
rect 40258 549922 40326 549978
rect 40382 549922 40478 549978
rect 39858 532350 40478 549922
rect 66858 597212 67478 598268
rect 66858 597156 66954 597212
rect 67010 597156 67078 597212
rect 67134 597156 67202 597212
rect 67258 597156 67326 597212
rect 67382 597156 67478 597212
rect 66858 597088 67478 597156
rect 66858 597032 66954 597088
rect 67010 597032 67078 597088
rect 67134 597032 67202 597088
rect 67258 597032 67326 597088
rect 67382 597032 67478 597088
rect 66858 596964 67478 597032
rect 66858 596908 66954 596964
rect 67010 596908 67078 596964
rect 67134 596908 67202 596964
rect 67258 596908 67326 596964
rect 67382 596908 67478 596964
rect 66858 596840 67478 596908
rect 66858 596784 66954 596840
rect 67010 596784 67078 596840
rect 67134 596784 67202 596840
rect 67258 596784 67326 596840
rect 67382 596784 67478 596840
rect 66858 580350 67478 596784
rect 66858 580294 66954 580350
rect 67010 580294 67078 580350
rect 67134 580294 67202 580350
rect 67258 580294 67326 580350
rect 67382 580294 67478 580350
rect 66858 580226 67478 580294
rect 66858 580170 66954 580226
rect 67010 580170 67078 580226
rect 67134 580170 67202 580226
rect 67258 580170 67326 580226
rect 67382 580170 67478 580226
rect 66858 580102 67478 580170
rect 66858 580046 66954 580102
rect 67010 580046 67078 580102
rect 67134 580046 67202 580102
rect 67258 580046 67326 580102
rect 67382 580046 67478 580102
rect 66858 579978 67478 580046
rect 66858 579922 66954 579978
rect 67010 579922 67078 579978
rect 67134 579922 67202 579978
rect 67258 579922 67326 579978
rect 67382 579922 67478 579978
rect 66858 562350 67478 579922
rect 66858 562294 66954 562350
rect 67010 562294 67078 562350
rect 67134 562294 67202 562350
rect 67258 562294 67326 562350
rect 67382 562294 67478 562350
rect 66858 562226 67478 562294
rect 66858 562170 66954 562226
rect 67010 562170 67078 562226
rect 67134 562170 67202 562226
rect 67258 562170 67326 562226
rect 67382 562170 67478 562226
rect 66858 562102 67478 562170
rect 66858 562046 66954 562102
rect 67010 562046 67078 562102
rect 67134 562046 67202 562102
rect 67258 562046 67326 562102
rect 67382 562046 67478 562102
rect 66858 561978 67478 562046
rect 66858 561922 66954 561978
rect 67010 561922 67078 561978
rect 67134 561922 67202 561978
rect 67258 561922 67326 561978
rect 67382 561922 67478 561978
rect 66858 544350 67478 561922
rect 66858 544294 66954 544350
rect 67010 544294 67078 544350
rect 67134 544294 67202 544350
rect 67258 544294 67326 544350
rect 67382 544294 67478 544350
rect 66858 544226 67478 544294
rect 66858 544170 66954 544226
rect 67010 544170 67078 544226
rect 67134 544170 67202 544226
rect 67258 544170 67326 544226
rect 67382 544170 67478 544226
rect 66858 544102 67478 544170
rect 66858 544046 66954 544102
rect 67010 544046 67078 544102
rect 67134 544046 67202 544102
rect 67258 544046 67326 544102
rect 67382 544046 67478 544102
rect 66858 543978 67478 544046
rect 66858 543922 66954 543978
rect 67010 543922 67078 543978
rect 67134 543922 67202 543978
rect 67258 543922 67326 543978
rect 67382 543922 67478 543978
rect 66858 532362 67478 543922
rect 70578 598172 71198 598268
rect 70578 598116 70674 598172
rect 70730 598116 70798 598172
rect 70854 598116 70922 598172
rect 70978 598116 71046 598172
rect 71102 598116 71198 598172
rect 70578 598048 71198 598116
rect 70578 597992 70674 598048
rect 70730 597992 70798 598048
rect 70854 597992 70922 598048
rect 70978 597992 71046 598048
rect 71102 597992 71198 598048
rect 70578 597924 71198 597992
rect 70578 597868 70674 597924
rect 70730 597868 70798 597924
rect 70854 597868 70922 597924
rect 70978 597868 71046 597924
rect 71102 597868 71198 597924
rect 70578 597800 71198 597868
rect 70578 597744 70674 597800
rect 70730 597744 70798 597800
rect 70854 597744 70922 597800
rect 70978 597744 71046 597800
rect 71102 597744 71198 597800
rect 70578 586350 71198 597744
rect 70578 586294 70674 586350
rect 70730 586294 70798 586350
rect 70854 586294 70922 586350
rect 70978 586294 71046 586350
rect 71102 586294 71198 586350
rect 70578 586226 71198 586294
rect 70578 586170 70674 586226
rect 70730 586170 70798 586226
rect 70854 586170 70922 586226
rect 70978 586170 71046 586226
rect 71102 586170 71198 586226
rect 70578 586102 71198 586170
rect 70578 586046 70674 586102
rect 70730 586046 70798 586102
rect 70854 586046 70922 586102
rect 70978 586046 71046 586102
rect 71102 586046 71198 586102
rect 70578 585978 71198 586046
rect 70578 585922 70674 585978
rect 70730 585922 70798 585978
rect 70854 585922 70922 585978
rect 70978 585922 71046 585978
rect 71102 585922 71198 585978
rect 70578 568350 71198 585922
rect 70578 568294 70674 568350
rect 70730 568294 70798 568350
rect 70854 568294 70922 568350
rect 70978 568294 71046 568350
rect 71102 568294 71198 568350
rect 70578 568226 71198 568294
rect 70578 568170 70674 568226
rect 70730 568170 70798 568226
rect 70854 568170 70922 568226
rect 70978 568170 71046 568226
rect 71102 568170 71198 568226
rect 70578 568102 71198 568170
rect 70578 568046 70674 568102
rect 70730 568046 70798 568102
rect 70854 568046 70922 568102
rect 70978 568046 71046 568102
rect 71102 568046 71198 568102
rect 70578 567978 71198 568046
rect 70578 567922 70674 567978
rect 70730 567922 70798 567978
rect 70854 567922 70922 567978
rect 70978 567922 71046 567978
rect 71102 567922 71198 567978
rect 70578 550350 71198 567922
rect 70578 550294 70674 550350
rect 70730 550294 70798 550350
rect 70854 550294 70922 550350
rect 70978 550294 71046 550350
rect 71102 550294 71198 550350
rect 70578 550226 71198 550294
rect 70578 550170 70674 550226
rect 70730 550170 70798 550226
rect 70854 550170 70922 550226
rect 70978 550170 71046 550226
rect 71102 550170 71198 550226
rect 70578 550102 71198 550170
rect 70578 550046 70674 550102
rect 70730 550046 70798 550102
rect 70854 550046 70922 550102
rect 70978 550046 71046 550102
rect 71102 550046 71198 550102
rect 70578 549978 71198 550046
rect 70578 549922 70674 549978
rect 70730 549922 70798 549978
rect 70854 549922 70922 549978
rect 70978 549922 71046 549978
rect 71102 549922 71198 549978
rect 70578 535962 71198 549922
rect 97578 597212 98198 598268
rect 97578 597156 97674 597212
rect 97730 597156 97798 597212
rect 97854 597156 97922 597212
rect 97978 597156 98046 597212
rect 98102 597156 98198 597212
rect 97578 597088 98198 597156
rect 97578 597032 97674 597088
rect 97730 597032 97798 597088
rect 97854 597032 97922 597088
rect 97978 597032 98046 597088
rect 98102 597032 98198 597088
rect 97578 596964 98198 597032
rect 97578 596908 97674 596964
rect 97730 596908 97798 596964
rect 97854 596908 97922 596964
rect 97978 596908 98046 596964
rect 98102 596908 98198 596964
rect 97578 596840 98198 596908
rect 97578 596784 97674 596840
rect 97730 596784 97798 596840
rect 97854 596784 97922 596840
rect 97978 596784 98046 596840
rect 98102 596784 98198 596840
rect 97578 580350 98198 596784
rect 97578 580294 97674 580350
rect 97730 580294 97798 580350
rect 97854 580294 97922 580350
rect 97978 580294 98046 580350
rect 98102 580294 98198 580350
rect 97578 580226 98198 580294
rect 97578 580170 97674 580226
rect 97730 580170 97798 580226
rect 97854 580170 97922 580226
rect 97978 580170 98046 580226
rect 98102 580170 98198 580226
rect 97578 580102 98198 580170
rect 97578 580046 97674 580102
rect 97730 580046 97798 580102
rect 97854 580046 97922 580102
rect 97978 580046 98046 580102
rect 98102 580046 98198 580102
rect 97578 579978 98198 580046
rect 97578 579922 97674 579978
rect 97730 579922 97798 579978
rect 97854 579922 97922 579978
rect 97978 579922 98046 579978
rect 98102 579922 98198 579978
rect 97578 562350 98198 579922
rect 97578 562294 97674 562350
rect 97730 562294 97798 562350
rect 97854 562294 97922 562350
rect 97978 562294 98046 562350
rect 98102 562294 98198 562350
rect 97578 562226 98198 562294
rect 97578 562170 97674 562226
rect 97730 562170 97798 562226
rect 97854 562170 97922 562226
rect 97978 562170 98046 562226
rect 98102 562170 98198 562226
rect 97578 562102 98198 562170
rect 97578 562046 97674 562102
rect 97730 562046 97798 562102
rect 97854 562046 97922 562102
rect 97978 562046 98046 562102
rect 98102 562046 98198 562102
rect 97578 561978 98198 562046
rect 97578 561922 97674 561978
rect 97730 561922 97798 561978
rect 97854 561922 97922 561978
rect 97978 561922 98046 561978
rect 98102 561922 98198 561978
rect 97578 544350 98198 561922
rect 101298 598172 101918 598268
rect 101298 598116 101394 598172
rect 101450 598116 101518 598172
rect 101574 598116 101642 598172
rect 101698 598116 101766 598172
rect 101822 598116 101918 598172
rect 101298 598048 101918 598116
rect 101298 597992 101394 598048
rect 101450 597992 101518 598048
rect 101574 597992 101642 598048
rect 101698 597992 101766 598048
rect 101822 597992 101918 598048
rect 101298 597924 101918 597992
rect 101298 597868 101394 597924
rect 101450 597868 101518 597924
rect 101574 597868 101642 597924
rect 101698 597868 101766 597924
rect 101822 597868 101918 597924
rect 101298 597800 101918 597868
rect 101298 597744 101394 597800
rect 101450 597744 101518 597800
rect 101574 597744 101642 597800
rect 101698 597744 101766 597800
rect 101822 597744 101918 597800
rect 101298 586350 101918 597744
rect 101298 586294 101394 586350
rect 101450 586294 101518 586350
rect 101574 586294 101642 586350
rect 101698 586294 101766 586350
rect 101822 586294 101918 586350
rect 101298 586226 101918 586294
rect 101298 586170 101394 586226
rect 101450 586170 101518 586226
rect 101574 586170 101642 586226
rect 101698 586170 101766 586226
rect 101822 586170 101918 586226
rect 101298 586102 101918 586170
rect 101298 586046 101394 586102
rect 101450 586046 101518 586102
rect 101574 586046 101642 586102
rect 101698 586046 101766 586102
rect 101822 586046 101918 586102
rect 101298 585978 101918 586046
rect 101298 585922 101394 585978
rect 101450 585922 101518 585978
rect 101574 585922 101642 585978
rect 101698 585922 101766 585978
rect 101822 585922 101918 585978
rect 101298 568350 101918 585922
rect 101298 568294 101394 568350
rect 101450 568294 101518 568350
rect 101574 568294 101642 568350
rect 101698 568294 101766 568350
rect 101822 568294 101918 568350
rect 101298 568226 101918 568294
rect 101298 568170 101394 568226
rect 101450 568170 101518 568226
rect 101574 568170 101642 568226
rect 101698 568170 101766 568226
rect 101822 568170 101918 568226
rect 101298 568102 101918 568170
rect 101298 568046 101394 568102
rect 101450 568046 101518 568102
rect 101574 568046 101642 568102
rect 101698 568046 101766 568102
rect 101822 568046 101918 568102
rect 101298 567978 101918 568046
rect 101298 567922 101394 567978
rect 101450 567922 101518 567978
rect 101574 567922 101642 567978
rect 101698 567922 101766 567978
rect 101822 567922 101918 567978
rect 101298 550350 101918 567922
rect 128298 597212 128918 598268
rect 128298 597156 128394 597212
rect 128450 597156 128518 597212
rect 128574 597156 128642 597212
rect 128698 597156 128766 597212
rect 128822 597156 128918 597212
rect 128298 597088 128918 597156
rect 128298 597032 128394 597088
rect 128450 597032 128518 597088
rect 128574 597032 128642 597088
rect 128698 597032 128766 597088
rect 128822 597032 128918 597088
rect 128298 596964 128918 597032
rect 128298 596908 128394 596964
rect 128450 596908 128518 596964
rect 128574 596908 128642 596964
rect 128698 596908 128766 596964
rect 128822 596908 128918 596964
rect 128298 596840 128918 596908
rect 128298 596784 128394 596840
rect 128450 596784 128518 596840
rect 128574 596784 128642 596840
rect 128698 596784 128766 596840
rect 128822 596784 128918 596840
rect 128298 580350 128918 596784
rect 128298 580294 128394 580350
rect 128450 580294 128518 580350
rect 128574 580294 128642 580350
rect 128698 580294 128766 580350
rect 128822 580294 128918 580350
rect 128298 580226 128918 580294
rect 128298 580170 128394 580226
rect 128450 580170 128518 580226
rect 128574 580170 128642 580226
rect 128698 580170 128766 580226
rect 128822 580170 128918 580226
rect 128298 580102 128918 580170
rect 128298 580046 128394 580102
rect 128450 580046 128518 580102
rect 128574 580046 128642 580102
rect 128698 580046 128766 580102
rect 128822 580046 128918 580102
rect 128298 579978 128918 580046
rect 128298 579922 128394 579978
rect 128450 579922 128518 579978
rect 128574 579922 128642 579978
rect 128698 579922 128766 579978
rect 128822 579922 128918 579978
rect 128298 562350 128918 579922
rect 128298 562294 128394 562350
rect 128450 562294 128518 562350
rect 128574 562294 128642 562350
rect 128698 562294 128766 562350
rect 128822 562294 128918 562350
rect 128298 562226 128918 562294
rect 128298 562170 128394 562226
rect 128450 562170 128518 562226
rect 128574 562170 128642 562226
rect 128698 562170 128766 562226
rect 128822 562170 128918 562226
rect 128298 562102 128918 562170
rect 114000 562003 120450 562050
rect 114000 561947 114035 562003
rect 114091 561947 114159 562003
rect 114215 561947 114283 562003
rect 114339 561947 114407 562003
rect 114463 561947 114531 562003
rect 114587 561947 114655 562003
rect 114711 561947 114779 562003
rect 114835 561947 114903 562003
rect 114959 561947 115027 562003
rect 115083 561947 115151 562003
rect 115207 561947 115275 562003
rect 115331 561947 115399 562003
rect 115455 561947 115523 562003
rect 115579 561947 115647 562003
rect 115703 561947 115771 562003
rect 115827 561947 115895 562003
rect 115951 561947 116019 562003
rect 116075 561947 116143 562003
rect 116199 561947 116267 562003
rect 116323 561947 116391 562003
rect 116447 561947 116515 562003
rect 116571 561947 116639 562003
rect 116695 561947 116763 562003
rect 116819 561947 116887 562003
rect 116943 561947 117011 562003
rect 117067 561947 117135 562003
rect 117191 561947 117259 562003
rect 117315 561947 117383 562003
rect 117439 561947 117507 562003
rect 117563 561947 117631 562003
rect 117687 561947 117755 562003
rect 117811 561947 117879 562003
rect 117935 561947 118003 562003
rect 118059 561947 118127 562003
rect 118183 561947 118251 562003
rect 118307 561947 118375 562003
rect 118431 561947 118499 562003
rect 118555 561947 118623 562003
rect 118679 561947 118747 562003
rect 118803 561947 118871 562003
rect 118927 561947 118995 562003
rect 119051 561947 119119 562003
rect 119175 561947 119243 562003
rect 119299 561947 119367 562003
rect 119423 561947 119491 562003
rect 119547 561947 119615 562003
rect 119671 561947 119739 562003
rect 119795 561947 119863 562003
rect 119919 561947 119987 562003
rect 120043 561947 120111 562003
rect 120167 561947 120235 562003
rect 120291 561947 120359 562003
rect 120415 561947 120450 562003
rect 114000 561900 120450 561947
rect 128298 562046 128394 562102
rect 128450 562046 128518 562102
rect 128574 562046 128642 562102
rect 128698 562046 128766 562102
rect 128822 562046 128918 562102
rect 128298 561978 128918 562046
rect 128298 561922 128394 561978
rect 128450 561922 128518 561978
rect 128574 561922 128642 561978
rect 128698 561922 128766 561978
rect 128822 561922 128918 561978
rect 101298 550294 101394 550350
rect 101450 550294 101518 550350
rect 101574 550294 101642 550350
rect 101698 550294 101766 550350
rect 101822 550294 101918 550350
rect 101298 550226 101918 550294
rect 101298 550170 101394 550226
rect 101450 550170 101518 550226
rect 101574 550170 101642 550226
rect 101698 550170 101766 550226
rect 101822 550170 101918 550226
rect 101298 550102 101918 550170
rect 101298 550046 101394 550102
rect 101450 550046 101518 550102
rect 101574 550046 101642 550102
rect 101698 550046 101766 550102
rect 101822 550046 101918 550102
rect 101298 549978 101918 550046
rect 101298 549922 101394 549978
rect 101450 549922 101518 549978
rect 101574 549922 101642 549978
rect 101698 549922 101766 549978
rect 101822 549922 101918 549978
rect 101298 547962 101918 549922
rect 128298 544350 128918 561922
rect 132018 598172 132638 598268
rect 132018 598116 132114 598172
rect 132170 598116 132238 598172
rect 132294 598116 132362 598172
rect 132418 598116 132486 598172
rect 132542 598116 132638 598172
rect 132018 598048 132638 598116
rect 132018 597992 132114 598048
rect 132170 597992 132238 598048
rect 132294 597992 132362 598048
rect 132418 597992 132486 598048
rect 132542 597992 132638 598048
rect 132018 597924 132638 597992
rect 132018 597868 132114 597924
rect 132170 597868 132238 597924
rect 132294 597868 132362 597924
rect 132418 597868 132486 597924
rect 132542 597868 132638 597924
rect 132018 597800 132638 597868
rect 132018 597744 132114 597800
rect 132170 597744 132238 597800
rect 132294 597744 132362 597800
rect 132418 597744 132486 597800
rect 132542 597744 132638 597800
rect 132018 586350 132638 597744
rect 132018 586294 132114 586350
rect 132170 586294 132238 586350
rect 132294 586294 132362 586350
rect 132418 586294 132486 586350
rect 132542 586294 132638 586350
rect 132018 586226 132638 586294
rect 132018 586170 132114 586226
rect 132170 586170 132238 586226
rect 132294 586170 132362 586226
rect 132418 586170 132486 586226
rect 132542 586170 132638 586226
rect 132018 586102 132638 586170
rect 132018 586046 132114 586102
rect 132170 586046 132238 586102
rect 132294 586046 132362 586102
rect 132418 586046 132486 586102
rect 132542 586046 132638 586102
rect 132018 585978 132638 586046
rect 132018 585922 132114 585978
rect 132170 585922 132238 585978
rect 132294 585922 132362 585978
rect 132418 585922 132486 585978
rect 132542 585922 132638 585978
rect 132018 568350 132638 585922
rect 132018 568294 132114 568350
rect 132170 568294 132238 568350
rect 132294 568294 132362 568350
rect 132418 568294 132486 568350
rect 132542 568294 132638 568350
rect 132018 568226 132638 568294
rect 132018 568170 132114 568226
rect 132170 568170 132238 568226
rect 132294 568170 132362 568226
rect 132418 568170 132486 568226
rect 132542 568170 132638 568226
rect 132018 568102 132638 568170
rect 132018 568046 132114 568102
rect 132170 568046 132238 568102
rect 132294 568046 132362 568102
rect 132418 568046 132486 568102
rect 132542 568046 132638 568102
rect 132018 567978 132638 568046
rect 132018 567922 132114 567978
rect 132170 567922 132238 567978
rect 132294 567922 132362 567978
rect 132418 567922 132486 567978
rect 132542 567922 132638 567978
rect 132018 550350 132638 567922
rect 132018 550294 132114 550350
rect 132170 550294 132238 550350
rect 132294 550294 132362 550350
rect 132418 550294 132486 550350
rect 132542 550294 132638 550350
rect 132018 550226 132638 550294
rect 132018 550170 132114 550226
rect 132170 550170 132238 550226
rect 132294 550170 132362 550226
rect 132418 550170 132486 550226
rect 132542 550170 132638 550226
rect 132018 550102 132638 550170
rect 132018 550046 132114 550102
rect 132170 550046 132238 550102
rect 132294 550046 132362 550102
rect 132418 550046 132486 550102
rect 132542 550046 132638 550102
rect 132018 549978 132638 550046
rect 132018 549922 132114 549978
rect 132170 549922 132238 549978
rect 132294 549922 132362 549978
rect 132418 549922 132486 549978
rect 132542 549922 132638 549978
rect 132018 544962 132638 549922
rect 159018 597212 159638 598268
rect 159018 597156 159114 597212
rect 159170 597156 159238 597212
rect 159294 597156 159362 597212
rect 159418 597156 159486 597212
rect 159542 597156 159638 597212
rect 159018 597088 159638 597156
rect 159018 597032 159114 597088
rect 159170 597032 159238 597088
rect 159294 597032 159362 597088
rect 159418 597032 159486 597088
rect 159542 597032 159638 597088
rect 159018 596964 159638 597032
rect 159018 596908 159114 596964
rect 159170 596908 159238 596964
rect 159294 596908 159362 596964
rect 159418 596908 159486 596964
rect 159542 596908 159638 596964
rect 159018 596840 159638 596908
rect 159018 596784 159114 596840
rect 159170 596784 159238 596840
rect 159294 596784 159362 596840
rect 159418 596784 159486 596840
rect 159542 596784 159638 596840
rect 159018 580350 159638 596784
rect 159018 580294 159114 580350
rect 159170 580294 159238 580350
rect 159294 580294 159362 580350
rect 159418 580294 159486 580350
rect 159542 580294 159638 580350
rect 159018 580226 159638 580294
rect 159018 580170 159114 580226
rect 159170 580170 159238 580226
rect 159294 580170 159362 580226
rect 159418 580170 159486 580226
rect 159542 580170 159638 580226
rect 159018 580102 159638 580170
rect 159018 580046 159114 580102
rect 159170 580046 159238 580102
rect 159294 580046 159362 580102
rect 159418 580046 159486 580102
rect 159542 580046 159638 580102
rect 159018 579978 159638 580046
rect 159018 579922 159114 579978
rect 159170 579922 159238 579978
rect 159294 579922 159362 579978
rect 159418 579922 159486 579978
rect 159542 579922 159638 579978
rect 159018 562350 159638 579922
rect 159018 562294 159114 562350
rect 159170 562294 159238 562350
rect 159294 562294 159362 562350
rect 159418 562294 159486 562350
rect 159542 562294 159638 562350
rect 159018 562226 159638 562294
rect 159018 562170 159114 562226
rect 159170 562170 159238 562226
rect 159294 562170 159362 562226
rect 159418 562170 159486 562226
rect 159542 562170 159638 562226
rect 159018 562102 159638 562170
rect 159018 562046 159114 562102
rect 159170 562046 159238 562102
rect 159294 562046 159362 562102
rect 159418 562046 159486 562102
rect 159542 562046 159638 562102
rect 159018 561978 159638 562046
rect 159018 561922 159114 561978
rect 159170 561922 159238 561978
rect 159294 561922 159362 561978
rect 159418 561922 159486 561978
rect 159542 561922 159638 561978
rect 97578 544294 97674 544350
rect 97730 544294 97798 544350
rect 97854 544294 97922 544350
rect 97978 544294 98046 544350
rect 98102 544294 98198 544350
rect 97578 544226 98198 544294
rect 97578 544170 97674 544226
rect 97730 544170 97798 544226
rect 97854 544170 97922 544226
rect 97978 544170 98046 544226
rect 98102 544170 98198 544226
rect 97578 544102 98198 544170
rect 97578 544046 97674 544102
rect 97730 544046 97798 544102
rect 97854 544046 97922 544102
rect 97978 544046 98046 544102
rect 98102 544046 98198 544102
rect 100950 544290 101036 544350
rect 100950 544234 100965 544290
rect 101021 544234 101036 544290
rect 100950 544166 101036 544234
rect 100950 544110 100965 544166
rect 101021 544110 101036 544166
rect 100950 544050 101036 544110
rect 101074 544290 101532 544350
rect 101074 544234 101089 544290
rect 101145 544234 101213 544290
rect 101269 544234 101337 544290
rect 101393 544234 101461 544290
rect 101517 544234 101532 544290
rect 101074 544166 101532 544234
rect 101074 544110 101089 544166
rect 101145 544110 101213 544166
rect 101269 544110 101337 544166
rect 101393 544110 101461 544166
rect 101517 544110 101532 544166
rect 101074 544050 101532 544110
rect 101570 544290 102028 544350
rect 101570 544234 101585 544290
rect 101641 544234 101709 544290
rect 101765 544234 101833 544290
rect 101889 544234 101957 544290
rect 102013 544234 102028 544290
rect 101570 544166 102028 544234
rect 101570 544110 101585 544166
rect 101641 544110 101709 544166
rect 101765 544110 101833 544166
rect 101889 544110 101957 544166
rect 102013 544110 102028 544166
rect 101570 544050 102028 544110
rect 102066 544290 102524 544350
rect 102066 544234 102081 544290
rect 102137 544234 102205 544290
rect 102261 544234 102329 544290
rect 102385 544234 102453 544290
rect 102509 544234 102524 544290
rect 102066 544166 102524 544234
rect 102066 544110 102081 544166
rect 102137 544110 102205 544166
rect 102261 544110 102329 544166
rect 102385 544110 102453 544166
rect 102509 544110 102524 544166
rect 102066 544050 102524 544110
rect 102562 544290 103020 544350
rect 102562 544234 102577 544290
rect 102633 544234 102701 544290
rect 102757 544234 102825 544290
rect 102881 544234 102949 544290
rect 103005 544234 103020 544290
rect 102562 544166 103020 544234
rect 102562 544110 102577 544166
rect 102633 544110 102701 544166
rect 102757 544110 102825 544166
rect 102881 544110 102949 544166
rect 103005 544110 103020 544166
rect 102562 544050 103020 544110
rect 103058 544290 103516 544350
rect 103058 544234 103073 544290
rect 103129 544234 103197 544290
rect 103253 544234 103321 544290
rect 103377 544234 103445 544290
rect 103501 544234 103516 544290
rect 103058 544166 103516 544234
rect 103058 544110 103073 544166
rect 103129 544110 103197 544166
rect 103253 544110 103321 544166
rect 103377 544110 103445 544166
rect 103501 544110 103516 544166
rect 103058 544050 103516 544110
rect 103554 544290 104012 544350
rect 103554 544234 103569 544290
rect 103625 544234 103693 544290
rect 103749 544234 103817 544290
rect 103873 544234 103941 544290
rect 103997 544234 104012 544290
rect 103554 544166 104012 544234
rect 103554 544110 103569 544166
rect 103625 544110 103693 544166
rect 103749 544110 103817 544166
rect 103873 544110 103941 544166
rect 103997 544110 104012 544166
rect 103554 544050 104012 544110
rect 104050 544290 104508 544350
rect 104050 544234 104065 544290
rect 104121 544234 104189 544290
rect 104245 544234 104313 544290
rect 104369 544234 104437 544290
rect 104493 544234 104508 544290
rect 104050 544166 104508 544234
rect 104050 544110 104065 544166
rect 104121 544110 104189 544166
rect 104245 544110 104313 544166
rect 104369 544110 104437 544166
rect 104493 544110 104508 544166
rect 104050 544050 104508 544110
rect 104546 544290 105004 544350
rect 104546 544234 104561 544290
rect 104617 544234 104685 544290
rect 104741 544234 104809 544290
rect 104865 544234 104933 544290
rect 104989 544234 105004 544290
rect 104546 544166 105004 544234
rect 104546 544110 104561 544166
rect 104617 544110 104685 544166
rect 104741 544110 104809 544166
rect 104865 544110 104933 544166
rect 104989 544110 105004 544166
rect 104546 544050 105004 544110
rect 105042 544290 105500 544350
rect 105042 544234 105057 544290
rect 105113 544234 105181 544290
rect 105237 544234 105305 544290
rect 105361 544234 105429 544290
rect 105485 544234 105500 544290
rect 105042 544166 105500 544234
rect 105042 544110 105057 544166
rect 105113 544110 105181 544166
rect 105237 544110 105305 544166
rect 105361 544110 105429 544166
rect 105485 544110 105500 544166
rect 105042 544050 105500 544110
rect 105538 544290 105996 544350
rect 105538 544234 105553 544290
rect 105609 544234 105677 544290
rect 105733 544234 105801 544290
rect 105857 544234 105925 544290
rect 105981 544234 105996 544290
rect 105538 544166 105996 544234
rect 105538 544110 105553 544166
rect 105609 544110 105677 544166
rect 105733 544110 105801 544166
rect 105857 544110 105925 544166
rect 105981 544110 105996 544166
rect 105538 544050 105996 544110
rect 106034 544290 106492 544350
rect 106034 544234 106049 544290
rect 106105 544234 106173 544290
rect 106229 544234 106297 544290
rect 106353 544234 106421 544290
rect 106477 544234 106492 544290
rect 106034 544166 106492 544234
rect 106034 544110 106049 544166
rect 106105 544110 106173 544166
rect 106229 544110 106297 544166
rect 106353 544110 106421 544166
rect 106477 544110 106492 544166
rect 106034 544050 106492 544110
rect 106530 544290 106988 544350
rect 106530 544234 106545 544290
rect 106601 544234 106669 544290
rect 106725 544234 106793 544290
rect 106849 544234 106917 544290
rect 106973 544234 106988 544290
rect 106530 544166 106988 544234
rect 106530 544110 106545 544166
rect 106601 544110 106669 544166
rect 106725 544110 106793 544166
rect 106849 544110 106917 544166
rect 106973 544110 106988 544166
rect 106530 544050 106988 544110
rect 107026 544290 107484 544350
rect 107026 544234 107041 544290
rect 107097 544234 107165 544290
rect 107221 544234 107289 544290
rect 107345 544234 107413 544290
rect 107469 544234 107484 544290
rect 107026 544166 107484 544234
rect 107026 544110 107041 544166
rect 107097 544110 107165 544166
rect 107221 544110 107289 544166
rect 107345 544110 107413 544166
rect 107469 544110 107484 544166
rect 107026 544050 107484 544110
rect 107522 544290 107980 544350
rect 107522 544234 107537 544290
rect 107593 544234 107661 544290
rect 107717 544234 107785 544290
rect 107841 544234 107909 544290
rect 107965 544234 107980 544290
rect 107522 544166 107980 544234
rect 107522 544110 107537 544166
rect 107593 544110 107661 544166
rect 107717 544110 107785 544166
rect 107841 544110 107909 544166
rect 107965 544110 107980 544166
rect 107522 544050 107980 544110
rect 108018 544290 108476 544350
rect 108018 544234 108033 544290
rect 108089 544234 108157 544290
rect 108213 544234 108281 544290
rect 108337 544234 108405 544290
rect 108461 544234 108476 544290
rect 108018 544166 108476 544234
rect 108018 544110 108033 544166
rect 108089 544110 108157 544166
rect 108213 544110 108281 544166
rect 108337 544110 108405 544166
rect 108461 544110 108476 544166
rect 108018 544050 108476 544110
rect 108514 544290 108972 544350
rect 108514 544234 108529 544290
rect 108585 544234 108653 544290
rect 108709 544234 108777 544290
rect 108833 544234 108901 544290
rect 108957 544234 108972 544290
rect 108514 544166 108972 544234
rect 108514 544110 108529 544166
rect 108585 544110 108653 544166
rect 108709 544110 108777 544166
rect 108833 544110 108901 544166
rect 108957 544110 108972 544166
rect 108514 544050 108972 544110
rect 109010 544290 109468 544350
rect 109010 544234 109025 544290
rect 109081 544234 109149 544290
rect 109205 544234 109273 544290
rect 109329 544234 109397 544290
rect 109453 544234 109468 544290
rect 109010 544166 109468 544234
rect 109010 544110 109025 544166
rect 109081 544110 109149 544166
rect 109205 544110 109273 544166
rect 109329 544110 109397 544166
rect 109453 544110 109468 544166
rect 109010 544050 109468 544110
rect 109506 544290 109964 544350
rect 109506 544234 109521 544290
rect 109577 544234 109645 544290
rect 109701 544234 109769 544290
rect 109825 544234 109893 544290
rect 109949 544234 109964 544290
rect 109506 544166 109964 544234
rect 109506 544110 109521 544166
rect 109577 544110 109645 544166
rect 109701 544110 109769 544166
rect 109825 544110 109893 544166
rect 109949 544110 109964 544166
rect 109506 544050 109964 544110
rect 110002 544290 110460 544350
rect 110002 544234 110017 544290
rect 110073 544234 110141 544290
rect 110197 544234 110265 544290
rect 110321 544234 110389 544290
rect 110445 544234 110460 544290
rect 110002 544166 110460 544234
rect 110002 544110 110017 544166
rect 110073 544110 110141 544166
rect 110197 544110 110265 544166
rect 110321 544110 110389 544166
rect 110445 544110 110460 544166
rect 110002 544050 110460 544110
rect 110498 544290 110956 544350
rect 110498 544234 110513 544290
rect 110569 544234 110637 544290
rect 110693 544234 110761 544290
rect 110817 544234 110885 544290
rect 110941 544234 110956 544290
rect 110498 544166 110956 544234
rect 110498 544110 110513 544166
rect 110569 544110 110637 544166
rect 110693 544110 110761 544166
rect 110817 544110 110885 544166
rect 110941 544110 110956 544166
rect 110498 544050 110956 544110
rect 110994 544290 111452 544350
rect 110994 544234 111009 544290
rect 111065 544234 111133 544290
rect 111189 544234 111257 544290
rect 111313 544234 111381 544290
rect 111437 544234 111452 544290
rect 110994 544166 111452 544234
rect 110994 544110 111009 544166
rect 111065 544110 111133 544166
rect 111189 544110 111257 544166
rect 111313 544110 111381 544166
rect 111437 544110 111452 544166
rect 110994 544050 111452 544110
rect 111490 544290 111948 544350
rect 111490 544234 111505 544290
rect 111561 544234 111629 544290
rect 111685 544234 111753 544290
rect 111809 544234 111877 544290
rect 111933 544234 111948 544290
rect 111490 544166 111948 544234
rect 111490 544110 111505 544166
rect 111561 544110 111629 544166
rect 111685 544110 111753 544166
rect 111809 544110 111877 544166
rect 111933 544110 111948 544166
rect 111490 544050 111948 544110
rect 111986 544290 112444 544350
rect 111986 544234 112001 544290
rect 112057 544234 112125 544290
rect 112181 544234 112249 544290
rect 112305 544234 112373 544290
rect 112429 544234 112444 544290
rect 111986 544166 112444 544234
rect 111986 544110 112001 544166
rect 112057 544110 112125 544166
rect 112181 544110 112249 544166
rect 112305 544110 112373 544166
rect 112429 544110 112444 544166
rect 111986 544050 112444 544110
rect 112482 544290 112940 544350
rect 112482 544234 112497 544290
rect 112553 544234 112621 544290
rect 112677 544234 112745 544290
rect 112801 544234 112869 544290
rect 112925 544234 112940 544290
rect 112482 544166 112940 544234
rect 112482 544110 112497 544166
rect 112553 544110 112621 544166
rect 112677 544110 112745 544166
rect 112801 544110 112869 544166
rect 112925 544110 112940 544166
rect 112482 544050 112940 544110
rect 112978 544290 113436 544350
rect 112978 544234 112993 544290
rect 113049 544234 113117 544290
rect 113173 544234 113241 544290
rect 113297 544234 113365 544290
rect 113421 544234 113436 544290
rect 112978 544166 113436 544234
rect 112978 544110 112993 544166
rect 113049 544110 113117 544166
rect 113173 544110 113241 544166
rect 113297 544110 113365 544166
rect 113421 544110 113436 544166
rect 112978 544050 113436 544110
rect 113474 544290 113932 544350
rect 113474 544234 113489 544290
rect 113545 544234 113613 544290
rect 113669 544234 113737 544290
rect 113793 544234 113861 544290
rect 113917 544234 113932 544290
rect 113474 544166 113932 544234
rect 113474 544110 113489 544166
rect 113545 544110 113613 544166
rect 113669 544110 113737 544166
rect 113793 544110 113861 544166
rect 113917 544110 113932 544166
rect 113474 544050 113932 544110
rect 113970 544290 114428 544350
rect 113970 544234 113985 544290
rect 114041 544234 114109 544290
rect 114165 544234 114233 544290
rect 114289 544234 114357 544290
rect 114413 544234 114428 544290
rect 113970 544166 114428 544234
rect 113970 544110 113985 544166
rect 114041 544110 114109 544166
rect 114165 544110 114233 544166
rect 114289 544110 114357 544166
rect 114413 544110 114428 544166
rect 113970 544050 114428 544110
rect 114466 544290 114924 544350
rect 114466 544234 114481 544290
rect 114537 544234 114605 544290
rect 114661 544234 114729 544290
rect 114785 544234 114853 544290
rect 114909 544234 114924 544290
rect 114466 544166 114924 544234
rect 114466 544110 114481 544166
rect 114537 544110 114605 544166
rect 114661 544110 114729 544166
rect 114785 544110 114853 544166
rect 114909 544110 114924 544166
rect 114466 544050 114924 544110
rect 114962 544290 115420 544350
rect 114962 544234 114977 544290
rect 115033 544234 115101 544290
rect 115157 544234 115225 544290
rect 115281 544234 115349 544290
rect 115405 544234 115420 544290
rect 114962 544166 115420 544234
rect 114962 544110 114977 544166
rect 115033 544110 115101 544166
rect 115157 544110 115225 544166
rect 115281 544110 115349 544166
rect 115405 544110 115420 544166
rect 114962 544050 115420 544110
rect 115458 544290 115916 544350
rect 115458 544234 115473 544290
rect 115529 544234 115597 544290
rect 115653 544234 115721 544290
rect 115777 544234 115845 544290
rect 115901 544234 115916 544290
rect 115458 544166 115916 544234
rect 115458 544110 115473 544166
rect 115529 544110 115597 544166
rect 115653 544110 115721 544166
rect 115777 544110 115845 544166
rect 115901 544110 115916 544166
rect 115458 544050 115916 544110
rect 115954 544290 116412 544350
rect 115954 544234 115969 544290
rect 116025 544234 116093 544290
rect 116149 544234 116217 544290
rect 116273 544234 116341 544290
rect 116397 544234 116412 544290
rect 115954 544166 116412 544234
rect 115954 544110 115969 544166
rect 116025 544110 116093 544166
rect 116149 544110 116217 544166
rect 116273 544110 116341 544166
rect 116397 544110 116412 544166
rect 115954 544050 116412 544110
rect 116450 544290 116908 544350
rect 116450 544234 116465 544290
rect 116521 544234 116589 544290
rect 116645 544234 116713 544290
rect 116769 544234 116837 544290
rect 116893 544234 116908 544290
rect 116450 544166 116908 544234
rect 116450 544110 116465 544166
rect 116521 544110 116589 544166
rect 116645 544110 116713 544166
rect 116769 544110 116837 544166
rect 116893 544110 116908 544166
rect 116450 544050 116908 544110
rect 116946 544290 117404 544350
rect 116946 544234 116961 544290
rect 117017 544234 117085 544290
rect 117141 544234 117209 544290
rect 117265 544234 117333 544290
rect 117389 544234 117404 544290
rect 116946 544166 117404 544234
rect 116946 544110 116961 544166
rect 117017 544110 117085 544166
rect 117141 544110 117209 544166
rect 117265 544110 117333 544166
rect 117389 544110 117404 544166
rect 116946 544050 117404 544110
rect 117442 544290 117900 544350
rect 117442 544234 117457 544290
rect 117513 544234 117581 544290
rect 117637 544234 117705 544290
rect 117761 544234 117829 544290
rect 117885 544234 117900 544290
rect 117442 544166 117900 544234
rect 117442 544110 117457 544166
rect 117513 544110 117581 544166
rect 117637 544110 117705 544166
rect 117761 544110 117829 544166
rect 117885 544110 117900 544166
rect 117442 544050 117900 544110
rect 128298 544294 128394 544350
rect 128450 544294 128518 544350
rect 128574 544294 128642 544350
rect 128698 544294 128766 544350
rect 128822 544294 128918 544350
rect 128298 544226 128918 544294
rect 128298 544170 128394 544226
rect 128450 544170 128518 544226
rect 128574 544170 128642 544226
rect 128698 544170 128766 544226
rect 128822 544170 128918 544226
rect 128298 544102 128918 544170
rect 97578 543978 98198 544046
rect 97578 543922 97674 543978
rect 97730 543922 97798 543978
rect 97854 543922 97922 543978
rect 97978 543922 98046 543978
rect 98102 543922 98198 543978
rect 97578 542112 98198 543922
rect 128298 544046 128394 544102
rect 128450 544046 128518 544102
rect 128574 544046 128642 544102
rect 128698 544046 128766 544102
rect 128822 544046 128918 544102
rect 128298 543978 128918 544046
rect 128298 543922 128394 543978
rect 128450 543922 128518 543978
rect 128574 543922 128642 543978
rect 128698 543922 128766 543978
rect 128822 543922 128918 543978
rect 100800 543891 117750 543900
rect 100800 543835 100823 543891
rect 100879 543835 100927 543891
rect 100983 543835 101031 543891
rect 101087 543835 101135 543891
rect 101191 543835 101239 543891
rect 101295 543835 101343 543891
rect 101399 543835 101447 543891
rect 101503 543835 101551 543891
rect 101607 543835 101655 543891
rect 101711 543835 101759 543891
rect 101815 543835 101863 543891
rect 101919 543835 101967 543891
rect 102023 543835 102071 543891
rect 102127 543835 102175 543891
rect 102231 543835 102279 543891
rect 102335 543835 102383 543891
rect 102439 543835 102487 543891
rect 102543 543835 102591 543891
rect 102647 543835 102695 543891
rect 102751 543835 102799 543891
rect 102855 543835 102903 543891
rect 102959 543835 103007 543891
rect 103063 543835 103111 543891
rect 103167 543835 103215 543891
rect 103271 543835 103319 543891
rect 103375 543835 103423 543891
rect 103479 543835 103527 543891
rect 103583 543835 103631 543891
rect 103687 543835 103735 543891
rect 103791 543835 103839 543891
rect 103895 543835 103943 543891
rect 103999 543835 104047 543891
rect 104103 543835 104151 543891
rect 104207 543835 104255 543891
rect 104311 543835 104359 543891
rect 104415 543835 104463 543891
rect 104519 543835 104567 543891
rect 104623 543835 104671 543891
rect 104727 543835 104775 543891
rect 104831 543835 104879 543891
rect 104935 543835 104983 543891
rect 105039 543835 105087 543891
rect 105143 543835 105191 543891
rect 105247 543835 105295 543891
rect 105351 543835 105399 543891
rect 105455 543835 105503 543891
rect 105559 543835 105607 543891
rect 105663 543835 105711 543891
rect 105767 543835 105815 543891
rect 105871 543835 105919 543891
rect 105975 543835 106023 543891
rect 106079 543835 106127 543891
rect 106183 543835 106231 543891
rect 106287 543835 106335 543891
rect 106391 543835 106439 543891
rect 106495 543835 106543 543891
rect 106599 543835 106647 543891
rect 106703 543835 106751 543891
rect 106807 543835 106855 543891
rect 106911 543835 106959 543891
rect 107015 543835 107063 543891
rect 107119 543835 107167 543891
rect 107223 543835 107271 543891
rect 107327 543835 107375 543891
rect 107431 543835 107479 543891
rect 107535 543835 107583 543891
rect 107639 543835 107687 543891
rect 107743 543835 107791 543891
rect 107847 543835 107895 543891
rect 107951 543835 107999 543891
rect 108055 543835 108103 543891
rect 108159 543835 108207 543891
rect 108263 543835 108311 543891
rect 108367 543835 108415 543891
rect 108471 543835 108519 543891
rect 108575 543835 108623 543891
rect 108679 543835 108727 543891
rect 108783 543835 108831 543891
rect 108887 543835 108935 543891
rect 108991 543835 109039 543891
rect 109095 543835 109143 543891
rect 109199 543835 109247 543891
rect 109303 543835 109351 543891
rect 109407 543835 109455 543891
rect 109511 543835 109559 543891
rect 109615 543835 109663 543891
rect 109719 543835 109767 543891
rect 109823 543835 109871 543891
rect 109927 543835 109975 543891
rect 110031 543835 110079 543891
rect 110135 543835 110183 543891
rect 110239 543835 110287 543891
rect 110343 543835 110391 543891
rect 110447 543835 110495 543891
rect 110551 543835 110599 543891
rect 110655 543835 110703 543891
rect 110759 543835 110807 543891
rect 110863 543835 110911 543891
rect 110967 543835 111015 543891
rect 111071 543835 111119 543891
rect 111175 543835 111223 543891
rect 111279 543835 111327 543891
rect 111383 543835 111431 543891
rect 111487 543835 111535 543891
rect 111591 543835 111639 543891
rect 111695 543835 111743 543891
rect 111799 543835 111847 543891
rect 111903 543835 111951 543891
rect 112007 543835 112055 543891
rect 112111 543835 112159 543891
rect 112215 543835 112263 543891
rect 112319 543835 112367 543891
rect 112423 543835 112471 543891
rect 112527 543835 112575 543891
rect 112631 543835 112679 543891
rect 112735 543835 112783 543891
rect 112839 543835 112887 543891
rect 112943 543835 112991 543891
rect 113047 543835 113095 543891
rect 113151 543835 113199 543891
rect 113255 543835 113303 543891
rect 113359 543835 113407 543891
rect 113463 543835 113511 543891
rect 113567 543835 113615 543891
rect 113671 543835 113719 543891
rect 113775 543835 113823 543891
rect 113879 543835 113927 543891
rect 113983 543835 114031 543891
rect 114087 543835 114135 543891
rect 114191 543835 114239 543891
rect 114295 543835 114343 543891
rect 114399 543835 114447 543891
rect 114503 543835 114551 543891
rect 114607 543835 114655 543891
rect 114711 543835 114759 543891
rect 114815 543835 114863 543891
rect 114919 543835 114967 543891
rect 115023 543835 115071 543891
rect 115127 543835 115175 543891
rect 115231 543835 115279 543891
rect 115335 543835 115383 543891
rect 115439 543835 115487 543891
rect 115543 543835 115591 543891
rect 115647 543835 115695 543891
rect 115751 543835 115799 543891
rect 115855 543835 115903 543891
rect 115959 543835 116007 543891
rect 116063 543835 116111 543891
rect 116167 543835 116215 543891
rect 116271 543835 116319 543891
rect 116375 543835 116423 543891
rect 116479 543835 116527 543891
rect 116583 543835 116631 543891
rect 116687 543835 116735 543891
rect 116791 543835 116839 543891
rect 116895 543835 116943 543891
rect 116999 543835 117047 543891
rect 117103 543835 117151 543891
rect 117207 543835 117255 543891
rect 117311 543835 117359 543891
rect 117415 543835 117463 543891
rect 117519 543835 117567 543891
rect 117623 543835 117671 543891
rect 117727 543835 117750 543891
rect 100800 543826 117750 543835
rect 128298 543612 128918 543922
rect 159018 544350 159638 561922
rect 159018 544294 159114 544350
rect 159170 544294 159238 544350
rect 159294 544294 159362 544350
rect 159418 544294 159486 544350
rect 159542 544294 159638 544350
rect 159018 544226 159638 544294
rect 159018 544170 159114 544226
rect 159170 544170 159238 544226
rect 159294 544170 159362 544226
rect 159418 544170 159486 544226
rect 159542 544170 159638 544226
rect 159018 544102 159638 544170
rect 159018 544046 159114 544102
rect 159170 544046 159238 544102
rect 159294 544046 159362 544102
rect 159418 544046 159486 544102
rect 159542 544046 159638 544102
rect 159018 543978 159638 544046
rect 159018 543922 159114 543978
rect 159170 543922 159238 543978
rect 159294 543922 159362 543978
rect 159418 543922 159486 543978
rect 159542 543922 159638 543978
rect 39858 532294 39954 532350
rect 40010 532294 40078 532350
rect 40134 532294 40202 532350
rect 40258 532294 40326 532350
rect 40382 532294 40478 532350
rect 39858 532226 40478 532294
rect 39858 532170 39954 532226
rect 40010 532170 40078 532226
rect 40134 532170 40202 532226
rect 40258 532170 40326 532226
rect 40382 532170 40478 532226
rect 69450 532303 78300 532350
rect 69450 532247 69507 532303
rect 69563 532247 69631 532303
rect 69687 532247 69755 532303
rect 69811 532247 69879 532303
rect 69935 532247 70003 532303
rect 70059 532247 70127 532303
rect 70183 532247 70251 532303
rect 70307 532247 70375 532303
rect 70431 532247 70499 532303
rect 70555 532247 70623 532303
rect 70679 532247 70747 532303
rect 70803 532247 70871 532303
rect 70927 532247 70995 532303
rect 71051 532247 71119 532303
rect 71175 532247 71243 532303
rect 71299 532247 71367 532303
rect 71423 532247 71491 532303
rect 71547 532247 71615 532303
rect 71671 532247 71739 532303
rect 71795 532247 71863 532303
rect 71919 532247 71987 532303
rect 72043 532247 72111 532303
rect 72167 532247 72235 532303
rect 72291 532247 72359 532303
rect 72415 532247 72483 532303
rect 72539 532247 72607 532303
rect 72663 532247 72731 532303
rect 72787 532247 72855 532303
rect 72911 532247 72979 532303
rect 73035 532247 73103 532303
rect 73159 532247 73227 532303
rect 73283 532247 73351 532303
rect 73407 532247 73475 532303
rect 73531 532247 73599 532303
rect 73655 532247 73723 532303
rect 73779 532247 73847 532303
rect 73903 532247 73971 532303
rect 74027 532247 74095 532303
rect 74151 532247 74219 532303
rect 74275 532247 74343 532303
rect 74399 532247 74467 532303
rect 74523 532247 74591 532303
rect 74647 532247 74715 532303
rect 74771 532247 74839 532303
rect 74895 532247 74963 532303
rect 75019 532247 75087 532303
rect 75143 532247 75211 532303
rect 75267 532247 75335 532303
rect 75391 532247 75459 532303
rect 75515 532247 75583 532303
rect 75639 532247 75707 532303
rect 75763 532247 75831 532303
rect 75887 532247 75955 532303
rect 76011 532247 76079 532303
rect 76135 532247 76203 532303
rect 76259 532247 76327 532303
rect 76383 532247 76451 532303
rect 76507 532247 76575 532303
rect 76631 532247 76699 532303
rect 76755 532247 76823 532303
rect 76879 532247 76947 532303
rect 77003 532247 77071 532303
rect 77127 532247 77195 532303
rect 77251 532247 77319 532303
rect 77375 532247 77443 532303
rect 77499 532247 77567 532303
rect 77623 532247 77691 532303
rect 77747 532247 77815 532303
rect 77871 532247 77939 532303
rect 77995 532247 78063 532303
rect 78119 532247 78187 532303
rect 78243 532247 78300 532303
rect 69450 532200 78300 532247
rect 39858 532102 40478 532170
rect 39858 532046 39954 532102
rect 40010 532046 40078 532102
rect 40134 532046 40202 532102
rect 40258 532046 40326 532102
rect 40382 532046 40478 532102
rect 39858 531978 40478 532046
rect 39858 531922 39954 531978
rect 40010 531922 40078 531978
rect 40134 531922 40202 531978
rect 40258 531922 40326 531978
rect 40382 531922 40478 531978
rect 39858 514350 40478 531922
rect 69150 532003 69268 532050
rect 69150 531947 69181 532003
rect 69237 531947 69268 532003
rect 69150 531900 69268 531947
rect 69274 532003 69764 532050
rect 69274 531947 69305 532003
rect 69361 531947 69429 532003
rect 69485 531947 69553 532003
rect 69609 531947 69677 532003
rect 69733 531947 69764 532003
rect 69274 531900 69764 531947
rect 69770 532003 70260 532050
rect 69770 531947 69801 532003
rect 69857 531947 69925 532003
rect 69981 531947 70049 532003
rect 70105 531947 70173 532003
rect 70229 531947 70260 532003
rect 69770 531900 70260 531947
rect 70266 532003 70756 532050
rect 70266 531947 70297 532003
rect 70353 531947 70421 532003
rect 70477 531947 70545 532003
rect 70601 531947 70669 532003
rect 70725 531947 70756 532003
rect 70266 531900 70756 531947
rect 70762 532003 71252 532050
rect 70762 531947 70793 532003
rect 70849 531947 70917 532003
rect 70973 531947 71041 532003
rect 71097 531947 71165 532003
rect 71221 531947 71252 532003
rect 70762 531900 71252 531947
rect 71258 532003 71748 532050
rect 71258 531947 71289 532003
rect 71345 531947 71413 532003
rect 71469 531947 71537 532003
rect 71593 531947 71661 532003
rect 71717 531947 71748 532003
rect 71258 531900 71748 531947
rect 71754 532003 72244 532050
rect 71754 531947 71785 532003
rect 71841 531947 71909 532003
rect 71965 531947 72033 532003
rect 72089 531947 72157 532003
rect 72213 531947 72244 532003
rect 71754 531900 72244 531947
rect 72250 532003 72740 532050
rect 72250 531947 72281 532003
rect 72337 531947 72405 532003
rect 72461 531947 72529 532003
rect 72585 531947 72653 532003
rect 72709 531947 72740 532003
rect 72250 531900 72740 531947
rect 72746 532003 73236 532050
rect 72746 531947 72777 532003
rect 72833 531947 72901 532003
rect 72957 531947 73025 532003
rect 73081 531947 73149 532003
rect 73205 531947 73236 532003
rect 72746 531900 73236 531947
rect 73242 532003 73732 532050
rect 73242 531947 73273 532003
rect 73329 531947 73397 532003
rect 73453 531947 73521 532003
rect 73577 531947 73645 532003
rect 73701 531947 73732 532003
rect 73242 531900 73732 531947
rect 73738 532003 74228 532050
rect 73738 531947 73769 532003
rect 73825 531947 73893 532003
rect 73949 531947 74017 532003
rect 74073 531947 74141 532003
rect 74197 531947 74228 532003
rect 73738 531900 74228 531947
rect 74234 532003 74724 532050
rect 74234 531947 74265 532003
rect 74321 531947 74389 532003
rect 74445 531947 74513 532003
rect 74569 531947 74637 532003
rect 74693 531947 74724 532003
rect 74234 531900 74724 531947
rect 74730 532003 75220 532050
rect 74730 531947 74761 532003
rect 74817 531947 74885 532003
rect 74941 531947 75009 532003
rect 75065 531947 75133 532003
rect 75189 531947 75220 532003
rect 74730 531900 75220 531947
rect 75226 532003 75716 532050
rect 75226 531947 75257 532003
rect 75313 531947 75381 532003
rect 75437 531947 75505 532003
rect 75561 531947 75629 532003
rect 75685 531947 75716 532003
rect 75226 531900 75716 531947
rect 75722 532003 76212 532050
rect 75722 531947 75753 532003
rect 75809 531947 75877 532003
rect 75933 531947 76001 532003
rect 76057 531947 76125 532003
rect 76181 531947 76212 532003
rect 75722 531900 76212 531947
rect 76218 532003 76708 532050
rect 76218 531947 76249 532003
rect 76305 531947 76373 532003
rect 76429 531947 76497 532003
rect 76553 531947 76621 532003
rect 76677 531947 76708 532003
rect 76218 531900 76708 531947
rect 76714 532003 77204 532050
rect 76714 531947 76745 532003
rect 76801 531947 76869 532003
rect 76925 531947 76993 532003
rect 77049 531947 77117 532003
rect 77173 531947 77204 532003
rect 76714 531900 77204 531947
rect 77210 532003 77700 532050
rect 77210 531947 77241 532003
rect 77297 531947 77365 532003
rect 77421 531947 77489 532003
rect 77545 531947 77613 532003
rect 77669 531947 77700 532003
rect 77210 531900 77700 531947
rect 159018 526350 159638 543922
rect 159018 526294 159114 526350
rect 159170 526294 159238 526350
rect 159294 526294 159362 526350
rect 159418 526294 159486 526350
rect 159542 526294 159638 526350
rect 159018 526226 159638 526294
rect 91350 526153 91840 526200
rect 91350 526097 91381 526153
rect 91437 526097 91505 526153
rect 91561 526097 91629 526153
rect 91685 526097 91753 526153
rect 91809 526097 91840 526153
rect 91350 526050 91840 526097
rect 91846 526153 92336 526200
rect 91846 526097 91877 526153
rect 91933 526097 92001 526153
rect 92057 526097 92125 526153
rect 92181 526097 92249 526153
rect 92305 526097 92336 526153
rect 91846 526050 92336 526097
rect 92342 526153 92832 526200
rect 92342 526097 92373 526153
rect 92429 526097 92497 526153
rect 92553 526097 92621 526153
rect 92677 526097 92745 526153
rect 92801 526097 92832 526153
rect 92342 526050 92832 526097
rect 92838 526153 93328 526200
rect 92838 526097 92869 526153
rect 92925 526097 92993 526153
rect 93049 526097 93117 526153
rect 93173 526097 93241 526153
rect 93297 526097 93328 526153
rect 92838 526050 93328 526097
rect 93334 526153 93824 526200
rect 93334 526097 93365 526153
rect 93421 526097 93489 526153
rect 93545 526097 93613 526153
rect 93669 526097 93737 526153
rect 93793 526097 93824 526153
rect 93334 526050 93824 526097
rect 93830 526153 94320 526200
rect 93830 526097 93861 526153
rect 93917 526097 93985 526153
rect 94041 526097 94109 526153
rect 94165 526097 94233 526153
rect 94289 526097 94320 526153
rect 93830 526050 94320 526097
rect 94326 526153 94816 526200
rect 94326 526097 94357 526153
rect 94413 526097 94481 526153
rect 94537 526097 94605 526153
rect 94661 526097 94729 526153
rect 94785 526097 94816 526153
rect 94326 526050 94816 526097
rect 94822 526153 95312 526200
rect 94822 526097 94853 526153
rect 94909 526097 94977 526153
rect 95033 526097 95101 526153
rect 95157 526097 95225 526153
rect 95281 526097 95312 526153
rect 94822 526050 95312 526097
rect 95318 526153 95808 526200
rect 95318 526097 95349 526153
rect 95405 526097 95473 526153
rect 95529 526097 95597 526153
rect 95653 526097 95721 526153
rect 95777 526097 95808 526153
rect 95318 526050 95808 526097
rect 95814 526153 96304 526200
rect 95814 526097 95845 526153
rect 95901 526097 95969 526153
rect 96025 526097 96093 526153
rect 96149 526097 96217 526153
rect 96273 526097 96304 526153
rect 95814 526050 96304 526097
rect 96310 526153 96800 526200
rect 96310 526097 96341 526153
rect 96397 526097 96465 526153
rect 96521 526097 96589 526153
rect 96645 526097 96713 526153
rect 96769 526097 96800 526153
rect 96310 526050 96800 526097
rect 96806 526153 97296 526200
rect 96806 526097 96837 526153
rect 96893 526097 96961 526153
rect 97017 526097 97085 526153
rect 97141 526097 97209 526153
rect 97265 526097 97296 526153
rect 96806 526050 97296 526097
rect 97302 526153 97792 526200
rect 97302 526097 97333 526153
rect 97389 526097 97457 526153
rect 97513 526097 97581 526153
rect 97637 526097 97705 526153
rect 97761 526097 97792 526153
rect 97302 526050 97792 526097
rect 97798 526153 98288 526200
rect 97798 526097 97829 526153
rect 97885 526097 97953 526153
rect 98009 526097 98077 526153
rect 98133 526097 98201 526153
rect 98257 526097 98288 526153
rect 97798 526050 98288 526097
rect 98294 526153 98784 526200
rect 98294 526097 98325 526153
rect 98381 526097 98449 526153
rect 98505 526097 98573 526153
rect 98629 526097 98697 526153
rect 98753 526097 98784 526153
rect 98294 526050 98784 526097
rect 98790 526153 99280 526200
rect 98790 526097 98821 526153
rect 98877 526097 98945 526153
rect 99001 526097 99069 526153
rect 99125 526097 99193 526153
rect 99249 526097 99280 526153
rect 98790 526050 99280 526097
rect 99286 526153 99776 526200
rect 99286 526097 99317 526153
rect 99373 526097 99441 526153
rect 99497 526097 99565 526153
rect 99621 526097 99689 526153
rect 99745 526097 99776 526153
rect 99286 526050 99776 526097
rect 99782 526153 100272 526200
rect 99782 526097 99813 526153
rect 99869 526097 99937 526153
rect 99993 526097 100061 526153
rect 100117 526097 100185 526153
rect 100241 526097 100272 526153
rect 99782 526050 100272 526097
rect 100278 526153 100768 526200
rect 100278 526097 100309 526153
rect 100365 526097 100433 526153
rect 100489 526097 100557 526153
rect 100613 526097 100681 526153
rect 100737 526097 100768 526153
rect 100278 526050 100768 526097
rect 100774 526153 101264 526200
rect 100774 526097 100805 526153
rect 100861 526097 100929 526153
rect 100985 526097 101053 526153
rect 101109 526097 101177 526153
rect 101233 526097 101264 526153
rect 100774 526050 101264 526097
rect 101270 526153 101760 526200
rect 101270 526097 101301 526153
rect 101357 526097 101425 526153
rect 101481 526097 101549 526153
rect 101605 526097 101673 526153
rect 101729 526097 101760 526153
rect 101270 526050 101760 526097
rect 101766 526153 102256 526200
rect 101766 526097 101797 526153
rect 101853 526097 101921 526153
rect 101977 526097 102045 526153
rect 102101 526097 102169 526153
rect 102225 526097 102256 526153
rect 101766 526050 102256 526097
rect 102262 526153 102752 526200
rect 102262 526097 102293 526153
rect 102349 526097 102417 526153
rect 102473 526097 102541 526153
rect 102597 526097 102665 526153
rect 102721 526097 102752 526153
rect 102262 526050 102752 526097
rect 102758 526153 103248 526200
rect 102758 526097 102789 526153
rect 102845 526097 102913 526153
rect 102969 526097 103037 526153
rect 103093 526097 103161 526153
rect 103217 526097 103248 526153
rect 102758 526050 103248 526097
rect 103254 526153 103744 526200
rect 103254 526097 103285 526153
rect 103341 526097 103409 526153
rect 103465 526097 103533 526153
rect 103589 526097 103657 526153
rect 103713 526097 103744 526153
rect 103254 526050 103744 526097
rect 103750 526153 104240 526200
rect 103750 526097 103781 526153
rect 103837 526097 103905 526153
rect 103961 526097 104029 526153
rect 104085 526097 104153 526153
rect 104209 526097 104240 526153
rect 103750 526050 104240 526097
rect 104246 526153 104736 526200
rect 104246 526097 104277 526153
rect 104333 526097 104401 526153
rect 104457 526097 104525 526153
rect 104581 526097 104649 526153
rect 104705 526097 104736 526153
rect 104246 526050 104736 526097
rect 104742 526153 105232 526200
rect 104742 526097 104773 526153
rect 104829 526097 104897 526153
rect 104953 526097 105021 526153
rect 105077 526097 105145 526153
rect 105201 526097 105232 526153
rect 104742 526050 105232 526097
rect 105238 526153 105728 526200
rect 105238 526097 105269 526153
rect 105325 526097 105393 526153
rect 105449 526097 105517 526153
rect 105573 526097 105641 526153
rect 105697 526097 105728 526153
rect 105238 526050 105728 526097
rect 105734 526153 106224 526200
rect 105734 526097 105765 526153
rect 105821 526097 105889 526153
rect 105945 526097 106013 526153
rect 106069 526097 106137 526153
rect 106193 526097 106224 526153
rect 105734 526050 106224 526097
rect 106230 526153 106720 526200
rect 106230 526097 106261 526153
rect 106317 526097 106385 526153
rect 106441 526097 106509 526153
rect 106565 526097 106633 526153
rect 106689 526097 106720 526153
rect 106230 526050 106720 526097
rect 106726 526153 107216 526200
rect 106726 526097 106757 526153
rect 106813 526097 106881 526153
rect 106937 526097 107005 526153
rect 107061 526097 107129 526153
rect 107185 526097 107216 526153
rect 106726 526050 107216 526097
rect 107222 526153 107712 526200
rect 107222 526097 107253 526153
rect 107309 526097 107377 526153
rect 107433 526097 107501 526153
rect 107557 526097 107625 526153
rect 107681 526097 107712 526153
rect 107222 526050 107712 526097
rect 107718 526153 108208 526200
rect 107718 526097 107749 526153
rect 107805 526097 107873 526153
rect 107929 526097 107997 526153
rect 108053 526097 108121 526153
rect 108177 526097 108208 526153
rect 107718 526050 108208 526097
rect 108214 526153 108704 526200
rect 108214 526097 108245 526153
rect 108301 526097 108369 526153
rect 108425 526097 108493 526153
rect 108549 526097 108617 526153
rect 108673 526097 108704 526153
rect 108214 526050 108704 526097
rect 108710 526153 109200 526200
rect 108710 526097 108741 526153
rect 108797 526097 108865 526153
rect 108921 526097 108989 526153
rect 109045 526097 109113 526153
rect 109169 526097 109200 526153
rect 108710 526050 109200 526097
rect 159018 526170 159114 526226
rect 159170 526170 159238 526226
rect 159294 526170 159362 526226
rect 159418 526170 159486 526226
rect 159542 526170 159638 526226
rect 159018 526102 159638 526170
rect 159018 526046 159114 526102
rect 159170 526046 159238 526102
rect 159294 526046 159362 526102
rect 159418 526046 159486 526102
rect 159542 526046 159638 526102
rect 159018 525978 159638 526046
rect 159018 525922 159114 525978
rect 159170 525922 159238 525978
rect 159294 525922 159362 525978
rect 159418 525922 159486 525978
rect 159542 525922 159638 525978
rect 91200 525891 108900 525900
rect 91200 525835 91234 525891
rect 91290 525835 91338 525891
rect 91394 525835 91442 525891
rect 91498 525835 91546 525891
rect 91602 525835 91650 525891
rect 91706 525835 91754 525891
rect 91810 525835 91858 525891
rect 91914 525835 91962 525891
rect 92018 525835 92066 525891
rect 92122 525835 92170 525891
rect 92226 525835 92274 525891
rect 92330 525835 92378 525891
rect 92434 525835 92482 525891
rect 92538 525835 92586 525891
rect 92642 525835 92690 525891
rect 92746 525835 92794 525891
rect 92850 525835 92898 525891
rect 92954 525835 93002 525891
rect 93058 525835 93106 525891
rect 93162 525835 93210 525891
rect 93266 525835 93314 525891
rect 93370 525835 93418 525891
rect 93474 525835 93522 525891
rect 93578 525835 93626 525891
rect 93682 525835 93730 525891
rect 93786 525835 93834 525891
rect 93890 525835 93938 525891
rect 93994 525835 94042 525891
rect 94098 525835 94146 525891
rect 94202 525835 94250 525891
rect 94306 525835 94354 525891
rect 94410 525835 94458 525891
rect 94514 525835 94562 525891
rect 94618 525835 94666 525891
rect 94722 525835 94770 525891
rect 94826 525835 94874 525891
rect 94930 525835 94978 525891
rect 95034 525835 95082 525891
rect 95138 525835 95186 525891
rect 95242 525835 95290 525891
rect 95346 525835 95394 525891
rect 95450 525835 95498 525891
rect 95554 525835 95602 525891
rect 95658 525835 95706 525891
rect 95762 525835 95810 525891
rect 95866 525835 95914 525891
rect 95970 525835 96018 525891
rect 96074 525835 96122 525891
rect 96178 525835 96226 525891
rect 96282 525835 96330 525891
rect 96386 525835 96434 525891
rect 96490 525835 96538 525891
rect 96594 525835 96642 525891
rect 96698 525835 96746 525891
rect 96802 525835 96850 525891
rect 96906 525835 96954 525891
rect 97010 525835 97058 525891
rect 97114 525835 97162 525891
rect 97218 525835 97266 525891
rect 97322 525835 97370 525891
rect 97426 525835 97474 525891
rect 97530 525835 97578 525891
rect 97634 525835 97682 525891
rect 97738 525835 97786 525891
rect 97842 525835 97890 525891
rect 97946 525835 97994 525891
rect 98050 525835 98098 525891
rect 98154 525835 98202 525891
rect 98258 525835 98306 525891
rect 98362 525835 98410 525891
rect 98466 525835 98514 525891
rect 98570 525835 98618 525891
rect 98674 525835 98722 525891
rect 98778 525835 98826 525891
rect 98882 525835 98930 525891
rect 98986 525835 99034 525891
rect 99090 525835 99138 525891
rect 99194 525835 99242 525891
rect 99298 525835 99346 525891
rect 99402 525835 99450 525891
rect 99506 525835 99554 525891
rect 99610 525835 99658 525891
rect 99714 525835 99762 525891
rect 99818 525835 99866 525891
rect 99922 525835 99970 525891
rect 100026 525835 100074 525891
rect 100130 525835 100178 525891
rect 100234 525835 100282 525891
rect 100338 525835 100386 525891
rect 100442 525835 100490 525891
rect 100546 525835 100594 525891
rect 100650 525835 100698 525891
rect 100754 525835 100802 525891
rect 100858 525835 100906 525891
rect 100962 525835 101010 525891
rect 101066 525835 101114 525891
rect 101170 525835 101218 525891
rect 101274 525835 101322 525891
rect 101378 525835 101426 525891
rect 101482 525835 101530 525891
rect 101586 525835 101634 525891
rect 101690 525835 101738 525891
rect 101794 525835 101842 525891
rect 101898 525835 101946 525891
rect 102002 525835 102050 525891
rect 102106 525835 102154 525891
rect 102210 525835 102258 525891
rect 102314 525835 102362 525891
rect 102418 525835 102466 525891
rect 102522 525835 102570 525891
rect 102626 525835 102674 525891
rect 102730 525835 102778 525891
rect 102834 525835 102882 525891
rect 102938 525835 102986 525891
rect 103042 525835 103090 525891
rect 103146 525835 103194 525891
rect 103250 525835 103298 525891
rect 103354 525835 103402 525891
rect 103458 525835 103506 525891
rect 103562 525835 103610 525891
rect 103666 525835 103714 525891
rect 103770 525835 103818 525891
rect 103874 525835 103922 525891
rect 103978 525835 104026 525891
rect 104082 525835 104130 525891
rect 104186 525835 104234 525891
rect 104290 525835 104338 525891
rect 104394 525835 104442 525891
rect 104498 525835 104546 525891
rect 104602 525835 104650 525891
rect 104706 525835 104754 525891
rect 104810 525835 104858 525891
rect 104914 525835 104962 525891
rect 105018 525835 105066 525891
rect 105122 525835 105170 525891
rect 105226 525835 105274 525891
rect 105330 525835 105378 525891
rect 105434 525835 105482 525891
rect 105538 525835 105586 525891
rect 105642 525835 105690 525891
rect 105746 525835 105794 525891
rect 105850 525835 105898 525891
rect 105954 525835 106002 525891
rect 106058 525835 106106 525891
rect 106162 525835 106210 525891
rect 106266 525835 106314 525891
rect 106370 525835 106418 525891
rect 106474 525835 106522 525891
rect 106578 525835 106626 525891
rect 106682 525835 106730 525891
rect 106786 525835 106834 525891
rect 106890 525835 106938 525891
rect 106994 525835 107042 525891
rect 107098 525835 107146 525891
rect 107202 525835 107250 525891
rect 107306 525835 107354 525891
rect 107410 525835 107458 525891
rect 107514 525835 107562 525891
rect 107618 525835 107666 525891
rect 107722 525835 107770 525891
rect 107826 525835 107874 525891
rect 107930 525835 107978 525891
rect 108034 525835 108082 525891
rect 108138 525835 108186 525891
rect 108242 525835 108290 525891
rect 108346 525835 108394 525891
rect 108450 525835 108498 525891
rect 108554 525835 108602 525891
rect 108658 525835 108706 525891
rect 108762 525835 108810 525891
rect 108866 525835 108900 525891
rect 91200 525826 108900 525835
rect 39858 514294 39954 514350
rect 40010 514294 40078 514350
rect 40134 514294 40202 514350
rect 40258 514294 40326 514350
rect 40382 514294 40478 514350
rect 39858 514226 40478 514294
rect 39858 514170 39954 514226
rect 40010 514170 40078 514226
rect 40134 514170 40202 514226
rect 40258 514170 40326 514226
rect 40382 514170 40478 514226
rect 39858 514102 40478 514170
rect 39858 514046 39954 514102
rect 40010 514046 40078 514102
rect 40134 514046 40202 514102
rect 40258 514046 40326 514102
rect 40382 514046 40478 514102
rect 39858 513978 40478 514046
rect 39858 513922 39954 513978
rect 40010 513922 40078 513978
rect 40134 513922 40202 513978
rect 40258 513922 40326 513978
rect 40382 513922 40478 513978
rect 39858 496350 40478 513922
rect 60300 514412 65550 514446
rect 60300 514356 60355 514412
rect 60411 514356 60479 514412
rect 60535 514356 60603 514412
rect 60659 514356 60727 514412
rect 60783 514356 60851 514412
rect 60907 514356 60975 514412
rect 61031 514356 61099 514412
rect 61155 514356 61223 514412
rect 61279 514356 61347 514412
rect 61403 514356 61471 514412
rect 61527 514356 61595 514412
rect 61651 514356 61719 514412
rect 61775 514356 61843 514412
rect 61899 514356 61967 514412
rect 62023 514356 62091 514412
rect 62147 514356 62215 514412
rect 62271 514356 62339 514412
rect 62395 514356 62463 514412
rect 62519 514356 62587 514412
rect 62643 514356 62711 514412
rect 62767 514356 62835 514412
rect 62891 514356 62959 514412
rect 63015 514356 63083 514412
rect 63139 514356 63207 514412
rect 63263 514356 63331 514412
rect 63387 514356 63455 514412
rect 63511 514356 63579 514412
rect 63635 514356 63703 514412
rect 63759 514356 63827 514412
rect 63883 514356 63951 514412
rect 64007 514356 64075 514412
rect 64131 514356 64199 514412
rect 64255 514356 64323 514412
rect 64379 514356 64447 514412
rect 64503 514356 64571 514412
rect 64627 514356 64695 514412
rect 64751 514356 64819 514412
rect 64875 514356 64943 514412
rect 64999 514356 65067 514412
rect 65123 514356 65191 514412
rect 65247 514356 65315 514412
rect 65371 514356 65439 514412
rect 65495 514356 65550 514412
rect 60300 514288 65550 514356
rect 60300 514232 60355 514288
rect 60411 514232 60479 514288
rect 60535 514232 60603 514288
rect 60659 514232 60727 514288
rect 60783 514232 60851 514288
rect 60907 514232 60975 514288
rect 61031 514232 61099 514288
rect 61155 514232 61223 514288
rect 61279 514232 61347 514288
rect 61403 514232 61471 514288
rect 61527 514232 61595 514288
rect 61651 514232 61719 514288
rect 61775 514232 61843 514288
rect 61899 514232 61967 514288
rect 62023 514232 62091 514288
rect 62147 514232 62215 514288
rect 62271 514232 62339 514288
rect 62395 514232 62463 514288
rect 62519 514232 62587 514288
rect 62643 514232 62711 514288
rect 62767 514232 62835 514288
rect 62891 514232 62959 514288
rect 63015 514232 63083 514288
rect 63139 514232 63207 514288
rect 63263 514232 63331 514288
rect 63387 514232 63455 514288
rect 63511 514232 63579 514288
rect 63635 514232 63703 514288
rect 63759 514232 63827 514288
rect 63883 514232 63951 514288
rect 64007 514232 64075 514288
rect 64131 514232 64199 514288
rect 64255 514232 64323 514288
rect 64379 514232 64447 514288
rect 64503 514232 64571 514288
rect 64627 514232 64695 514288
rect 64751 514232 64819 514288
rect 64875 514232 64943 514288
rect 64999 514232 65067 514288
rect 65123 514232 65191 514288
rect 65247 514232 65315 514288
rect 65371 514232 65439 514288
rect 65495 514232 65550 514288
rect 60300 514164 65550 514232
rect 60300 514108 60355 514164
rect 60411 514108 60479 514164
rect 60535 514108 60603 514164
rect 60659 514108 60727 514164
rect 60783 514108 60851 514164
rect 60907 514108 60975 514164
rect 61031 514108 61099 514164
rect 61155 514108 61223 514164
rect 61279 514108 61347 514164
rect 61403 514108 61471 514164
rect 61527 514108 61595 514164
rect 61651 514108 61719 514164
rect 61775 514108 61843 514164
rect 61899 514108 61967 514164
rect 62023 514108 62091 514164
rect 62147 514108 62215 514164
rect 62271 514108 62339 514164
rect 62395 514108 62463 514164
rect 62519 514108 62587 514164
rect 62643 514108 62711 514164
rect 62767 514108 62835 514164
rect 62891 514108 62959 514164
rect 63015 514108 63083 514164
rect 63139 514108 63207 514164
rect 63263 514108 63331 514164
rect 63387 514108 63455 514164
rect 63511 514108 63579 514164
rect 63635 514108 63703 514164
rect 63759 514108 63827 514164
rect 63883 514108 63951 514164
rect 64007 514108 64075 514164
rect 64131 514108 64199 514164
rect 64255 514108 64323 514164
rect 64379 514108 64447 514164
rect 64503 514108 64571 514164
rect 64627 514108 64695 514164
rect 64751 514108 64819 514164
rect 64875 514108 64943 514164
rect 64999 514108 65067 514164
rect 65123 514108 65191 514164
rect 65247 514108 65315 514164
rect 65371 514108 65439 514164
rect 65495 514108 65550 514164
rect 60300 514040 65550 514108
rect 60300 513984 60355 514040
rect 60411 513984 60479 514040
rect 60535 513984 60603 514040
rect 60659 513984 60727 514040
rect 60783 513984 60851 514040
rect 60907 513984 60975 514040
rect 61031 513984 61099 514040
rect 61155 513984 61223 514040
rect 61279 513984 61347 514040
rect 61403 513984 61471 514040
rect 61527 513984 61595 514040
rect 61651 513984 61719 514040
rect 61775 513984 61843 514040
rect 61899 513984 61967 514040
rect 62023 513984 62091 514040
rect 62147 513984 62215 514040
rect 62271 513984 62339 514040
rect 62395 513984 62463 514040
rect 62519 513984 62587 514040
rect 62643 513984 62711 514040
rect 62767 513984 62835 514040
rect 62891 513984 62959 514040
rect 63015 513984 63083 514040
rect 63139 513984 63207 514040
rect 63263 513984 63331 514040
rect 63387 513984 63455 514040
rect 63511 513984 63579 514040
rect 63635 513984 63703 514040
rect 63759 513984 63827 514040
rect 63883 513984 63951 514040
rect 64007 513984 64075 514040
rect 64131 513984 64199 514040
rect 64255 513984 64323 514040
rect 64379 513984 64447 514040
rect 64503 513984 64571 514040
rect 64627 513984 64695 514040
rect 64751 513984 64819 514040
rect 64875 513984 64943 514040
rect 64999 513984 65067 514040
rect 65123 513984 65191 514040
rect 65247 513984 65315 514040
rect 65371 513984 65439 514040
rect 65495 513984 65550 514040
rect 60300 513916 65550 513984
rect 60300 513860 60355 513916
rect 60411 513860 60479 513916
rect 60535 513860 60603 513916
rect 60659 513860 60727 513916
rect 60783 513860 60851 513916
rect 60907 513860 60975 513916
rect 61031 513860 61099 513916
rect 61155 513860 61223 513916
rect 61279 513860 61347 513916
rect 61403 513860 61471 513916
rect 61527 513860 61595 513916
rect 61651 513860 61719 513916
rect 61775 513860 61843 513916
rect 61899 513860 61967 513916
rect 62023 513860 62091 513916
rect 62147 513860 62215 513916
rect 62271 513860 62339 513916
rect 62395 513860 62463 513916
rect 62519 513860 62587 513916
rect 62643 513860 62711 513916
rect 62767 513860 62835 513916
rect 62891 513860 62959 513916
rect 63015 513860 63083 513916
rect 63139 513860 63207 513916
rect 63263 513860 63331 513916
rect 63387 513860 63455 513916
rect 63511 513860 63579 513916
rect 63635 513860 63703 513916
rect 63759 513860 63827 513916
rect 63883 513860 63951 513916
rect 64007 513860 64075 513916
rect 64131 513860 64199 513916
rect 64255 513860 64323 513916
rect 64379 513860 64447 513916
rect 64503 513860 64571 513916
rect 64627 513860 64695 513916
rect 64751 513860 64819 513916
rect 64875 513860 64943 513916
rect 64999 513860 65067 513916
rect 65123 513860 65191 513916
rect 65247 513860 65315 513916
rect 65371 513860 65439 513916
rect 65495 513860 65550 513916
rect 60300 513826 65550 513860
rect 159018 508350 159638 525922
rect 85200 508290 85318 508350
rect 85200 508234 85231 508290
rect 85287 508234 85318 508290
rect 85200 508166 85318 508234
rect 85200 508110 85231 508166
rect 85287 508110 85318 508166
rect 85200 508050 85318 508110
rect 85324 508290 85814 508350
rect 85324 508234 85355 508290
rect 85411 508234 85479 508290
rect 85535 508234 85603 508290
rect 85659 508234 85727 508290
rect 85783 508234 85814 508290
rect 85324 508166 85814 508234
rect 85324 508110 85355 508166
rect 85411 508110 85479 508166
rect 85535 508110 85603 508166
rect 85659 508110 85727 508166
rect 85783 508110 85814 508166
rect 85324 508050 85814 508110
rect 85820 508290 86310 508350
rect 85820 508234 85851 508290
rect 85907 508234 85975 508290
rect 86031 508234 86099 508290
rect 86155 508234 86223 508290
rect 86279 508234 86310 508290
rect 85820 508166 86310 508234
rect 85820 508110 85851 508166
rect 85907 508110 85975 508166
rect 86031 508110 86099 508166
rect 86155 508110 86223 508166
rect 86279 508110 86310 508166
rect 85820 508050 86310 508110
rect 86316 508290 86806 508350
rect 86316 508234 86347 508290
rect 86403 508234 86471 508290
rect 86527 508234 86595 508290
rect 86651 508234 86719 508290
rect 86775 508234 86806 508290
rect 86316 508166 86806 508234
rect 86316 508110 86347 508166
rect 86403 508110 86471 508166
rect 86527 508110 86595 508166
rect 86651 508110 86719 508166
rect 86775 508110 86806 508166
rect 86316 508050 86806 508110
rect 86812 508290 87302 508350
rect 86812 508234 86843 508290
rect 86899 508234 86967 508290
rect 87023 508234 87091 508290
rect 87147 508234 87215 508290
rect 87271 508234 87302 508290
rect 86812 508166 87302 508234
rect 86812 508110 86843 508166
rect 86899 508110 86967 508166
rect 87023 508110 87091 508166
rect 87147 508110 87215 508166
rect 87271 508110 87302 508166
rect 86812 508050 87302 508110
rect 87308 508290 87798 508350
rect 87308 508234 87339 508290
rect 87395 508234 87463 508290
rect 87519 508234 87587 508290
rect 87643 508234 87711 508290
rect 87767 508234 87798 508290
rect 87308 508166 87798 508234
rect 87308 508110 87339 508166
rect 87395 508110 87463 508166
rect 87519 508110 87587 508166
rect 87643 508110 87711 508166
rect 87767 508110 87798 508166
rect 87308 508050 87798 508110
rect 87804 508290 88294 508350
rect 87804 508234 87835 508290
rect 87891 508234 87959 508290
rect 88015 508234 88083 508290
rect 88139 508234 88207 508290
rect 88263 508234 88294 508290
rect 87804 508166 88294 508234
rect 87804 508110 87835 508166
rect 87891 508110 87959 508166
rect 88015 508110 88083 508166
rect 88139 508110 88207 508166
rect 88263 508110 88294 508166
rect 87804 508050 88294 508110
rect 88300 508290 88790 508350
rect 88300 508234 88331 508290
rect 88387 508234 88455 508290
rect 88511 508234 88579 508290
rect 88635 508234 88703 508290
rect 88759 508234 88790 508290
rect 88300 508166 88790 508234
rect 88300 508110 88331 508166
rect 88387 508110 88455 508166
rect 88511 508110 88579 508166
rect 88635 508110 88703 508166
rect 88759 508110 88790 508166
rect 88300 508050 88790 508110
rect 88796 508290 89286 508350
rect 88796 508234 88827 508290
rect 88883 508234 88951 508290
rect 89007 508234 89075 508290
rect 89131 508234 89199 508290
rect 89255 508234 89286 508290
rect 88796 508166 89286 508234
rect 88796 508110 88827 508166
rect 88883 508110 88951 508166
rect 89007 508110 89075 508166
rect 89131 508110 89199 508166
rect 89255 508110 89286 508166
rect 88796 508050 89286 508110
rect 89292 508290 89782 508350
rect 89292 508234 89323 508290
rect 89379 508234 89447 508290
rect 89503 508234 89571 508290
rect 89627 508234 89695 508290
rect 89751 508234 89782 508290
rect 89292 508166 89782 508234
rect 89292 508110 89323 508166
rect 89379 508110 89447 508166
rect 89503 508110 89571 508166
rect 89627 508110 89695 508166
rect 89751 508110 89782 508166
rect 89292 508050 89782 508110
rect 89788 508290 90278 508350
rect 89788 508234 89819 508290
rect 89875 508234 89943 508290
rect 89999 508234 90067 508290
rect 90123 508234 90191 508290
rect 90247 508234 90278 508290
rect 89788 508166 90278 508234
rect 89788 508110 89819 508166
rect 89875 508110 89943 508166
rect 89999 508110 90067 508166
rect 90123 508110 90191 508166
rect 90247 508110 90278 508166
rect 89788 508050 90278 508110
rect 90284 508290 90774 508350
rect 90284 508234 90315 508290
rect 90371 508234 90439 508290
rect 90495 508234 90563 508290
rect 90619 508234 90687 508290
rect 90743 508234 90774 508290
rect 90284 508166 90774 508234
rect 90284 508110 90315 508166
rect 90371 508110 90439 508166
rect 90495 508110 90563 508166
rect 90619 508110 90687 508166
rect 90743 508110 90774 508166
rect 90284 508050 90774 508110
rect 90780 508290 91270 508350
rect 90780 508234 90811 508290
rect 90867 508234 90935 508290
rect 90991 508234 91059 508290
rect 91115 508234 91183 508290
rect 91239 508234 91270 508290
rect 90780 508166 91270 508234
rect 90780 508110 90811 508166
rect 90867 508110 90935 508166
rect 90991 508110 91059 508166
rect 91115 508110 91183 508166
rect 91239 508110 91270 508166
rect 90780 508050 91270 508110
rect 91276 508290 91766 508350
rect 91276 508234 91307 508290
rect 91363 508234 91431 508290
rect 91487 508234 91555 508290
rect 91611 508234 91679 508290
rect 91735 508234 91766 508290
rect 91276 508166 91766 508234
rect 91276 508110 91307 508166
rect 91363 508110 91431 508166
rect 91487 508110 91555 508166
rect 91611 508110 91679 508166
rect 91735 508110 91766 508166
rect 91276 508050 91766 508110
rect 91772 508290 92262 508350
rect 91772 508234 91803 508290
rect 91859 508234 91927 508290
rect 91983 508234 92051 508290
rect 92107 508234 92175 508290
rect 92231 508234 92262 508290
rect 91772 508166 92262 508234
rect 91772 508110 91803 508166
rect 91859 508110 91927 508166
rect 91983 508110 92051 508166
rect 92107 508110 92175 508166
rect 92231 508110 92262 508166
rect 91772 508050 92262 508110
rect 92268 508290 92758 508350
rect 92268 508234 92299 508290
rect 92355 508234 92423 508290
rect 92479 508234 92547 508290
rect 92603 508234 92671 508290
rect 92727 508234 92758 508290
rect 92268 508166 92758 508234
rect 92268 508110 92299 508166
rect 92355 508110 92423 508166
rect 92479 508110 92547 508166
rect 92603 508110 92671 508166
rect 92727 508110 92758 508166
rect 92268 508050 92758 508110
rect 92764 508290 93254 508350
rect 92764 508234 92795 508290
rect 92851 508234 92919 508290
rect 92975 508234 93043 508290
rect 93099 508234 93167 508290
rect 93223 508234 93254 508290
rect 92764 508166 93254 508234
rect 92764 508110 92795 508166
rect 92851 508110 92919 508166
rect 92975 508110 93043 508166
rect 93099 508110 93167 508166
rect 93223 508110 93254 508166
rect 92764 508050 93254 508110
rect 93260 508290 93750 508350
rect 93260 508234 93291 508290
rect 93347 508234 93415 508290
rect 93471 508234 93539 508290
rect 93595 508234 93663 508290
rect 93719 508234 93750 508290
rect 93260 508166 93750 508234
rect 93260 508110 93291 508166
rect 93347 508110 93415 508166
rect 93471 508110 93539 508166
rect 93595 508110 93663 508166
rect 93719 508110 93750 508166
rect 93260 508050 93750 508110
rect 159018 508294 159114 508350
rect 159170 508294 159238 508350
rect 159294 508294 159362 508350
rect 159418 508294 159486 508350
rect 159542 508294 159638 508350
rect 159018 508226 159638 508294
rect 159018 508170 159114 508226
rect 159170 508170 159238 508226
rect 159294 508170 159362 508226
rect 159418 508170 159486 508226
rect 159542 508170 159638 508226
rect 159018 508102 159638 508170
rect 159018 508046 159114 508102
rect 159170 508046 159238 508102
rect 159294 508046 159362 508102
rect 159418 508046 159486 508102
rect 159542 508046 159638 508102
rect 159018 507978 159638 508046
rect 159018 507922 159114 507978
rect 159170 507922 159238 507978
rect 159294 507922 159362 507978
rect 159418 507922 159486 507978
rect 159542 507922 159638 507978
rect 85050 507891 93450 507900
rect 85050 507835 85062 507891
rect 85118 507835 85166 507891
rect 85222 507835 85270 507891
rect 85326 507835 85374 507891
rect 85430 507835 85478 507891
rect 85534 507835 85582 507891
rect 85638 507835 85686 507891
rect 85742 507835 85790 507891
rect 85846 507835 85894 507891
rect 85950 507835 85998 507891
rect 86054 507835 86102 507891
rect 86158 507835 86206 507891
rect 86262 507835 86310 507891
rect 86366 507835 86414 507891
rect 86470 507835 86518 507891
rect 86574 507835 86622 507891
rect 86678 507835 86726 507891
rect 86782 507835 86830 507891
rect 86886 507835 86934 507891
rect 86990 507835 87038 507891
rect 87094 507835 87142 507891
rect 87198 507835 87246 507891
rect 87302 507835 87350 507891
rect 87406 507835 87454 507891
rect 87510 507835 87558 507891
rect 87614 507835 87662 507891
rect 87718 507835 87766 507891
rect 87822 507835 87870 507891
rect 87926 507835 87974 507891
rect 88030 507835 88078 507891
rect 88134 507835 88182 507891
rect 88238 507835 88286 507891
rect 88342 507835 88390 507891
rect 88446 507835 88494 507891
rect 88550 507835 88598 507891
rect 88654 507835 88702 507891
rect 88758 507835 88806 507891
rect 88862 507835 88910 507891
rect 88966 507835 89014 507891
rect 89070 507835 89118 507891
rect 89174 507835 89222 507891
rect 89278 507835 89326 507891
rect 89382 507835 89430 507891
rect 89486 507835 89534 507891
rect 89590 507835 89638 507891
rect 89694 507835 89742 507891
rect 89798 507835 89846 507891
rect 89902 507835 89950 507891
rect 90006 507835 90054 507891
rect 90110 507835 90158 507891
rect 90214 507835 90262 507891
rect 90318 507835 90366 507891
rect 90422 507835 90470 507891
rect 90526 507835 90574 507891
rect 90630 507835 90678 507891
rect 90734 507835 90782 507891
rect 90838 507835 90886 507891
rect 90942 507835 90990 507891
rect 91046 507835 91094 507891
rect 91150 507835 91198 507891
rect 91254 507835 91302 507891
rect 91358 507835 91406 507891
rect 91462 507835 91510 507891
rect 91566 507835 91614 507891
rect 91670 507835 91718 507891
rect 91774 507835 91822 507891
rect 91878 507835 91926 507891
rect 91982 507835 92030 507891
rect 92086 507835 92134 507891
rect 92190 507835 92238 507891
rect 92294 507835 92342 507891
rect 92398 507835 92446 507891
rect 92502 507835 92550 507891
rect 92606 507835 92654 507891
rect 92710 507835 92758 507891
rect 92814 507835 92862 507891
rect 92918 507835 92966 507891
rect 93022 507835 93070 507891
rect 93126 507835 93174 507891
rect 93230 507835 93278 507891
rect 93334 507835 93382 507891
rect 93438 507835 93450 507891
rect 85050 507826 93450 507835
rect 39858 496294 39954 496350
rect 40010 496294 40078 496350
rect 40134 496294 40202 496350
rect 40258 496294 40326 496350
rect 40382 496294 40478 496350
rect 39858 496226 40478 496294
rect 39858 496170 39954 496226
rect 40010 496170 40078 496226
rect 40134 496170 40202 496226
rect 40258 496170 40326 496226
rect 40382 496170 40478 496226
rect 39858 496102 40478 496170
rect 39858 496046 39954 496102
rect 40010 496046 40078 496102
rect 40134 496046 40202 496102
rect 40258 496046 40326 496102
rect 40382 496046 40478 496102
rect 39858 495978 40478 496046
rect 39858 495922 39954 495978
rect 40010 495922 40078 495978
rect 40134 495922 40202 495978
rect 40258 495922 40326 495978
rect 40382 495922 40478 495978
rect 39858 478350 40478 495922
rect 39858 478294 39954 478350
rect 40010 478294 40078 478350
rect 40134 478294 40202 478350
rect 40258 478294 40326 478350
rect 40382 478294 40478 478350
rect 39858 478226 40478 478294
rect 39858 478170 39954 478226
rect 40010 478170 40078 478226
rect 40134 478170 40202 478226
rect 40258 478170 40326 478226
rect 40382 478170 40478 478226
rect 39858 478102 40478 478170
rect 39858 478046 39954 478102
rect 40010 478046 40078 478102
rect 40134 478046 40202 478102
rect 40258 478046 40326 478102
rect 40382 478046 40478 478102
rect 39858 477978 40478 478046
rect 39858 477922 39954 477978
rect 40010 477922 40078 477978
rect 40134 477922 40202 477978
rect 40258 477922 40326 477978
rect 40382 477922 40478 477978
rect 39858 460350 40478 477922
rect 39858 460294 39954 460350
rect 40010 460294 40078 460350
rect 40134 460294 40202 460350
rect 40258 460294 40326 460350
rect 40382 460294 40478 460350
rect 39858 460226 40478 460294
rect 39858 460170 39954 460226
rect 40010 460170 40078 460226
rect 40134 460170 40202 460226
rect 40258 460170 40326 460226
rect 40382 460170 40478 460226
rect 39858 460102 40478 460170
rect 39858 460046 39954 460102
rect 40010 460046 40078 460102
rect 40134 460046 40202 460102
rect 40258 460046 40326 460102
rect 40382 460046 40478 460102
rect 39858 459978 40478 460046
rect 39858 459922 39954 459978
rect 40010 459922 40078 459978
rect 40134 459922 40202 459978
rect 40258 459922 40326 459978
rect 40382 459922 40478 459978
rect 39858 442350 40478 459922
rect 39858 442294 39954 442350
rect 40010 442294 40078 442350
rect 40134 442294 40202 442350
rect 40258 442294 40326 442350
rect 40382 442294 40478 442350
rect 39858 442226 40478 442294
rect 39858 442170 39954 442226
rect 40010 442170 40078 442226
rect 40134 442170 40202 442226
rect 40258 442170 40326 442226
rect 40382 442170 40478 442226
rect 39858 442102 40478 442170
rect 39858 442046 39954 442102
rect 40010 442046 40078 442102
rect 40134 442046 40202 442102
rect 40258 442046 40326 442102
rect 40382 442046 40478 442102
rect 39858 441978 40478 442046
rect 39858 441922 39954 441978
rect 40010 441922 40078 441978
rect 40134 441922 40202 441978
rect 40258 441922 40326 441978
rect 40382 441922 40478 441978
rect 39858 424350 40478 441922
rect 39858 424294 39954 424350
rect 40010 424294 40078 424350
rect 40134 424294 40202 424350
rect 40258 424294 40326 424350
rect 40382 424294 40478 424350
rect 39858 424226 40478 424294
rect 39858 424170 39954 424226
rect 40010 424170 40078 424226
rect 40134 424170 40202 424226
rect 40258 424170 40326 424226
rect 40382 424170 40478 424226
rect 39858 424102 40478 424170
rect 39858 424046 39954 424102
rect 40010 424046 40078 424102
rect 40134 424046 40202 424102
rect 40258 424046 40326 424102
rect 40382 424046 40478 424102
rect 39858 423978 40478 424046
rect 39858 423922 39954 423978
rect 40010 423922 40078 423978
rect 40134 423922 40202 423978
rect 40258 423922 40326 423978
rect 40382 423922 40478 423978
rect 39858 406350 40478 423922
rect 57932 502516 57988 502526
rect 57932 409258 57988 502460
rect 63450 496413 69450 496446
rect 63450 496357 63508 496413
rect 63564 496357 63632 496413
rect 63688 496357 63756 496413
rect 63812 496357 63880 496413
rect 63936 496357 64004 496413
rect 64060 496357 64128 496413
rect 64184 496357 64252 496413
rect 64308 496357 64376 496413
rect 64432 496357 64500 496413
rect 64556 496357 64624 496413
rect 64680 496357 64748 496413
rect 64804 496357 64872 496413
rect 64928 496357 64996 496413
rect 65052 496357 65120 496413
rect 65176 496357 65244 496413
rect 65300 496357 65368 496413
rect 65424 496357 65492 496413
rect 65548 496357 65616 496413
rect 65672 496357 65740 496413
rect 65796 496357 65864 496413
rect 65920 496357 65988 496413
rect 66044 496357 66112 496413
rect 66168 496357 66236 496413
rect 66292 496357 66360 496413
rect 66416 496357 66484 496413
rect 66540 496357 66608 496413
rect 66664 496357 66732 496413
rect 66788 496357 66856 496413
rect 66912 496357 66980 496413
rect 67036 496357 67104 496413
rect 67160 496357 67228 496413
rect 67284 496357 67352 496413
rect 67408 496357 67476 496413
rect 67532 496357 67600 496413
rect 67656 496357 67724 496413
rect 67780 496357 67848 496413
rect 67904 496357 67972 496413
rect 68028 496357 68096 496413
rect 68152 496357 68220 496413
rect 68276 496357 68344 496413
rect 68400 496357 68468 496413
rect 68524 496357 68592 496413
rect 68648 496357 68716 496413
rect 68772 496357 68840 496413
rect 68896 496357 68964 496413
rect 69020 496357 69088 496413
rect 69144 496357 69212 496413
rect 69268 496357 69336 496413
rect 69392 496357 69450 496413
rect 63450 496289 69450 496357
rect 63450 496233 63508 496289
rect 63564 496233 63632 496289
rect 63688 496233 63756 496289
rect 63812 496233 63880 496289
rect 63936 496233 64004 496289
rect 64060 496233 64128 496289
rect 64184 496233 64252 496289
rect 64308 496233 64376 496289
rect 64432 496233 64500 496289
rect 64556 496233 64624 496289
rect 64680 496233 64748 496289
rect 64804 496233 64872 496289
rect 64928 496233 64996 496289
rect 65052 496233 65120 496289
rect 65176 496233 65244 496289
rect 65300 496233 65368 496289
rect 65424 496233 65492 496289
rect 65548 496233 65616 496289
rect 65672 496233 65740 496289
rect 65796 496233 65864 496289
rect 65920 496233 65988 496289
rect 66044 496233 66112 496289
rect 66168 496233 66236 496289
rect 66292 496233 66360 496289
rect 66416 496233 66484 496289
rect 66540 496233 66608 496289
rect 66664 496233 66732 496289
rect 66788 496233 66856 496289
rect 66912 496233 66980 496289
rect 67036 496233 67104 496289
rect 67160 496233 67228 496289
rect 67284 496233 67352 496289
rect 67408 496233 67476 496289
rect 67532 496233 67600 496289
rect 67656 496233 67724 496289
rect 67780 496233 67848 496289
rect 67904 496233 67972 496289
rect 68028 496233 68096 496289
rect 68152 496233 68220 496289
rect 68276 496233 68344 496289
rect 68400 496233 68468 496289
rect 68524 496233 68592 496289
rect 68648 496233 68716 496289
rect 68772 496233 68840 496289
rect 68896 496233 68964 496289
rect 69020 496233 69088 496289
rect 69144 496233 69212 496289
rect 69268 496233 69336 496289
rect 69392 496233 69450 496289
rect 63450 496200 69450 496233
rect 63600 496003 69750 496050
rect 63600 495947 63671 496003
rect 63727 495947 63795 496003
rect 63851 495947 63919 496003
rect 63975 495947 64043 496003
rect 64099 495947 64167 496003
rect 64223 495947 64291 496003
rect 64347 495947 64415 496003
rect 64471 495947 64539 496003
rect 64595 495947 64663 496003
rect 64719 495947 64787 496003
rect 64843 495947 64911 496003
rect 64967 495947 65035 496003
rect 65091 495947 65159 496003
rect 65215 495947 65283 496003
rect 65339 495947 65407 496003
rect 65463 495947 65531 496003
rect 65587 495947 65655 496003
rect 65711 495947 65779 496003
rect 65835 495947 65903 496003
rect 65959 495947 66027 496003
rect 66083 495947 66151 496003
rect 66207 495947 66275 496003
rect 66331 495947 66399 496003
rect 66455 495947 66523 496003
rect 66579 495947 66647 496003
rect 66703 495947 66771 496003
rect 66827 495947 66895 496003
rect 66951 495947 67019 496003
rect 67075 495947 67143 496003
rect 67199 495947 67267 496003
rect 67323 495947 67391 496003
rect 67447 495947 67515 496003
rect 67571 495947 67639 496003
rect 67695 495947 67763 496003
rect 67819 495947 67887 496003
rect 67943 495947 68011 496003
rect 68067 495947 68135 496003
rect 68191 495947 68259 496003
rect 68315 495947 68383 496003
rect 68439 495947 68507 496003
rect 68563 495947 68631 496003
rect 68687 495947 68755 496003
rect 68811 495947 68879 496003
rect 68935 495947 69003 496003
rect 69059 495947 69127 496003
rect 69183 495947 69251 496003
rect 69307 495947 69375 496003
rect 69431 495947 69499 496003
rect 69555 495947 69623 496003
rect 69679 495947 69750 496003
rect 63600 495900 69750 495947
rect 128298 490350 128918 497538
rect 80550 490290 82800 490350
rect 80550 490234 80593 490290
rect 80649 490234 80717 490290
rect 80773 490234 80841 490290
rect 80897 490234 80965 490290
rect 81021 490234 81089 490290
rect 81145 490234 81213 490290
rect 81269 490234 81337 490290
rect 81393 490234 81461 490290
rect 81517 490234 81585 490290
rect 81641 490234 81709 490290
rect 81765 490234 81833 490290
rect 81889 490234 81957 490290
rect 82013 490234 82081 490290
rect 82137 490234 82205 490290
rect 82261 490234 82329 490290
rect 82385 490234 82453 490290
rect 82509 490234 82577 490290
rect 82633 490234 82701 490290
rect 82757 490234 82800 490290
rect 80550 490166 82800 490234
rect 80550 490110 80593 490166
rect 80649 490110 80717 490166
rect 80773 490110 80841 490166
rect 80897 490110 80965 490166
rect 81021 490110 81089 490166
rect 81145 490110 81213 490166
rect 81269 490110 81337 490166
rect 81393 490110 81461 490166
rect 81517 490110 81585 490166
rect 81641 490110 81709 490166
rect 81765 490110 81833 490166
rect 81889 490110 81957 490166
rect 82013 490110 82081 490166
rect 82137 490110 82205 490166
rect 82261 490110 82329 490166
rect 82385 490110 82453 490166
rect 82509 490110 82577 490166
rect 82633 490110 82701 490166
rect 82757 490110 82800 490166
rect 80550 490050 82800 490110
rect 128298 490294 128394 490350
rect 128450 490294 128518 490350
rect 128574 490294 128642 490350
rect 128698 490294 128766 490350
rect 128822 490294 128918 490350
rect 128298 490226 128918 490294
rect 128298 490170 128394 490226
rect 128450 490170 128518 490226
rect 128574 490170 128642 490226
rect 128698 490170 128766 490226
rect 128822 490170 128918 490226
rect 128298 490102 128918 490170
rect 128298 490046 128394 490102
rect 128450 490046 128518 490102
rect 128574 490046 128642 490102
rect 128698 490046 128766 490102
rect 128822 490046 128918 490102
rect 128298 489978 128918 490046
rect 128298 489922 128394 489978
rect 128450 489922 128518 489978
rect 128574 489922 128642 489978
rect 128698 489922 128766 489978
rect 128822 489922 128918 489978
rect 80400 489891 82650 489900
rect 80400 489835 80457 489891
rect 80513 489835 80561 489891
rect 80617 489835 80665 489891
rect 80721 489835 80769 489891
rect 80825 489835 80873 489891
rect 80929 489835 80977 489891
rect 81033 489835 81081 489891
rect 81137 489835 81185 489891
rect 81241 489835 81289 489891
rect 81345 489835 81393 489891
rect 81449 489835 81497 489891
rect 81553 489835 81601 489891
rect 81657 489835 81705 489891
rect 81761 489835 81809 489891
rect 81865 489835 81913 489891
rect 81969 489835 82017 489891
rect 82073 489835 82121 489891
rect 82177 489835 82225 489891
rect 82281 489835 82329 489891
rect 82385 489835 82433 489891
rect 82489 489835 82537 489891
rect 82593 489835 82650 489891
rect 80400 489826 82650 489835
rect 57932 409192 57988 409202
rect 66858 472350 67478 488238
rect 66858 472294 66954 472350
rect 67010 472294 67078 472350
rect 67134 472294 67202 472350
rect 67258 472294 67326 472350
rect 67382 472294 67478 472350
rect 66858 472226 67478 472294
rect 66858 472170 66954 472226
rect 67010 472170 67078 472226
rect 67134 472170 67202 472226
rect 67258 472170 67326 472226
rect 67382 472170 67478 472226
rect 66858 472102 67478 472170
rect 66858 472046 66954 472102
rect 67010 472046 67078 472102
rect 67134 472046 67202 472102
rect 67258 472046 67326 472102
rect 67382 472046 67478 472102
rect 66858 471978 67478 472046
rect 66858 471922 66954 471978
rect 67010 471922 67078 471978
rect 67134 471922 67202 471978
rect 67258 471922 67326 471978
rect 67382 471922 67478 471978
rect 66858 454350 67478 471922
rect 66858 454294 66954 454350
rect 67010 454294 67078 454350
rect 67134 454294 67202 454350
rect 67258 454294 67326 454350
rect 67382 454294 67478 454350
rect 66858 454226 67478 454294
rect 66858 454170 66954 454226
rect 67010 454170 67078 454226
rect 67134 454170 67202 454226
rect 67258 454170 67326 454226
rect 67382 454170 67478 454226
rect 66858 454102 67478 454170
rect 66858 454046 66954 454102
rect 67010 454046 67078 454102
rect 67134 454046 67202 454102
rect 67258 454046 67326 454102
rect 67382 454046 67478 454102
rect 66858 453978 67478 454046
rect 66858 453922 66954 453978
rect 67010 453922 67078 453978
rect 67134 453922 67202 453978
rect 67258 453922 67326 453978
rect 67382 453922 67478 453978
rect 66858 436350 67478 453922
rect 66858 436294 66954 436350
rect 67010 436294 67078 436350
rect 67134 436294 67202 436350
rect 67258 436294 67326 436350
rect 67382 436294 67478 436350
rect 66858 436226 67478 436294
rect 66858 436170 66954 436226
rect 67010 436170 67078 436226
rect 67134 436170 67202 436226
rect 67258 436170 67326 436226
rect 67382 436170 67478 436226
rect 66858 436102 67478 436170
rect 66858 436046 66954 436102
rect 67010 436046 67078 436102
rect 67134 436046 67202 436102
rect 67258 436046 67326 436102
rect 67382 436046 67478 436102
rect 66858 435978 67478 436046
rect 66858 435922 66954 435978
rect 67010 435922 67078 435978
rect 67134 435922 67202 435978
rect 67258 435922 67326 435978
rect 67382 435922 67478 435978
rect 66858 418350 67478 435922
rect 66858 418294 66954 418350
rect 67010 418294 67078 418350
rect 67134 418294 67202 418350
rect 67258 418294 67326 418350
rect 67382 418294 67478 418350
rect 66858 418226 67478 418294
rect 66858 418170 66954 418226
rect 67010 418170 67078 418226
rect 67134 418170 67202 418226
rect 67258 418170 67326 418226
rect 67382 418170 67478 418226
rect 66858 418102 67478 418170
rect 66858 418046 66954 418102
rect 67010 418046 67078 418102
rect 67134 418046 67202 418102
rect 67258 418046 67326 418102
rect 67382 418046 67478 418102
rect 66858 417978 67478 418046
rect 66858 417922 66954 417978
rect 67010 417922 67078 417978
rect 67134 417922 67202 417978
rect 67258 417922 67326 417978
rect 67382 417922 67478 417978
rect 39858 406294 39954 406350
rect 40010 406294 40078 406350
rect 40134 406294 40202 406350
rect 40258 406294 40326 406350
rect 40382 406294 40478 406350
rect 39858 406226 40478 406294
rect 39858 406170 39954 406226
rect 40010 406170 40078 406226
rect 40134 406170 40202 406226
rect 40258 406170 40326 406226
rect 40382 406170 40478 406226
rect 39858 406102 40478 406170
rect 39858 406046 39954 406102
rect 40010 406046 40078 406102
rect 40134 406046 40202 406102
rect 40258 406046 40326 406102
rect 40382 406046 40478 406102
rect 39858 405978 40478 406046
rect 39858 405922 39954 405978
rect 40010 405922 40078 405978
rect 40134 405922 40202 405978
rect 40258 405922 40326 405978
rect 40382 405922 40478 405978
rect 39858 388350 40478 405922
rect 39858 388294 39954 388350
rect 40010 388294 40078 388350
rect 40134 388294 40202 388350
rect 40258 388294 40326 388350
rect 40382 388294 40478 388350
rect 39858 388226 40478 388294
rect 39858 388170 39954 388226
rect 40010 388170 40078 388226
rect 40134 388170 40202 388226
rect 40258 388170 40326 388226
rect 40382 388170 40478 388226
rect 39858 388102 40478 388170
rect 39858 388046 39954 388102
rect 40010 388046 40078 388102
rect 40134 388046 40202 388102
rect 40258 388046 40326 388102
rect 40382 388046 40478 388102
rect 39858 387978 40478 388046
rect 39858 387922 39954 387978
rect 40010 387922 40078 387978
rect 40134 387922 40202 387978
rect 40258 387922 40326 387978
rect 40382 387922 40478 387978
rect 39858 370350 40478 387922
rect 39858 370294 39954 370350
rect 40010 370294 40078 370350
rect 40134 370294 40202 370350
rect 40258 370294 40326 370350
rect 40382 370294 40478 370350
rect 39858 370226 40478 370294
rect 39858 370170 39954 370226
rect 40010 370170 40078 370226
rect 40134 370170 40202 370226
rect 40258 370170 40326 370226
rect 40382 370170 40478 370226
rect 39858 370102 40478 370170
rect 39858 370046 39954 370102
rect 40010 370046 40078 370102
rect 40134 370046 40202 370102
rect 40258 370046 40326 370102
rect 40382 370046 40478 370102
rect 39858 369978 40478 370046
rect 39858 369922 39954 369978
rect 40010 369922 40078 369978
rect 40134 369922 40202 369978
rect 40258 369922 40326 369978
rect 40382 369922 40478 369978
rect 39858 352350 40478 369922
rect 39858 352294 39954 352350
rect 40010 352294 40078 352350
rect 40134 352294 40202 352350
rect 40258 352294 40326 352350
rect 40382 352294 40478 352350
rect 39858 352226 40478 352294
rect 39858 352170 39954 352226
rect 40010 352170 40078 352226
rect 40134 352170 40202 352226
rect 40258 352170 40326 352226
rect 40382 352170 40478 352226
rect 39858 352102 40478 352170
rect 39858 352046 39954 352102
rect 40010 352046 40078 352102
rect 40134 352046 40202 352102
rect 40258 352046 40326 352102
rect 40382 352046 40478 352102
rect 39858 351978 40478 352046
rect 39858 351922 39954 351978
rect 40010 351922 40078 351978
rect 40134 351922 40202 351978
rect 40258 351922 40326 351978
rect 40382 351922 40478 351978
rect 39858 334350 40478 351922
rect 39858 334294 39954 334350
rect 40010 334294 40078 334350
rect 40134 334294 40202 334350
rect 40258 334294 40326 334350
rect 40382 334294 40478 334350
rect 39858 334226 40478 334294
rect 39858 334170 39954 334226
rect 40010 334170 40078 334226
rect 40134 334170 40202 334226
rect 40258 334170 40326 334226
rect 40382 334170 40478 334226
rect 39858 334102 40478 334170
rect 39858 334046 39954 334102
rect 40010 334046 40078 334102
rect 40134 334046 40202 334102
rect 40258 334046 40326 334102
rect 40382 334046 40478 334102
rect 39858 333978 40478 334046
rect 39858 333922 39954 333978
rect 40010 333922 40078 333978
rect 40134 333922 40202 333978
rect 40258 333922 40326 333978
rect 40382 333922 40478 333978
rect 39858 316350 40478 333922
rect 39858 316294 39954 316350
rect 40010 316294 40078 316350
rect 40134 316294 40202 316350
rect 40258 316294 40326 316350
rect 40382 316294 40478 316350
rect 39858 316226 40478 316294
rect 39858 316170 39954 316226
rect 40010 316170 40078 316226
rect 40134 316170 40202 316226
rect 40258 316170 40326 316226
rect 40382 316170 40478 316226
rect 39858 316102 40478 316170
rect 39858 316046 39954 316102
rect 40010 316046 40078 316102
rect 40134 316046 40202 316102
rect 40258 316046 40326 316102
rect 40382 316046 40478 316102
rect 39858 315978 40478 316046
rect 39858 315922 39954 315978
rect 40010 315922 40078 315978
rect 40134 315922 40202 315978
rect 40258 315922 40326 315978
rect 40382 315922 40478 315978
rect 39858 298350 40478 315922
rect 66858 400350 67478 417922
rect 66858 400294 66954 400350
rect 67010 400294 67078 400350
rect 67134 400294 67202 400350
rect 67258 400294 67326 400350
rect 67382 400294 67478 400350
rect 66858 400226 67478 400294
rect 66858 400170 66954 400226
rect 67010 400170 67078 400226
rect 67134 400170 67202 400226
rect 67258 400170 67326 400226
rect 67382 400170 67478 400226
rect 66858 400102 67478 400170
rect 66858 400046 66954 400102
rect 67010 400046 67078 400102
rect 67134 400046 67202 400102
rect 67258 400046 67326 400102
rect 67382 400046 67478 400102
rect 66858 399978 67478 400046
rect 66858 399922 66954 399978
rect 67010 399922 67078 399978
rect 67134 399922 67202 399978
rect 67258 399922 67326 399978
rect 67382 399922 67478 399978
rect 66858 382350 67478 399922
rect 66858 382294 66954 382350
rect 67010 382294 67078 382350
rect 67134 382294 67202 382350
rect 67258 382294 67326 382350
rect 67382 382294 67478 382350
rect 66858 382226 67478 382294
rect 66858 382170 66954 382226
rect 67010 382170 67078 382226
rect 67134 382170 67202 382226
rect 67258 382170 67326 382226
rect 67382 382170 67478 382226
rect 66858 382102 67478 382170
rect 66858 382046 66954 382102
rect 67010 382046 67078 382102
rect 67134 382046 67202 382102
rect 67258 382046 67326 382102
rect 67382 382046 67478 382102
rect 66858 381978 67478 382046
rect 66858 381922 66954 381978
rect 67010 381922 67078 381978
rect 67134 381922 67202 381978
rect 67258 381922 67326 381978
rect 67382 381922 67478 381978
rect 66858 364350 67478 381922
rect 66858 364294 66954 364350
rect 67010 364294 67078 364350
rect 67134 364294 67202 364350
rect 67258 364294 67326 364350
rect 67382 364294 67478 364350
rect 66858 364226 67478 364294
rect 66858 364170 66954 364226
rect 67010 364170 67078 364226
rect 67134 364170 67202 364226
rect 67258 364170 67326 364226
rect 67382 364170 67478 364226
rect 66858 364102 67478 364170
rect 66858 364046 66954 364102
rect 67010 364046 67078 364102
rect 67134 364046 67202 364102
rect 67258 364046 67326 364102
rect 67382 364046 67478 364102
rect 66858 363978 67478 364046
rect 66858 363922 66954 363978
rect 67010 363922 67078 363978
rect 67134 363922 67202 363978
rect 67258 363922 67326 363978
rect 67382 363922 67478 363978
rect 66858 346350 67478 363922
rect 66858 346294 66954 346350
rect 67010 346294 67078 346350
rect 67134 346294 67202 346350
rect 67258 346294 67326 346350
rect 67382 346294 67478 346350
rect 66858 346226 67478 346294
rect 66858 346170 66954 346226
rect 67010 346170 67078 346226
rect 67134 346170 67202 346226
rect 67258 346170 67326 346226
rect 67382 346170 67478 346226
rect 66858 346102 67478 346170
rect 66858 346046 66954 346102
rect 67010 346046 67078 346102
rect 67134 346046 67202 346102
rect 67258 346046 67326 346102
rect 67382 346046 67478 346102
rect 66858 345978 67478 346046
rect 66858 345922 66954 345978
rect 67010 345922 67078 345978
rect 67134 345922 67202 345978
rect 67258 345922 67326 345978
rect 67382 345922 67478 345978
rect 66858 328350 67478 345922
rect 66858 328294 66954 328350
rect 67010 328294 67078 328350
rect 67134 328294 67202 328350
rect 67258 328294 67326 328350
rect 67382 328294 67478 328350
rect 66858 328226 67478 328294
rect 66858 328170 66954 328226
rect 67010 328170 67078 328226
rect 67134 328170 67202 328226
rect 67258 328170 67326 328226
rect 67382 328170 67478 328226
rect 66858 328102 67478 328170
rect 66858 328046 66954 328102
rect 67010 328046 67078 328102
rect 67134 328046 67202 328102
rect 67258 328046 67326 328102
rect 67382 328046 67478 328102
rect 66858 327978 67478 328046
rect 66858 327922 66954 327978
rect 67010 327922 67078 327978
rect 67134 327922 67202 327978
rect 67258 327922 67326 327978
rect 67382 327922 67478 327978
rect 66858 310350 67478 327922
rect 66858 310294 66954 310350
rect 67010 310294 67078 310350
rect 67134 310294 67202 310350
rect 67258 310294 67326 310350
rect 67382 310294 67478 310350
rect 66858 310226 67478 310294
rect 66858 310170 66954 310226
rect 67010 310170 67078 310226
rect 67134 310170 67202 310226
rect 67258 310170 67326 310226
rect 67382 310170 67478 310226
rect 66858 310102 67478 310170
rect 66858 310046 66954 310102
rect 67010 310046 67078 310102
rect 67134 310046 67202 310102
rect 67258 310046 67326 310102
rect 67382 310046 67478 310102
rect 66858 309978 67478 310046
rect 66858 309922 66954 309978
rect 67010 309922 67078 309978
rect 67134 309922 67202 309978
rect 67258 309922 67326 309978
rect 67382 309922 67478 309978
rect 39858 298294 39954 298350
rect 40010 298294 40078 298350
rect 40134 298294 40202 298350
rect 40258 298294 40326 298350
rect 40382 298294 40478 298350
rect 39858 298226 40478 298294
rect 39858 298170 39954 298226
rect 40010 298170 40078 298226
rect 40134 298170 40202 298226
rect 40258 298170 40326 298226
rect 40382 298170 40478 298226
rect 39858 298102 40478 298170
rect 39858 298046 39954 298102
rect 40010 298046 40078 298102
rect 40134 298046 40202 298102
rect 40258 298046 40326 298102
rect 40382 298046 40478 298102
rect 39858 297978 40478 298046
rect 39858 297922 39954 297978
rect 40010 297922 40078 297978
rect 40134 297922 40202 297978
rect 40258 297922 40326 297978
rect 40382 297922 40478 297978
rect 39858 280350 40478 297922
rect 47404 299348 47460 299358
rect 47404 297444 47460 299292
rect 66858 298094 67478 309922
rect 70578 478350 71198 484638
rect 70578 478294 70674 478350
rect 70730 478294 70798 478350
rect 70854 478294 70922 478350
rect 70978 478294 71046 478350
rect 71102 478294 71198 478350
rect 101298 478350 101918 479238
rect 70578 478226 71198 478294
rect 70578 478170 70674 478226
rect 70730 478170 70798 478226
rect 70854 478170 70922 478226
rect 70978 478170 71046 478226
rect 71102 478170 71198 478226
rect 70578 478102 71198 478170
rect 70578 478046 70674 478102
rect 70730 478046 70798 478102
rect 70854 478046 70922 478102
rect 70978 478046 71046 478102
rect 71102 478046 71198 478102
rect 70578 477978 71198 478046
rect 70578 477922 70674 477978
rect 70730 477922 70798 477978
rect 70854 477922 70922 477978
rect 70978 477922 71046 477978
rect 71102 477922 71198 477978
rect 70578 460350 71198 477922
rect 70578 460294 70674 460350
rect 70730 460294 70798 460350
rect 70854 460294 70922 460350
rect 70978 460294 71046 460350
rect 71102 460294 71198 460350
rect 70578 460226 71198 460294
rect 70578 460170 70674 460226
rect 70730 460170 70798 460226
rect 70854 460170 70922 460226
rect 70978 460170 71046 460226
rect 71102 460170 71198 460226
rect 70578 460102 71198 460170
rect 70578 460046 70674 460102
rect 70730 460046 70798 460102
rect 70854 460046 70922 460102
rect 70978 460046 71046 460102
rect 71102 460046 71198 460102
rect 70578 459978 71198 460046
rect 70578 459922 70674 459978
rect 70730 459922 70798 459978
rect 70854 459922 70922 459978
rect 70978 459922 71046 459978
rect 71102 459922 71198 459978
rect 70578 442350 71198 459922
rect 70578 442294 70674 442350
rect 70730 442294 70798 442350
rect 70854 442294 70922 442350
rect 70978 442294 71046 442350
rect 71102 442294 71198 442350
rect 70578 442226 71198 442294
rect 70578 442170 70674 442226
rect 70730 442170 70798 442226
rect 70854 442170 70922 442226
rect 70978 442170 71046 442226
rect 71102 442170 71198 442226
rect 70578 442102 71198 442170
rect 70578 442046 70674 442102
rect 70730 442046 70798 442102
rect 70854 442046 70922 442102
rect 70978 442046 71046 442102
rect 71102 442046 71198 442102
rect 70578 441978 71198 442046
rect 70578 441922 70674 441978
rect 70730 441922 70798 441978
rect 70854 441922 70922 441978
rect 70978 441922 71046 441978
rect 71102 441922 71198 441978
rect 70578 424350 71198 441922
rect 70578 424294 70674 424350
rect 70730 424294 70798 424350
rect 70854 424294 70922 424350
rect 70978 424294 71046 424350
rect 71102 424294 71198 424350
rect 70578 424226 71198 424294
rect 70578 424170 70674 424226
rect 70730 424170 70798 424226
rect 70854 424170 70922 424226
rect 70978 424170 71046 424226
rect 71102 424170 71198 424226
rect 70578 424102 71198 424170
rect 70578 424046 70674 424102
rect 70730 424046 70798 424102
rect 70854 424046 70922 424102
rect 70978 424046 71046 424102
rect 71102 424046 71198 424102
rect 70578 423978 71198 424046
rect 70578 423922 70674 423978
rect 70730 423922 70798 423978
rect 70854 423922 70922 423978
rect 70978 423922 71046 423978
rect 71102 423922 71198 423978
rect 70578 406350 71198 423922
rect 70578 406294 70674 406350
rect 70730 406294 70798 406350
rect 70854 406294 70922 406350
rect 70978 406294 71046 406350
rect 71102 406294 71198 406350
rect 70578 406226 71198 406294
rect 70578 406170 70674 406226
rect 70730 406170 70798 406226
rect 70854 406170 70922 406226
rect 70978 406170 71046 406226
rect 71102 406170 71198 406226
rect 70578 406102 71198 406170
rect 70578 406046 70674 406102
rect 70730 406046 70798 406102
rect 70854 406046 70922 406102
rect 70978 406046 71046 406102
rect 71102 406046 71198 406102
rect 70578 405978 71198 406046
rect 70578 405922 70674 405978
rect 70730 405922 70798 405978
rect 70854 405922 70922 405978
rect 70978 405922 71046 405978
rect 71102 405922 71198 405978
rect 70578 388350 71198 405922
rect 70578 388294 70674 388350
rect 70730 388294 70798 388350
rect 70854 388294 70922 388350
rect 70978 388294 71046 388350
rect 71102 388294 71198 388350
rect 70578 388226 71198 388294
rect 70578 388170 70674 388226
rect 70730 388170 70798 388226
rect 70854 388170 70922 388226
rect 70978 388170 71046 388226
rect 71102 388170 71198 388226
rect 70578 388102 71198 388170
rect 70578 388046 70674 388102
rect 70730 388046 70798 388102
rect 70854 388046 70922 388102
rect 70978 388046 71046 388102
rect 71102 388046 71198 388102
rect 70578 387978 71198 388046
rect 70578 387922 70674 387978
rect 70730 387922 70798 387978
rect 70854 387922 70922 387978
rect 70978 387922 71046 387978
rect 71102 387922 71198 387978
rect 70578 370350 71198 387922
rect 70578 370294 70674 370350
rect 70730 370294 70798 370350
rect 70854 370294 70922 370350
rect 70978 370294 71046 370350
rect 71102 370294 71198 370350
rect 70578 370226 71198 370294
rect 70578 370170 70674 370226
rect 70730 370170 70798 370226
rect 70854 370170 70922 370226
rect 70978 370170 71046 370226
rect 71102 370170 71198 370226
rect 70578 370102 71198 370170
rect 70578 370046 70674 370102
rect 70730 370046 70798 370102
rect 70854 370046 70922 370102
rect 70978 370046 71046 370102
rect 71102 370046 71198 370102
rect 70578 369978 71198 370046
rect 70578 369922 70674 369978
rect 70730 369922 70798 369978
rect 70854 369922 70922 369978
rect 70978 369922 71046 369978
rect 71102 369922 71198 369978
rect 70578 352350 71198 369922
rect 70578 352294 70674 352350
rect 70730 352294 70798 352350
rect 70854 352294 70922 352350
rect 70978 352294 71046 352350
rect 71102 352294 71198 352350
rect 70578 352226 71198 352294
rect 70578 352170 70674 352226
rect 70730 352170 70798 352226
rect 70854 352170 70922 352226
rect 70978 352170 71046 352226
rect 71102 352170 71198 352226
rect 70578 352102 71198 352170
rect 70578 352046 70674 352102
rect 70730 352046 70798 352102
rect 70854 352046 70922 352102
rect 70978 352046 71046 352102
rect 71102 352046 71198 352102
rect 70578 351978 71198 352046
rect 70578 351922 70674 351978
rect 70730 351922 70798 351978
rect 70854 351922 70922 351978
rect 70978 351922 71046 351978
rect 71102 351922 71198 351978
rect 70578 334350 71198 351922
rect 70578 334294 70674 334350
rect 70730 334294 70798 334350
rect 70854 334294 70922 334350
rect 70978 334294 71046 334350
rect 71102 334294 71198 334350
rect 70578 334226 71198 334294
rect 70578 334170 70674 334226
rect 70730 334170 70798 334226
rect 70854 334170 70922 334226
rect 70978 334170 71046 334226
rect 71102 334170 71198 334226
rect 70578 334102 71198 334170
rect 70578 334046 70674 334102
rect 70730 334046 70798 334102
rect 70854 334046 70922 334102
rect 70978 334046 71046 334102
rect 71102 334046 71198 334102
rect 70578 333978 71198 334046
rect 70578 333922 70674 333978
rect 70730 333922 70798 333978
rect 70854 333922 70922 333978
rect 70978 333922 71046 333978
rect 71102 333922 71198 333978
rect 70578 316350 71198 333922
rect 70578 316294 70674 316350
rect 70730 316294 70798 316350
rect 70854 316294 70922 316350
rect 70978 316294 71046 316350
rect 71102 316294 71198 316350
rect 70578 316226 71198 316294
rect 70578 316170 70674 316226
rect 70730 316170 70798 316226
rect 70854 316170 70922 316226
rect 70978 316170 71046 316226
rect 71102 316170 71198 316226
rect 70578 316102 71198 316170
rect 70578 316046 70674 316102
rect 70730 316046 70798 316102
rect 70854 316046 70922 316102
rect 70978 316046 71046 316102
rect 71102 316046 71198 316102
rect 70578 315978 71198 316046
rect 70578 315922 70674 315978
rect 70730 315922 70798 315978
rect 70854 315922 70922 315978
rect 70978 315922 71046 315978
rect 71102 315922 71198 315978
rect 70578 298422 71198 315922
rect 70578 298366 70674 298422
rect 70730 298366 70798 298422
rect 70854 298366 70922 298422
rect 70978 298366 71046 298422
rect 71102 298366 71198 298422
rect 70578 298298 71198 298366
rect 70578 298242 70674 298298
rect 70730 298242 70798 298298
rect 70854 298242 70922 298298
rect 70978 298242 71046 298298
rect 71102 298242 71198 298298
rect 70578 298174 71198 298242
rect 70578 298118 70674 298174
rect 70730 298118 70798 298174
rect 70854 298118 70922 298174
rect 70978 298118 71046 298174
rect 71102 298118 71198 298174
rect 70578 298094 71198 298118
rect 97578 472350 98198 478338
rect 97578 472294 97674 472350
rect 97730 472294 97798 472350
rect 97854 472294 97922 472350
rect 97978 472294 98046 472350
rect 98102 472294 98198 472350
rect 97578 472226 98198 472294
rect 97578 472170 97674 472226
rect 97730 472170 97798 472226
rect 97854 472170 97922 472226
rect 97978 472170 98046 472226
rect 98102 472170 98198 472226
rect 97578 472102 98198 472170
rect 97578 472046 97674 472102
rect 97730 472046 97798 472102
rect 97854 472046 97922 472102
rect 97978 472046 98046 472102
rect 98102 472046 98198 472102
rect 97578 471978 98198 472046
rect 97578 471922 97674 471978
rect 97730 471922 97798 471978
rect 97854 471922 97922 471978
rect 97978 471922 98046 471978
rect 98102 471922 98198 471978
rect 97578 454350 98198 471922
rect 97578 454294 97674 454350
rect 97730 454294 97798 454350
rect 97854 454294 97922 454350
rect 97978 454294 98046 454350
rect 98102 454294 98198 454350
rect 97578 454226 98198 454294
rect 97578 454170 97674 454226
rect 97730 454170 97798 454226
rect 97854 454170 97922 454226
rect 97978 454170 98046 454226
rect 98102 454170 98198 454226
rect 97578 454102 98198 454170
rect 97578 454046 97674 454102
rect 97730 454046 97798 454102
rect 97854 454046 97922 454102
rect 97978 454046 98046 454102
rect 98102 454046 98198 454102
rect 97578 453978 98198 454046
rect 97578 453922 97674 453978
rect 97730 453922 97798 453978
rect 97854 453922 97922 453978
rect 97978 453922 98046 453978
rect 98102 453922 98198 453978
rect 97578 436350 98198 453922
rect 97578 436294 97674 436350
rect 97730 436294 97798 436350
rect 97854 436294 97922 436350
rect 97978 436294 98046 436350
rect 98102 436294 98198 436350
rect 97578 436226 98198 436294
rect 97578 436170 97674 436226
rect 97730 436170 97798 436226
rect 97854 436170 97922 436226
rect 97978 436170 98046 436226
rect 98102 436170 98198 436226
rect 97578 436102 98198 436170
rect 97578 436046 97674 436102
rect 97730 436046 97798 436102
rect 97854 436046 97922 436102
rect 97978 436046 98046 436102
rect 98102 436046 98198 436102
rect 97578 435978 98198 436046
rect 97578 435922 97674 435978
rect 97730 435922 97798 435978
rect 97854 435922 97922 435978
rect 97978 435922 98046 435978
rect 98102 435922 98198 435978
rect 97578 418350 98198 435922
rect 97578 418294 97674 418350
rect 97730 418294 97798 418350
rect 97854 418294 97922 418350
rect 97978 418294 98046 418350
rect 98102 418294 98198 418350
rect 97578 418226 98198 418294
rect 97578 418170 97674 418226
rect 97730 418170 97798 418226
rect 97854 418170 97922 418226
rect 97978 418170 98046 418226
rect 98102 418170 98198 418226
rect 97578 418102 98198 418170
rect 97578 418046 97674 418102
rect 97730 418046 97798 418102
rect 97854 418046 97922 418102
rect 97978 418046 98046 418102
rect 98102 418046 98198 418102
rect 97578 417978 98198 418046
rect 97578 417922 97674 417978
rect 97730 417922 97798 417978
rect 97854 417922 97922 417978
rect 97978 417922 98046 417978
rect 98102 417922 98198 417978
rect 97578 400350 98198 417922
rect 97578 400294 97674 400350
rect 97730 400294 97798 400350
rect 97854 400294 97922 400350
rect 97978 400294 98046 400350
rect 98102 400294 98198 400350
rect 97578 400226 98198 400294
rect 97578 400170 97674 400226
rect 97730 400170 97798 400226
rect 97854 400170 97922 400226
rect 97978 400170 98046 400226
rect 98102 400170 98198 400226
rect 97578 400102 98198 400170
rect 97578 400046 97674 400102
rect 97730 400046 97798 400102
rect 97854 400046 97922 400102
rect 97978 400046 98046 400102
rect 98102 400046 98198 400102
rect 97578 399978 98198 400046
rect 97578 399922 97674 399978
rect 97730 399922 97798 399978
rect 97854 399922 97922 399978
rect 97978 399922 98046 399978
rect 98102 399922 98198 399978
rect 97578 382350 98198 399922
rect 101298 478294 101394 478350
rect 101450 478294 101518 478350
rect 101574 478294 101642 478350
rect 101698 478294 101766 478350
rect 101822 478294 101918 478350
rect 101298 478226 101918 478294
rect 101298 478170 101394 478226
rect 101450 478170 101518 478226
rect 101574 478170 101642 478226
rect 101698 478170 101766 478226
rect 101822 478170 101918 478226
rect 101298 478102 101918 478170
rect 101298 478046 101394 478102
rect 101450 478046 101518 478102
rect 101574 478046 101642 478102
rect 101698 478046 101766 478102
rect 101822 478046 101918 478102
rect 101298 477978 101918 478046
rect 101298 477922 101394 477978
rect 101450 477922 101518 477978
rect 101574 477922 101642 477978
rect 101698 477922 101766 477978
rect 101822 477922 101918 477978
rect 101298 460350 101918 477922
rect 101298 460294 101394 460350
rect 101450 460294 101518 460350
rect 101574 460294 101642 460350
rect 101698 460294 101766 460350
rect 101822 460294 101918 460350
rect 101298 460226 101918 460294
rect 101298 460170 101394 460226
rect 101450 460170 101518 460226
rect 101574 460170 101642 460226
rect 101698 460170 101766 460226
rect 101822 460170 101918 460226
rect 101298 460102 101918 460170
rect 101298 460046 101394 460102
rect 101450 460046 101518 460102
rect 101574 460046 101642 460102
rect 101698 460046 101766 460102
rect 101822 460046 101918 460102
rect 101298 459978 101918 460046
rect 101298 459922 101394 459978
rect 101450 459922 101518 459978
rect 101574 459922 101642 459978
rect 101698 459922 101766 459978
rect 101822 459922 101918 459978
rect 101298 442350 101918 459922
rect 101298 442294 101394 442350
rect 101450 442294 101518 442350
rect 101574 442294 101642 442350
rect 101698 442294 101766 442350
rect 101822 442294 101918 442350
rect 101298 442226 101918 442294
rect 101298 442170 101394 442226
rect 101450 442170 101518 442226
rect 101574 442170 101642 442226
rect 101698 442170 101766 442226
rect 101822 442170 101918 442226
rect 101298 442102 101918 442170
rect 101298 442046 101394 442102
rect 101450 442046 101518 442102
rect 101574 442046 101642 442102
rect 101698 442046 101766 442102
rect 101822 442046 101918 442102
rect 101298 441978 101918 442046
rect 101298 441922 101394 441978
rect 101450 441922 101518 441978
rect 101574 441922 101642 441978
rect 101698 441922 101766 441978
rect 101822 441922 101918 441978
rect 101298 424350 101918 441922
rect 101298 424294 101394 424350
rect 101450 424294 101518 424350
rect 101574 424294 101642 424350
rect 101698 424294 101766 424350
rect 101822 424294 101918 424350
rect 101298 424226 101918 424294
rect 101298 424170 101394 424226
rect 101450 424170 101518 424226
rect 101574 424170 101642 424226
rect 101698 424170 101766 424226
rect 101822 424170 101918 424226
rect 101298 424102 101918 424170
rect 101298 424046 101394 424102
rect 101450 424046 101518 424102
rect 101574 424046 101642 424102
rect 101698 424046 101766 424102
rect 101822 424046 101918 424102
rect 101298 423978 101918 424046
rect 101298 423922 101394 423978
rect 101450 423922 101518 423978
rect 101574 423922 101642 423978
rect 101698 423922 101766 423978
rect 101822 423922 101918 423978
rect 101298 406350 101918 423922
rect 101298 406294 101394 406350
rect 101450 406294 101518 406350
rect 101574 406294 101642 406350
rect 101698 406294 101766 406350
rect 101822 406294 101918 406350
rect 101298 406226 101918 406294
rect 101298 406170 101394 406226
rect 101450 406170 101518 406226
rect 101574 406170 101642 406226
rect 101698 406170 101766 406226
rect 101822 406170 101918 406226
rect 101298 406102 101918 406170
rect 101298 406046 101394 406102
rect 101450 406046 101518 406102
rect 101574 406046 101642 406102
rect 101698 406046 101766 406102
rect 101822 406046 101918 406102
rect 101298 405978 101918 406046
rect 101298 405922 101394 405978
rect 101450 405922 101518 405978
rect 101574 405922 101642 405978
rect 101698 405922 101766 405978
rect 101822 405922 101918 405978
rect 101298 388350 101918 405922
rect 128298 472350 128918 489922
rect 128298 472294 128394 472350
rect 128450 472294 128518 472350
rect 128574 472294 128642 472350
rect 128698 472294 128766 472350
rect 128822 472294 128918 472350
rect 128298 472226 128918 472294
rect 128298 472170 128394 472226
rect 128450 472170 128518 472226
rect 128574 472170 128642 472226
rect 128698 472170 128766 472226
rect 128822 472170 128918 472226
rect 128298 472102 128918 472170
rect 128298 472046 128394 472102
rect 128450 472046 128518 472102
rect 128574 472046 128642 472102
rect 128698 472046 128766 472102
rect 128822 472046 128918 472102
rect 128298 471978 128918 472046
rect 128298 471922 128394 471978
rect 128450 471922 128518 471978
rect 128574 471922 128642 471978
rect 128698 471922 128766 471978
rect 128822 471922 128918 471978
rect 128298 454350 128918 471922
rect 128298 454294 128394 454350
rect 128450 454294 128518 454350
rect 128574 454294 128642 454350
rect 128698 454294 128766 454350
rect 128822 454294 128918 454350
rect 128298 454226 128918 454294
rect 128298 454170 128394 454226
rect 128450 454170 128518 454226
rect 128574 454170 128642 454226
rect 128698 454170 128766 454226
rect 128822 454170 128918 454226
rect 128298 454102 128918 454170
rect 128298 454046 128394 454102
rect 128450 454046 128518 454102
rect 128574 454046 128642 454102
rect 128698 454046 128766 454102
rect 128822 454046 128918 454102
rect 128298 453978 128918 454046
rect 128298 453922 128394 453978
rect 128450 453922 128518 453978
rect 128574 453922 128642 453978
rect 128698 453922 128766 453978
rect 128822 453922 128918 453978
rect 128298 436350 128918 453922
rect 128298 436294 128394 436350
rect 128450 436294 128518 436350
rect 128574 436294 128642 436350
rect 128698 436294 128766 436350
rect 128822 436294 128918 436350
rect 128298 436226 128918 436294
rect 128298 436170 128394 436226
rect 128450 436170 128518 436226
rect 128574 436170 128642 436226
rect 128698 436170 128766 436226
rect 128822 436170 128918 436226
rect 128298 436102 128918 436170
rect 128298 436046 128394 436102
rect 128450 436046 128518 436102
rect 128574 436046 128642 436102
rect 128698 436046 128766 436102
rect 128822 436046 128918 436102
rect 128298 435978 128918 436046
rect 128298 435922 128394 435978
rect 128450 435922 128518 435978
rect 128574 435922 128642 435978
rect 128698 435922 128766 435978
rect 128822 435922 128918 435978
rect 128298 418350 128918 435922
rect 128298 418294 128394 418350
rect 128450 418294 128518 418350
rect 128574 418294 128642 418350
rect 128698 418294 128766 418350
rect 128822 418294 128918 418350
rect 128298 418226 128918 418294
rect 128298 418170 128394 418226
rect 128450 418170 128518 418226
rect 128574 418170 128642 418226
rect 128698 418170 128766 418226
rect 128822 418170 128918 418226
rect 128298 418102 128918 418170
rect 128298 418046 128394 418102
rect 128450 418046 128518 418102
rect 128574 418046 128642 418102
rect 128698 418046 128766 418102
rect 128822 418046 128918 418102
rect 128298 417978 128918 418046
rect 128298 417922 128394 417978
rect 128450 417922 128518 417978
rect 128574 417922 128642 417978
rect 128698 417922 128766 417978
rect 128822 417922 128918 417978
rect 128298 400350 128918 417922
rect 128298 400294 128394 400350
rect 128450 400294 128518 400350
rect 128574 400294 128642 400350
rect 128698 400294 128766 400350
rect 128822 400294 128918 400350
rect 128298 400226 128918 400294
rect 128298 400170 128394 400226
rect 128450 400170 128518 400226
rect 128574 400170 128642 400226
rect 128698 400170 128766 400226
rect 128822 400170 128918 400226
rect 128298 400102 128918 400170
rect 128298 400046 128394 400102
rect 128450 400046 128518 400102
rect 128574 400046 128642 400102
rect 128698 400046 128766 400102
rect 128822 400046 128918 400102
rect 128298 399978 128918 400046
rect 128298 399922 128394 399978
rect 128450 399922 128518 399978
rect 128574 399922 128642 399978
rect 128698 399922 128766 399978
rect 128822 399922 128918 399978
rect 101298 388294 101394 388350
rect 101450 388294 101518 388350
rect 101574 388294 101642 388350
rect 101698 388294 101766 388350
rect 101822 388294 101918 388350
rect 101298 388226 101918 388294
rect 101298 388170 101394 388226
rect 101450 388170 101518 388226
rect 101574 388170 101642 388226
rect 101698 388170 101766 388226
rect 101822 388170 101918 388226
rect 101298 388102 101918 388170
rect 101298 388046 101394 388102
rect 101450 388046 101518 388102
rect 101574 388046 101642 388102
rect 101698 388046 101766 388102
rect 101822 388046 101918 388102
rect 101298 387978 101918 388046
rect 101298 387922 101394 387978
rect 101450 387922 101518 387978
rect 101574 387922 101642 387978
rect 101698 387922 101766 387978
rect 101822 387922 101918 387978
rect 97578 382294 97674 382350
rect 97730 382294 97798 382350
rect 97854 382294 97922 382350
rect 97978 382294 98046 382350
rect 98102 382294 98198 382350
rect 97578 382226 98198 382294
rect 97578 382170 97674 382226
rect 97730 382170 97798 382226
rect 97854 382170 97922 382226
rect 97978 382170 98046 382226
rect 98102 382170 98198 382226
rect 97578 382102 98198 382170
rect 97578 382046 97674 382102
rect 97730 382046 97798 382102
rect 97854 382046 97922 382102
rect 97978 382046 98046 382102
rect 98102 382046 98198 382102
rect 97578 381978 98198 382046
rect 97578 381922 97674 381978
rect 97730 381922 97798 381978
rect 97854 381922 97922 381978
rect 97978 381922 98046 381978
rect 98102 381922 98198 381978
rect 97578 364350 98198 381922
rect 97578 364294 97674 364350
rect 97730 364294 97798 364350
rect 97854 364294 97922 364350
rect 97978 364294 98046 364350
rect 98102 364294 98198 364350
rect 97578 364226 98198 364294
rect 97578 364170 97674 364226
rect 97730 364170 97798 364226
rect 97854 364170 97922 364226
rect 97978 364170 98046 364226
rect 98102 364170 98198 364226
rect 97578 364102 98198 364170
rect 97578 364046 97674 364102
rect 97730 364046 97798 364102
rect 97854 364046 97922 364102
rect 97978 364046 98046 364102
rect 98102 364046 98198 364102
rect 97578 363978 98198 364046
rect 97578 363922 97674 363978
rect 97730 363922 97798 363978
rect 97854 363922 97922 363978
rect 97978 363922 98046 363978
rect 98102 363922 98198 363978
rect 97578 346350 98198 363922
rect 97578 346294 97674 346350
rect 97730 346294 97798 346350
rect 97854 346294 97922 346350
rect 97978 346294 98046 346350
rect 98102 346294 98198 346350
rect 97578 346226 98198 346294
rect 97578 346170 97674 346226
rect 97730 346170 97798 346226
rect 97854 346170 97922 346226
rect 97978 346170 98046 346226
rect 98102 346170 98198 346226
rect 97578 346102 98198 346170
rect 97578 346046 97674 346102
rect 97730 346046 97798 346102
rect 97854 346046 97922 346102
rect 97978 346046 98046 346102
rect 98102 346046 98198 346102
rect 97578 345978 98198 346046
rect 97578 345922 97674 345978
rect 97730 345922 97798 345978
rect 97854 345922 97922 345978
rect 97978 345922 98046 345978
rect 98102 345922 98198 345978
rect 97578 328350 98198 345922
rect 97578 328294 97674 328350
rect 97730 328294 97798 328350
rect 97854 328294 97922 328350
rect 97978 328294 98046 328350
rect 98102 328294 98198 328350
rect 97578 328226 98198 328294
rect 97578 328170 97674 328226
rect 97730 328170 97798 328226
rect 97854 328170 97922 328226
rect 97978 328170 98046 328226
rect 98102 328170 98198 328226
rect 97578 328102 98198 328170
rect 97578 328046 97674 328102
rect 97730 328046 97798 328102
rect 97854 328046 97922 328102
rect 97978 328046 98046 328102
rect 98102 328046 98198 328102
rect 97578 327978 98198 328046
rect 97578 327922 97674 327978
rect 97730 327922 97798 327978
rect 97854 327922 97922 327978
rect 97978 327922 98046 327978
rect 98102 327922 98198 327978
rect 97578 310350 98198 327922
rect 97578 310294 97674 310350
rect 97730 310294 97798 310350
rect 97854 310294 97922 310350
rect 97978 310294 98046 310350
rect 98102 310294 98198 310350
rect 97578 310226 98198 310294
rect 97578 310170 97674 310226
rect 97730 310170 97798 310226
rect 97854 310170 97922 310226
rect 97978 310170 98046 310226
rect 98102 310170 98198 310226
rect 97578 310102 98198 310170
rect 97578 310046 97674 310102
rect 97730 310046 97798 310102
rect 97854 310046 97922 310102
rect 97978 310046 98046 310102
rect 98102 310046 98198 310102
rect 97578 309978 98198 310046
rect 97578 309922 97674 309978
rect 97730 309922 97798 309978
rect 97854 309922 97922 309978
rect 97978 309922 98046 309978
rect 98102 309922 98198 309978
rect 47404 297378 47460 297388
rect 48524 297444 48580 297454
rect 44448 292350 44768 292384
rect 44448 292294 44518 292350
rect 44574 292294 44642 292350
rect 44698 292294 44768 292350
rect 44448 292226 44768 292294
rect 44448 292170 44518 292226
rect 44574 292170 44642 292226
rect 44698 292170 44768 292226
rect 44448 292102 44768 292170
rect 44448 292046 44518 292102
rect 44574 292046 44642 292102
rect 44698 292046 44768 292102
rect 44448 291978 44768 292046
rect 44448 291922 44518 291978
rect 44574 291922 44642 291978
rect 44698 291922 44768 291978
rect 44448 291888 44768 291922
rect 39858 280294 39954 280350
rect 40010 280294 40078 280350
rect 40134 280294 40202 280350
rect 40258 280294 40326 280350
rect 40382 280294 40478 280350
rect 39858 280226 40478 280294
rect 39858 280170 39954 280226
rect 40010 280170 40078 280226
rect 40134 280170 40202 280226
rect 40258 280170 40326 280226
rect 40382 280170 40478 280226
rect 39858 280102 40478 280170
rect 39858 280046 39954 280102
rect 40010 280046 40078 280102
rect 40134 280046 40202 280102
rect 40258 280046 40326 280102
rect 40382 280046 40478 280102
rect 39858 279978 40478 280046
rect 39858 279922 39954 279978
rect 40010 279922 40078 279978
rect 40134 279922 40202 279978
rect 40258 279922 40326 279978
rect 40382 279922 40478 279978
rect 39858 262350 40478 279922
rect 44448 274350 44768 274384
rect 44448 274294 44518 274350
rect 44574 274294 44642 274350
rect 44698 274294 44768 274350
rect 44448 274226 44768 274294
rect 44448 274170 44518 274226
rect 44574 274170 44642 274226
rect 44698 274170 44768 274226
rect 44448 274102 44768 274170
rect 44448 274046 44518 274102
rect 44574 274046 44642 274102
rect 44698 274046 44768 274102
rect 44448 273978 44768 274046
rect 44448 273922 44518 273978
rect 44574 273922 44642 273978
rect 44698 273922 44768 273978
rect 44448 273888 44768 273922
rect 39858 262294 39954 262350
rect 40010 262294 40078 262350
rect 40134 262294 40202 262350
rect 40258 262294 40326 262350
rect 40382 262294 40478 262350
rect 39858 262226 40478 262294
rect 39858 262170 39954 262226
rect 40010 262170 40078 262226
rect 40134 262170 40202 262226
rect 40258 262170 40326 262226
rect 40382 262170 40478 262226
rect 39858 262102 40478 262170
rect 39858 262046 39954 262102
rect 40010 262046 40078 262102
rect 40134 262046 40202 262102
rect 40258 262046 40326 262102
rect 40382 262046 40478 262102
rect 39858 261978 40478 262046
rect 39858 261922 39954 261978
rect 40010 261922 40078 261978
rect 40134 261922 40202 261978
rect 40258 261922 40326 261978
rect 40382 261922 40478 261978
rect 39858 244350 40478 261922
rect 44448 256350 44768 256384
rect 44448 256294 44518 256350
rect 44574 256294 44642 256350
rect 44698 256294 44768 256350
rect 44448 256226 44768 256294
rect 44448 256170 44518 256226
rect 44574 256170 44642 256226
rect 44698 256170 44768 256226
rect 44448 256102 44768 256170
rect 44448 256046 44518 256102
rect 44574 256046 44642 256102
rect 44698 256046 44768 256102
rect 44448 255978 44768 256046
rect 44448 255922 44518 255978
rect 44574 255922 44642 255978
rect 44698 255922 44768 255978
rect 44448 255888 44768 255922
rect 39858 244294 39954 244350
rect 40010 244294 40078 244350
rect 40134 244294 40202 244350
rect 40258 244294 40326 244350
rect 40382 244294 40478 244350
rect 39858 244226 40478 244294
rect 39858 244170 39954 244226
rect 40010 244170 40078 244226
rect 40134 244170 40202 244226
rect 40258 244170 40326 244226
rect 40382 244170 40478 244226
rect 39858 244102 40478 244170
rect 39858 244046 39954 244102
rect 40010 244046 40078 244102
rect 40134 244046 40202 244102
rect 40258 244046 40326 244102
rect 40382 244046 40478 244102
rect 39858 243978 40478 244046
rect 39858 243922 39954 243978
rect 40010 243922 40078 243978
rect 40134 243922 40202 243978
rect 40258 243922 40326 243978
rect 40382 243922 40478 243978
rect 39858 226350 40478 243922
rect 46172 247078 46228 247088
rect 46172 242564 46228 247022
rect 46172 242498 46228 242508
rect 39858 226294 39954 226350
rect 40010 226294 40078 226350
rect 40134 226294 40202 226350
rect 40258 226294 40326 226350
rect 40382 226294 40478 226350
rect 39858 226226 40478 226294
rect 39858 226170 39954 226226
rect 40010 226170 40078 226226
rect 40134 226170 40202 226226
rect 40258 226170 40326 226226
rect 40382 226170 40478 226226
rect 39858 226102 40478 226170
rect 39858 226046 39954 226102
rect 40010 226046 40078 226102
rect 40134 226046 40202 226102
rect 40258 226046 40326 226102
rect 40382 226046 40478 226102
rect 39858 225978 40478 226046
rect 39858 225922 39954 225978
rect 40010 225922 40078 225978
rect 40134 225922 40202 225978
rect 40258 225922 40326 225978
rect 40382 225922 40478 225978
rect 39858 208350 40478 225922
rect 39858 208294 39954 208350
rect 40010 208294 40078 208350
rect 40134 208294 40202 208350
rect 40258 208294 40326 208350
rect 40382 208294 40478 208350
rect 39858 208226 40478 208294
rect 39858 208170 39954 208226
rect 40010 208170 40078 208226
rect 40134 208170 40202 208226
rect 40258 208170 40326 208226
rect 40382 208170 40478 208226
rect 39858 208102 40478 208170
rect 39858 208046 39954 208102
rect 40010 208046 40078 208102
rect 40134 208046 40202 208102
rect 40258 208046 40326 208102
rect 40382 208046 40478 208102
rect 39858 207978 40478 208046
rect 39858 207922 39954 207978
rect 40010 207922 40078 207978
rect 40134 207922 40202 207978
rect 40258 207922 40326 207978
rect 40382 207922 40478 207978
rect 39858 190350 40478 207922
rect 44448 202350 44768 202384
rect 44448 202294 44518 202350
rect 44574 202294 44642 202350
rect 44698 202294 44768 202350
rect 44448 202226 44768 202294
rect 44448 202170 44518 202226
rect 44574 202170 44642 202226
rect 44698 202170 44768 202226
rect 44448 202102 44768 202170
rect 44448 202046 44518 202102
rect 44574 202046 44642 202102
rect 44698 202046 44768 202102
rect 44448 201978 44768 202046
rect 44448 201922 44518 201978
rect 44574 201922 44642 201978
rect 44698 201922 44768 201978
rect 44448 201888 44768 201922
rect 39858 190294 39954 190350
rect 40010 190294 40078 190350
rect 40134 190294 40202 190350
rect 40258 190294 40326 190350
rect 40382 190294 40478 190350
rect 39858 190226 40478 190294
rect 39858 190170 39954 190226
rect 40010 190170 40078 190226
rect 40134 190170 40202 190226
rect 40258 190170 40326 190226
rect 40382 190170 40478 190226
rect 39858 190102 40478 190170
rect 39858 190046 39954 190102
rect 40010 190046 40078 190102
rect 40134 190046 40202 190102
rect 40258 190046 40326 190102
rect 40382 190046 40478 190102
rect 39858 189978 40478 190046
rect 39858 189922 39954 189978
rect 40010 189922 40078 189978
rect 40134 189922 40202 189978
rect 40258 189922 40326 189978
rect 40382 189922 40478 189978
rect 39858 172350 40478 189922
rect 44448 184350 44768 184384
rect 44448 184294 44518 184350
rect 44574 184294 44642 184350
rect 44698 184294 44768 184350
rect 44448 184226 44768 184294
rect 44448 184170 44518 184226
rect 44574 184170 44642 184226
rect 44698 184170 44768 184226
rect 44448 184102 44768 184170
rect 44448 184046 44518 184102
rect 44574 184046 44642 184102
rect 44698 184046 44768 184102
rect 44448 183978 44768 184046
rect 44448 183922 44518 183978
rect 44574 183922 44642 183978
rect 44698 183922 44768 183978
rect 44448 183888 44768 183922
rect 39858 172294 39954 172350
rect 40010 172294 40078 172350
rect 40134 172294 40202 172350
rect 40258 172294 40326 172350
rect 40382 172294 40478 172350
rect 39858 172226 40478 172294
rect 39858 172170 39954 172226
rect 40010 172170 40078 172226
rect 40134 172170 40202 172226
rect 40258 172170 40326 172226
rect 40382 172170 40478 172226
rect 39858 172102 40478 172170
rect 39858 172046 39954 172102
rect 40010 172046 40078 172102
rect 40134 172046 40202 172102
rect 40258 172046 40326 172102
rect 40382 172046 40478 172102
rect 39858 171978 40478 172046
rect 39858 171922 39954 171978
rect 40010 171922 40078 171978
rect 40134 171922 40202 171978
rect 40258 171922 40326 171978
rect 40382 171922 40478 171978
rect 39858 154350 40478 171922
rect 44448 166350 44768 166384
rect 44448 166294 44518 166350
rect 44574 166294 44642 166350
rect 44698 166294 44768 166350
rect 44448 166226 44768 166294
rect 44448 166170 44518 166226
rect 44574 166170 44642 166226
rect 44698 166170 44768 166226
rect 44448 166102 44768 166170
rect 44448 166046 44518 166102
rect 44574 166046 44642 166102
rect 44698 166046 44768 166102
rect 44448 165978 44768 166046
rect 44448 165922 44518 165978
rect 44574 165922 44642 165978
rect 44698 165922 44768 165978
rect 44448 165888 44768 165922
rect 39858 154294 39954 154350
rect 40010 154294 40078 154350
rect 40134 154294 40202 154350
rect 40258 154294 40326 154350
rect 40382 154294 40478 154350
rect 39858 154226 40478 154294
rect 39858 154170 39954 154226
rect 40010 154170 40078 154226
rect 40134 154170 40202 154226
rect 40258 154170 40326 154226
rect 40382 154170 40478 154226
rect 39858 154102 40478 154170
rect 39858 154046 39954 154102
rect 40010 154046 40078 154102
rect 40134 154046 40202 154102
rect 40258 154046 40326 154102
rect 40382 154046 40478 154102
rect 39858 153978 40478 154046
rect 39858 153922 39954 153978
rect 40010 153922 40078 153978
rect 40134 153922 40202 153978
rect 40258 153922 40326 153978
rect 40382 153922 40478 153978
rect 39858 136350 40478 153922
rect 44448 148350 44768 148384
rect 44448 148294 44518 148350
rect 44574 148294 44642 148350
rect 44698 148294 44768 148350
rect 44448 148226 44768 148294
rect 44448 148170 44518 148226
rect 44574 148170 44642 148226
rect 44698 148170 44768 148226
rect 44448 148102 44768 148170
rect 44448 148046 44518 148102
rect 44574 148046 44642 148102
rect 44698 148046 44768 148102
rect 44448 147978 44768 148046
rect 44448 147922 44518 147978
rect 44574 147922 44642 147978
rect 44698 147922 44768 147978
rect 44448 147888 44768 147922
rect 39858 136294 39954 136350
rect 40010 136294 40078 136350
rect 40134 136294 40202 136350
rect 40258 136294 40326 136350
rect 40382 136294 40478 136350
rect 39858 136226 40478 136294
rect 39858 136170 39954 136226
rect 40010 136170 40078 136226
rect 40134 136170 40202 136226
rect 40258 136170 40326 136226
rect 40382 136170 40478 136226
rect 39858 136102 40478 136170
rect 39858 136046 39954 136102
rect 40010 136046 40078 136102
rect 40134 136046 40202 136102
rect 40258 136046 40326 136102
rect 40382 136046 40478 136102
rect 39858 135978 40478 136046
rect 39858 135922 39954 135978
rect 40010 135922 40078 135978
rect 40134 135922 40202 135978
rect 40258 135922 40326 135978
rect 40382 135922 40478 135978
rect 39858 118350 40478 135922
rect 44448 130350 44768 130384
rect 44448 130294 44518 130350
rect 44574 130294 44642 130350
rect 44698 130294 44768 130350
rect 44448 130226 44768 130294
rect 44448 130170 44518 130226
rect 44574 130170 44642 130226
rect 44698 130170 44768 130226
rect 44448 130102 44768 130170
rect 44448 130046 44518 130102
rect 44574 130046 44642 130102
rect 44698 130046 44768 130102
rect 44448 129978 44768 130046
rect 44448 129922 44518 129978
rect 44574 129922 44642 129978
rect 44698 129922 44768 129978
rect 44448 129888 44768 129922
rect 39858 118294 39954 118350
rect 40010 118294 40078 118350
rect 40134 118294 40202 118350
rect 40258 118294 40326 118350
rect 40382 118294 40478 118350
rect 39858 118226 40478 118294
rect 39858 118170 39954 118226
rect 40010 118170 40078 118226
rect 40134 118170 40202 118226
rect 40258 118170 40326 118226
rect 40382 118170 40478 118226
rect 39858 118102 40478 118170
rect 39858 118046 39954 118102
rect 40010 118046 40078 118102
rect 40134 118046 40202 118102
rect 40258 118046 40326 118102
rect 40382 118046 40478 118102
rect 39858 117978 40478 118046
rect 39858 117922 39954 117978
rect 40010 117922 40078 117978
rect 40134 117922 40202 117978
rect 40258 117922 40326 117978
rect 40382 117922 40478 117978
rect 39858 100350 40478 117922
rect 44448 112350 44768 112384
rect 44448 112294 44518 112350
rect 44574 112294 44642 112350
rect 44698 112294 44768 112350
rect 44448 112226 44768 112294
rect 44448 112170 44518 112226
rect 44574 112170 44642 112226
rect 44698 112170 44768 112226
rect 44448 112102 44768 112170
rect 44448 112046 44518 112102
rect 44574 112046 44642 112102
rect 44698 112046 44768 112102
rect 44448 111978 44768 112046
rect 44448 111922 44518 111978
rect 44574 111922 44642 111978
rect 44698 111922 44768 111978
rect 44448 111888 44768 111922
rect 39858 100294 39954 100350
rect 40010 100294 40078 100350
rect 40134 100294 40202 100350
rect 40258 100294 40326 100350
rect 40382 100294 40478 100350
rect 39858 100226 40478 100294
rect 39858 100170 39954 100226
rect 40010 100170 40078 100226
rect 40134 100170 40202 100226
rect 40258 100170 40326 100226
rect 40382 100170 40478 100226
rect 39858 100102 40478 100170
rect 39858 100046 39954 100102
rect 40010 100046 40078 100102
rect 40134 100046 40202 100102
rect 40258 100046 40326 100102
rect 40382 100046 40478 100102
rect 39858 99978 40478 100046
rect 39858 99922 39954 99978
rect 40010 99922 40078 99978
rect 40134 99922 40202 99978
rect 40258 99922 40326 99978
rect 40382 99922 40478 99978
rect 39858 82350 40478 99922
rect 44448 94350 44768 94384
rect 44448 94294 44518 94350
rect 44574 94294 44642 94350
rect 44698 94294 44768 94350
rect 44448 94226 44768 94294
rect 44448 94170 44518 94226
rect 44574 94170 44642 94226
rect 44698 94170 44768 94226
rect 44448 94102 44768 94170
rect 44448 94046 44518 94102
rect 44574 94046 44642 94102
rect 44698 94046 44768 94102
rect 44448 93978 44768 94046
rect 44448 93922 44518 93978
rect 44574 93922 44642 93978
rect 44698 93922 44768 93978
rect 44448 93888 44768 93922
rect 39858 82294 39954 82350
rect 40010 82294 40078 82350
rect 40134 82294 40202 82350
rect 40258 82294 40326 82350
rect 40382 82294 40478 82350
rect 39858 82226 40478 82294
rect 39858 82170 39954 82226
rect 40010 82170 40078 82226
rect 40134 82170 40202 82226
rect 40258 82170 40326 82226
rect 40382 82170 40478 82226
rect 39858 82102 40478 82170
rect 39858 82046 39954 82102
rect 40010 82046 40078 82102
rect 40134 82046 40202 82102
rect 40258 82046 40326 82102
rect 40382 82046 40478 82102
rect 39858 81978 40478 82046
rect 39858 81922 39954 81978
rect 40010 81922 40078 81978
rect 40134 81922 40202 81978
rect 40258 81922 40326 81978
rect 40382 81922 40478 81978
rect 39858 64350 40478 81922
rect 44448 76350 44768 76384
rect 44448 76294 44518 76350
rect 44574 76294 44642 76350
rect 44698 76294 44768 76350
rect 44448 76226 44768 76294
rect 44448 76170 44518 76226
rect 44574 76170 44642 76226
rect 44698 76170 44768 76226
rect 44448 76102 44768 76170
rect 44448 76046 44518 76102
rect 44574 76046 44642 76102
rect 44698 76046 44768 76102
rect 44448 75978 44768 76046
rect 44448 75922 44518 75978
rect 44574 75922 44642 75978
rect 44698 75922 44768 75978
rect 44448 75888 44768 75922
rect 39858 64294 39954 64350
rect 40010 64294 40078 64350
rect 40134 64294 40202 64350
rect 40258 64294 40326 64350
rect 40382 64294 40478 64350
rect 39858 64226 40478 64294
rect 39858 64170 39954 64226
rect 40010 64170 40078 64226
rect 40134 64170 40202 64226
rect 40258 64170 40326 64226
rect 40382 64170 40478 64226
rect 39858 64102 40478 64170
rect 39858 64046 39954 64102
rect 40010 64046 40078 64102
rect 40134 64046 40202 64102
rect 40258 64046 40326 64102
rect 40382 64046 40478 64102
rect 39858 63978 40478 64046
rect 39858 63922 39954 63978
rect 40010 63922 40078 63978
rect 40134 63922 40202 63978
rect 40258 63922 40326 63978
rect 40382 63922 40478 63978
rect 39858 46350 40478 63922
rect 44448 58350 44768 58384
rect 44448 58294 44518 58350
rect 44574 58294 44642 58350
rect 44698 58294 44768 58350
rect 44448 58226 44768 58294
rect 44448 58170 44518 58226
rect 44574 58170 44642 58226
rect 44698 58170 44768 58226
rect 44448 58102 44768 58170
rect 44448 58046 44518 58102
rect 44574 58046 44642 58102
rect 44698 58046 44768 58102
rect 44448 57978 44768 58046
rect 44448 57922 44518 57978
rect 44574 57922 44642 57978
rect 44698 57922 44768 57978
rect 44448 57888 44768 57922
rect 48524 48692 48580 297388
rect 75168 292350 75488 292384
rect 75168 292294 75238 292350
rect 75294 292294 75362 292350
rect 75418 292294 75488 292350
rect 75168 292226 75488 292294
rect 75168 292170 75238 292226
rect 75294 292170 75362 292226
rect 75418 292170 75488 292226
rect 75168 292102 75488 292170
rect 75168 292046 75238 292102
rect 75294 292046 75362 292102
rect 75418 292046 75488 292102
rect 75168 291978 75488 292046
rect 75168 291922 75238 291978
rect 75294 291922 75362 291978
rect 75418 291922 75488 291978
rect 75168 291888 75488 291922
rect 97578 292350 98198 309922
rect 97578 292294 97674 292350
rect 97730 292294 97798 292350
rect 97854 292294 97922 292350
rect 97978 292294 98046 292350
rect 98102 292294 98198 292350
rect 97578 292226 98198 292294
rect 97578 292170 97674 292226
rect 97730 292170 97798 292226
rect 97854 292170 97922 292226
rect 97978 292170 98046 292226
rect 98102 292170 98198 292226
rect 97578 292102 98198 292170
rect 97578 292046 97674 292102
rect 97730 292046 97798 292102
rect 97854 292046 97922 292102
rect 97978 292046 98046 292102
rect 98102 292046 98198 292102
rect 97578 291978 98198 292046
rect 97578 291922 97674 291978
rect 97730 291922 97798 291978
rect 97854 291922 97922 291978
rect 97978 291922 98046 291978
rect 98102 291922 98198 291978
rect 59808 280350 60128 280384
rect 59808 280294 59878 280350
rect 59934 280294 60002 280350
rect 60058 280294 60128 280350
rect 59808 280226 60128 280294
rect 59808 280170 59878 280226
rect 59934 280170 60002 280226
rect 60058 280170 60128 280226
rect 59808 280102 60128 280170
rect 59808 280046 59878 280102
rect 59934 280046 60002 280102
rect 60058 280046 60128 280102
rect 59808 279978 60128 280046
rect 59808 279922 59878 279978
rect 59934 279922 60002 279978
rect 60058 279922 60128 279978
rect 59808 279888 60128 279922
rect 90528 280350 90848 280384
rect 90528 280294 90598 280350
rect 90654 280294 90722 280350
rect 90778 280294 90848 280350
rect 90528 280226 90848 280294
rect 90528 280170 90598 280226
rect 90654 280170 90722 280226
rect 90778 280170 90848 280226
rect 90528 280102 90848 280170
rect 90528 280046 90598 280102
rect 90654 280046 90722 280102
rect 90778 280046 90848 280102
rect 90528 279978 90848 280046
rect 90528 279922 90598 279978
rect 90654 279922 90722 279978
rect 90778 279922 90848 279978
rect 90528 279888 90848 279922
rect 75168 274350 75488 274384
rect 75168 274294 75238 274350
rect 75294 274294 75362 274350
rect 75418 274294 75488 274350
rect 75168 274226 75488 274294
rect 75168 274170 75238 274226
rect 75294 274170 75362 274226
rect 75418 274170 75488 274226
rect 75168 274102 75488 274170
rect 75168 274046 75238 274102
rect 75294 274046 75362 274102
rect 75418 274046 75488 274102
rect 75168 273978 75488 274046
rect 75168 273922 75238 273978
rect 75294 273922 75362 273978
rect 75418 273922 75488 273978
rect 75168 273888 75488 273922
rect 97578 274350 98198 291922
rect 97578 274294 97674 274350
rect 97730 274294 97798 274350
rect 97854 274294 97922 274350
rect 97978 274294 98046 274350
rect 98102 274294 98198 274350
rect 97578 274226 98198 274294
rect 97578 274170 97674 274226
rect 97730 274170 97798 274226
rect 97854 274170 97922 274226
rect 97978 274170 98046 274226
rect 98102 274170 98198 274226
rect 97578 274102 98198 274170
rect 97578 274046 97674 274102
rect 97730 274046 97798 274102
rect 97854 274046 97922 274102
rect 97978 274046 98046 274102
rect 98102 274046 98198 274102
rect 97578 273978 98198 274046
rect 97578 273922 97674 273978
rect 97730 273922 97798 273978
rect 97854 273922 97922 273978
rect 97978 273922 98046 273978
rect 98102 273922 98198 273978
rect 59808 262350 60128 262384
rect 59808 262294 59878 262350
rect 59934 262294 60002 262350
rect 60058 262294 60128 262350
rect 59808 262226 60128 262294
rect 59808 262170 59878 262226
rect 59934 262170 60002 262226
rect 60058 262170 60128 262226
rect 59808 262102 60128 262170
rect 59808 262046 59878 262102
rect 59934 262046 60002 262102
rect 60058 262046 60128 262102
rect 59808 261978 60128 262046
rect 59808 261922 59878 261978
rect 59934 261922 60002 261978
rect 60058 261922 60128 261978
rect 59808 261888 60128 261922
rect 90528 262350 90848 262384
rect 90528 262294 90598 262350
rect 90654 262294 90722 262350
rect 90778 262294 90848 262350
rect 90528 262226 90848 262294
rect 90528 262170 90598 262226
rect 90654 262170 90722 262226
rect 90778 262170 90848 262226
rect 90528 262102 90848 262170
rect 90528 262046 90598 262102
rect 90654 262046 90722 262102
rect 90778 262046 90848 262102
rect 90528 261978 90848 262046
rect 90528 261922 90598 261978
rect 90654 261922 90722 261978
rect 90778 261922 90848 261978
rect 90528 261888 90848 261922
rect 75168 256350 75488 256384
rect 75168 256294 75238 256350
rect 75294 256294 75362 256350
rect 75418 256294 75488 256350
rect 75168 256226 75488 256294
rect 75168 256170 75238 256226
rect 75294 256170 75362 256226
rect 75418 256170 75488 256226
rect 75168 256102 75488 256170
rect 75168 256046 75238 256102
rect 75294 256046 75362 256102
rect 75418 256046 75488 256102
rect 75168 255978 75488 256046
rect 75168 255922 75238 255978
rect 75294 255922 75362 255978
rect 75418 255922 75488 255978
rect 75168 255888 75488 255922
rect 97578 256350 98198 273922
rect 97578 256294 97674 256350
rect 97730 256294 97798 256350
rect 97854 256294 97922 256350
rect 97978 256294 98046 256350
rect 98102 256294 98198 256350
rect 97578 256226 98198 256294
rect 97578 256170 97674 256226
rect 97730 256170 97798 256226
rect 97854 256170 97922 256226
rect 97978 256170 98046 256226
rect 98102 256170 98198 256226
rect 97578 256102 98198 256170
rect 97578 256046 97674 256102
rect 97730 256046 97798 256102
rect 97854 256046 97922 256102
rect 97978 256046 98046 256102
rect 98102 256046 98198 256102
rect 97578 255978 98198 256046
rect 97578 255922 97674 255978
rect 97730 255922 97798 255978
rect 97854 255922 97922 255978
rect 97978 255922 98046 255978
rect 98102 255922 98198 255978
rect 59808 244350 60128 244384
rect 59808 244294 59878 244350
rect 59934 244294 60002 244350
rect 60058 244294 60128 244350
rect 59808 244226 60128 244294
rect 59808 244170 59878 244226
rect 59934 244170 60002 244226
rect 60058 244170 60128 244226
rect 59808 244102 60128 244170
rect 59808 244046 59878 244102
rect 59934 244046 60002 244102
rect 60058 244046 60128 244102
rect 59808 243978 60128 244046
rect 59808 243922 59878 243978
rect 59934 243922 60002 243978
rect 60058 243922 60128 243978
rect 59808 243888 60128 243922
rect 66858 238350 67478 245074
rect 66858 238294 66954 238350
rect 67010 238294 67078 238350
rect 67134 238294 67202 238350
rect 67258 238294 67326 238350
rect 67382 238294 67478 238350
rect 66858 238226 67478 238294
rect 66858 238170 66954 238226
rect 67010 238170 67078 238226
rect 67134 238170 67202 238226
rect 67258 238170 67326 238226
rect 67382 238170 67478 238226
rect 66858 238102 67478 238170
rect 66858 238046 66954 238102
rect 67010 238046 67078 238102
rect 67134 238046 67202 238102
rect 67258 238046 67326 238102
rect 67382 238046 67478 238102
rect 66858 237978 67478 238046
rect 66858 237922 66954 237978
rect 67010 237922 67078 237978
rect 67134 237922 67202 237978
rect 67258 237922 67326 237978
rect 67382 237922 67478 237978
rect 51996 231140 52052 231150
rect 51884 216020 51940 216030
rect 50316 210196 50372 210206
rect 49532 210084 49588 210094
rect 49532 164638 49588 210028
rect 50316 206578 50372 210140
rect 50316 206512 50372 206522
rect 49532 164572 49588 164582
rect 48524 48626 48580 48636
rect 39858 46294 39954 46350
rect 40010 46294 40078 46350
rect 40134 46294 40202 46350
rect 40258 46294 40326 46350
rect 40382 46294 40478 46350
rect 39858 46226 40478 46294
rect 39858 46170 39954 46226
rect 40010 46170 40078 46226
rect 40134 46170 40202 46226
rect 40258 46170 40326 46226
rect 40382 46170 40478 46226
rect 39858 46102 40478 46170
rect 39858 46046 39954 46102
rect 40010 46046 40078 46102
rect 40134 46046 40202 46102
rect 40258 46046 40326 46102
rect 40382 46046 40478 46102
rect 39858 45978 40478 46046
rect 39858 45922 39954 45978
rect 40010 45922 40078 45978
rect 40134 45922 40202 45978
rect 40258 45922 40326 45978
rect 40382 45922 40478 45978
rect 39858 28350 40478 45922
rect 39858 28294 39954 28350
rect 40010 28294 40078 28350
rect 40134 28294 40202 28350
rect 40258 28294 40326 28350
rect 40382 28294 40478 28350
rect 39858 28226 40478 28294
rect 39858 28170 39954 28226
rect 40010 28170 40078 28226
rect 40134 28170 40202 28226
rect 40258 28170 40326 28226
rect 40382 28170 40478 28226
rect 39858 28102 40478 28170
rect 39858 28046 39954 28102
rect 40010 28046 40078 28102
rect 40134 28046 40202 28102
rect 40258 28046 40326 28102
rect 40382 28046 40478 28102
rect 39858 27978 40478 28046
rect 39858 27922 39954 27978
rect 40010 27922 40078 27978
rect 40134 27922 40202 27978
rect 40258 27922 40326 27978
rect 40382 27922 40478 27978
rect 39858 10350 40478 27922
rect 39858 10294 39954 10350
rect 40010 10294 40078 10350
rect 40134 10294 40202 10350
rect 40258 10294 40326 10350
rect 40382 10294 40478 10350
rect 39858 10226 40478 10294
rect 39858 10170 39954 10226
rect 40010 10170 40078 10226
rect 40134 10170 40202 10226
rect 40258 10170 40326 10226
rect 40382 10170 40478 10226
rect 39858 10102 40478 10170
rect 39858 10046 39954 10102
rect 40010 10046 40078 10102
rect 40134 10046 40202 10102
rect 40258 10046 40326 10102
rect 40382 10046 40478 10102
rect 39858 9978 40478 10046
rect 39858 9922 39954 9978
rect 40010 9922 40078 9978
rect 40134 9922 40202 9978
rect 40258 9922 40326 9978
rect 40382 9922 40478 9978
rect 39858 -1120 40478 9922
rect 51884 4452 51940 215964
rect 51996 4564 52052 231084
rect 66858 220350 67478 237922
rect 66858 220294 66954 220350
rect 67010 220294 67078 220350
rect 67134 220294 67202 220350
rect 67258 220294 67326 220350
rect 67382 220294 67478 220350
rect 66858 220226 67478 220294
rect 66858 220170 66954 220226
rect 67010 220170 67078 220226
rect 67134 220170 67202 220226
rect 67258 220170 67326 220226
rect 67382 220170 67478 220226
rect 66858 220102 67478 220170
rect 66858 220046 66954 220102
rect 67010 220046 67078 220102
rect 67134 220046 67202 220102
rect 67258 220046 67326 220102
rect 67382 220046 67478 220102
rect 66858 219978 67478 220046
rect 66858 219922 66954 219978
rect 67010 219922 67078 219978
rect 67134 219922 67202 219978
rect 67258 219922 67326 219978
rect 67382 219922 67478 219978
rect 66858 210462 67478 219922
rect 70578 244350 71198 245074
rect 70578 244294 70674 244350
rect 70730 244294 70798 244350
rect 70854 244294 70922 244350
rect 70978 244294 71046 244350
rect 71102 244294 71198 244350
rect 70578 244226 71198 244294
rect 70578 244170 70674 244226
rect 70730 244170 70798 244226
rect 70854 244170 70922 244226
rect 70978 244170 71046 244226
rect 71102 244170 71198 244226
rect 70578 244102 71198 244170
rect 70578 244046 70674 244102
rect 70730 244046 70798 244102
rect 70854 244046 70922 244102
rect 70978 244046 71046 244102
rect 71102 244046 71198 244102
rect 70578 243978 71198 244046
rect 70578 243922 70674 243978
rect 70730 243922 70798 243978
rect 70854 243922 70922 243978
rect 70978 243922 71046 243978
rect 71102 243922 71198 243978
rect 70578 226350 71198 243922
rect 90528 244350 90848 244384
rect 90528 244294 90598 244350
rect 90654 244294 90722 244350
rect 90778 244294 90848 244350
rect 90528 244226 90848 244294
rect 90528 244170 90598 244226
rect 90654 244170 90722 244226
rect 90778 244170 90848 244226
rect 90528 244102 90848 244170
rect 90528 244046 90598 244102
rect 90654 244046 90722 244102
rect 90778 244046 90848 244102
rect 90528 243978 90848 244046
rect 90528 243922 90598 243978
rect 90654 243922 90722 243978
rect 90778 243922 90848 243978
rect 90528 243888 90848 243922
rect 74956 238532 75012 238542
rect 74956 237538 75012 238476
rect 76972 238532 77028 238542
rect 76972 237718 77028 238476
rect 97578 238350 98198 255922
rect 97578 238294 97674 238350
rect 97730 238294 97798 238350
rect 97854 238294 97922 238350
rect 97978 238294 98046 238350
rect 98102 238294 98198 238350
rect 97578 238226 98198 238294
rect 95452 238196 95508 238206
rect 95452 237748 95508 238140
rect 95452 237682 95508 237692
rect 97578 238170 97674 238226
rect 97730 238170 97798 238226
rect 97854 238170 97922 238226
rect 97978 238170 98046 238226
rect 98102 238170 98198 238226
rect 97578 238102 98198 238170
rect 97578 238046 97674 238102
rect 97730 238046 97798 238102
rect 97854 238046 97922 238102
rect 97978 238046 98046 238102
rect 98102 238046 98198 238102
rect 97578 237978 98198 238046
rect 97578 237922 97674 237978
rect 97730 237922 97798 237978
rect 97854 237922 97922 237978
rect 97978 237922 98046 237978
rect 98102 237922 98198 237978
rect 76972 237652 77028 237662
rect 74956 237472 75012 237482
rect 70578 226294 70674 226350
rect 70730 226294 70798 226350
rect 70854 226294 70922 226350
rect 70978 226294 71046 226350
rect 71102 226294 71198 226350
rect 70578 226226 71198 226294
rect 70578 226170 70674 226226
rect 70730 226170 70798 226226
rect 70854 226170 70922 226226
rect 70978 226170 71046 226226
rect 71102 226170 71198 226226
rect 70578 226102 71198 226170
rect 70578 226046 70674 226102
rect 70730 226046 70798 226102
rect 70854 226046 70922 226102
rect 70978 226046 71046 226102
rect 71102 226046 71198 226102
rect 70578 225978 71198 226046
rect 70578 225922 70674 225978
rect 70730 225922 70798 225978
rect 70854 225922 70922 225978
rect 70978 225922 71046 225978
rect 71102 225922 71198 225978
rect 70578 210462 71198 225922
rect 97578 220350 98198 237922
rect 99932 386932 99988 386942
rect 99932 237538 99988 386876
rect 99932 237472 99988 237482
rect 101298 370350 101918 387922
rect 101298 370294 101394 370350
rect 101450 370294 101518 370350
rect 101574 370294 101642 370350
rect 101698 370294 101766 370350
rect 101822 370294 101918 370350
rect 101298 370226 101918 370294
rect 101298 370170 101394 370226
rect 101450 370170 101518 370226
rect 101574 370170 101642 370226
rect 101698 370170 101766 370226
rect 101822 370170 101918 370226
rect 101298 370102 101918 370170
rect 101298 370046 101394 370102
rect 101450 370046 101518 370102
rect 101574 370046 101642 370102
rect 101698 370046 101766 370102
rect 101822 370046 101918 370102
rect 101298 369978 101918 370046
rect 101298 369922 101394 369978
rect 101450 369922 101518 369978
rect 101574 369922 101642 369978
rect 101698 369922 101766 369978
rect 101822 369922 101918 369978
rect 101298 352350 101918 369922
rect 101298 352294 101394 352350
rect 101450 352294 101518 352350
rect 101574 352294 101642 352350
rect 101698 352294 101766 352350
rect 101822 352294 101918 352350
rect 101298 352226 101918 352294
rect 101298 352170 101394 352226
rect 101450 352170 101518 352226
rect 101574 352170 101642 352226
rect 101698 352170 101766 352226
rect 101822 352170 101918 352226
rect 101298 352102 101918 352170
rect 101298 352046 101394 352102
rect 101450 352046 101518 352102
rect 101574 352046 101642 352102
rect 101698 352046 101766 352102
rect 101822 352046 101918 352102
rect 101298 351978 101918 352046
rect 101298 351922 101394 351978
rect 101450 351922 101518 351978
rect 101574 351922 101642 351978
rect 101698 351922 101766 351978
rect 101822 351922 101918 351978
rect 101298 334350 101918 351922
rect 101298 334294 101394 334350
rect 101450 334294 101518 334350
rect 101574 334294 101642 334350
rect 101698 334294 101766 334350
rect 101822 334294 101918 334350
rect 101298 334226 101918 334294
rect 101298 334170 101394 334226
rect 101450 334170 101518 334226
rect 101574 334170 101642 334226
rect 101698 334170 101766 334226
rect 101822 334170 101918 334226
rect 101298 334102 101918 334170
rect 101298 334046 101394 334102
rect 101450 334046 101518 334102
rect 101574 334046 101642 334102
rect 101698 334046 101766 334102
rect 101822 334046 101918 334102
rect 101298 333978 101918 334046
rect 101298 333922 101394 333978
rect 101450 333922 101518 333978
rect 101574 333922 101642 333978
rect 101698 333922 101766 333978
rect 101822 333922 101918 333978
rect 101298 316350 101918 333922
rect 101298 316294 101394 316350
rect 101450 316294 101518 316350
rect 101574 316294 101642 316350
rect 101698 316294 101766 316350
rect 101822 316294 101918 316350
rect 101298 316226 101918 316294
rect 101298 316170 101394 316226
rect 101450 316170 101518 316226
rect 101574 316170 101642 316226
rect 101698 316170 101766 316226
rect 101822 316170 101918 316226
rect 101298 316102 101918 316170
rect 101298 316046 101394 316102
rect 101450 316046 101518 316102
rect 101574 316046 101642 316102
rect 101698 316046 101766 316102
rect 101822 316046 101918 316102
rect 101298 315978 101918 316046
rect 101298 315922 101394 315978
rect 101450 315922 101518 315978
rect 101574 315922 101642 315978
rect 101698 315922 101766 315978
rect 101822 315922 101918 315978
rect 101298 298350 101918 315922
rect 101298 298294 101394 298350
rect 101450 298294 101518 298350
rect 101574 298294 101642 298350
rect 101698 298294 101766 298350
rect 101822 298294 101918 298350
rect 101298 298226 101918 298294
rect 101298 298170 101394 298226
rect 101450 298170 101518 298226
rect 101574 298170 101642 298226
rect 101698 298170 101766 298226
rect 101822 298170 101918 298226
rect 101298 298102 101918 298170
rect 101298 298046 101394 298102
rect 101450 298046 101518 298102
rect 101574 298046 101642 298102
rect 101698 298046 101766 298102
rect 101822 298046 101918 298102
rect 101298 297978 101918 298046
rect 101298 297922 101394 297978
rect 101450 297922 101518 297978
rect 101574 297922 101642 297978
rect 101698 297922 101766 297978
rect 101822 297922 101918 297978
rect 101298 280350 101918 297922
rect 101298 280294 101394 280350
rect 101450 280294 101518 280350
rect 101574 280294 101642 280350
rect 101698 280294 101766 280350
rect 101822 280294 101918 280350
rect 101298 280226 101918 280294
rect 101298 280170 101394 280226
rect 101450 280170 101518 280226
rect 101574 280170 101642 280226
rect 101698 280170 101766 280226
rect 101822 280170 101918 280226
rect 101298 280102 101918 280170
rect 101298 280046 101394 280102
rect 101450 280046 101518 280102
rect 101574 280046 101642 280102
rect 101698 280046 101766 280102
rect 101822 280046 101918 280102
rect 101298 279978 101918 280046
rect 101298 279922 101394 279978
rect 101450 279922 101518 279978
rect 101574 279922 101642 279978
rect 101698 279922 101766 279978
rect 101822 279922 101918 279978
rect 101298 262350 101918 279922
rect 101298 262294 101394 262350
rect 101450 262294 101518 262350
rect 101574 262294 101642 262350
rect 101698 262294 101766 262350
rect 101822 262294 101918 262350
rect 101298 262226 101918 262294
rect 101298 262170 101394 262226
rect 101450 262170 101518 262226
rect 101574 262170 101642 262226
rect 101698 262170 101766 262226
rect 101822 262170 101918 262226
rect 101298 262102 101918 262170
rect 101298 262046 101394 262102
rect 101450 262046 101518 262102
rect 101574 262046 101642 262102
rect 101698 262046 101766 262102
rect 101822 262046 101918 262102
rect 101298 261978 101918 262046
rect 101298 261922 101394 261978
rect 101450 261922 101518 261978
rect 101574 261922 101642 261978
rect 101698 261922 101766 261978
rect 101822 261922 101918 261978
rect 101298 244350 101918 261922
rect 101298 244294 101394 244350
rect 101450 244294 101518 244350
rect 101574 244294 101642 244350
rect 101698 244294 101766 244350
rect 101822 244294 101918 244350
rect 101298 244226 101918 244294
rect 101298 244170 101394 244226
rect 101450 244170 101518 244226
rect 101574 244170 101642 244226
rect 101698 244170 101766 244226
rect 101822 244170 101918 244226
rect 101298 244102 101918 244170
rect 101298 244046 101394 244102
rect 101450 244046 101518 244102
rect 101574 244046 101642 244102
rect 101698 244046 101766 244102
rect 101822 244046 101918 244102
rect 101298 243978 101918 244046
rect 101298 243922 101394 243978
rect 101450 243922 101518 243978
rect 101574 243922 101642 243978
rect 101698 243922 101766 243978
rect 101822 243922 101918 243978
rect 97578 220294 97674 220350
rect 97730 220294 97798 220350
rect 97854 220294 97922 220350
rect 97978 220294 98046 220350
rect 98102 220294 98198 220350
rect 97578 220226 98198 220294
rect 97578 220170 97674 220226
rect 97730 220170 97798 220226
rect 97854 220170 97922 220226
rect 97978 220170 98046 220226
rect 98102 220170 98198 220226
rect 97578 220102 98198 220170
rect 97578 220046 97674 220102
rect 97730 220046 97798 220102
rect 97854 220046 97922 220102
rect 97978 220046 98046 220102
rect 98102 220046 98198 220102
rect 97578 219978 98198 220046
rect 97578 219922 97674 219978
rect 97730 219922 97798 219978
rect 97854 219922 97922 219978
rect 97978 219922 98046 219978
rect 98102 219922 98198 219978
rect 97578 210462 98198 219922
rect 101298 226350 101918 243922
rect 103292 391748 103348 391758
rect 103292 237718 103348 391692
rect 103292 237652 103348 237662
rect 128298 382350 128918 399922
rect 128298 382294 128394 382350
rect 128450 382294 128518 382350
rect 128574 382294 128642 382350
rect 128698 382294 128766 382350
rect 128822 382294 128918 382350
rect 128298 382226 128918 382294
rect 128298 382170 128394 382226
rect 128450 382170 128518 382226
rect 128574 382170 128642 382226
rect 128698 382170 128766 382226
rect 128822 382170 128918 382226
rect 128298 382102 128918 382170
rect 128298 382046 128394 382102
rect 128450 382046 128518 382102
rect 128574 382046 128642 382102
rect 128698 382046 128766 382102
rect 128822 382046 128918 382102
rect 128298 381978 128918 382046
rect 128298 381922 128394 381978
rect 128450 381922 128518 381978
rect 128574 381922 128642 381978
rect 128698 381922 128766 381978
rect 128822 381922 128918 381978
rect 128298 364350 128918 381922
rect 128298 364294 128394 364350
rect 128450 364294 128518 364350
rect 128574 364294 128642 364350
rect 128698 364294 128766 364350
rect 128822 364294 128918 364350
rect 128298 364226 128918 364294
rect 128298 364170 128394 364226
rect 128450 364170 128518 364226
rect 128574 364170 128642 364226
rect 128698 364170 128766 364226
rect 128822 364170 128918 364226
rect 128298 364102 128918 364170
rect 128298 364046 128394 364102
rect 128450 364046 128518 364102
rect 128574 364046 128642 364102
rect 128698 364046 128766 364102
rect 128822 364046 128918 364102
rect 128298 363978 128918 364046
rect 128298 363922 128394 363978
rect 128450 363922 128518 363978
rect 128574 363922 128642 363978
rect 128698 363922 128766 363978
rect 128822 363922 128918 363978
rect 128298 346350 128918 363922
rect 128298 346294 128394 346350
rect 128450 346294 128518 346350
rect 128574 346294 128642 346350
rect 128698 346294 128766 346350
rect 128822 346294 128918 346350
rect 128298 346226 128918 346294
rect 128298 346170 128394 346226
rect 128450 346170 128518 346226
rect 128574 346170 128642 346226
rect 128698 346170 128766 346226
rect 128822 346170 128918 346226
rect 128298 346102 128918 346170
rect 128298 346046 128394 346102
rect 128450 346046 128518 346102
rect 128574 346046 128642 346102
rect 128698 346046 128766 346102
rect 128822 346046 128918 346102
rect 128298 345978 128918 346046
rect 128298 345922 128394 345978
rect 128450 345922 128518 345978
rect 128574 345922 128642 345978
rect 128698 345922 128766 345978
rect 128822 345922 128918 345978
rect 128298 328350 128918 345922
rect 128298 328294 128394 328350
rect 128450 328294 128518 328350
rect 128574 328294 128642 328350
rect 128698 328294 128766 328350
rect 128822 328294 128918 328350
rect 128298 328226 128918 328294
rect 128298 328170 128394 328226
rect 128450 328170 128518 328226
rect 128574 328170 128642 328226
rect 128698 328170 128766 328226
rect 128822 328170 128918 328226
rect 128298 328102 128918 328170
rect 128298 328046 128394 328102
rect 128450 328046 128518 328102
rect 128574 328046 128642 328102
rect 128698 328046 128766 328102
rect 128822 328046 128918 328102
rect 128298 327978 128918 328046
rect 128298 327922 128394 327978
rect 128450 327922 128518 327978
rect 128574 327922 128642 327978
rect 128698 327922 128766 327978
rect 128822 327922 128918 327978
rect 128298 310350 128918 327922
rect 128298 310294 128394 310350
rect 128450 310294 128518 310350
rect 128574 310294 128642 310350
rect 128698 310294 128766 310350
rect 128822 310294 128918 310350
rect 128298 310226 128918 310294
rect 128298 310170 128394 310226
rect 128450 310170 128518 310226
rect 128574 310170 128642 310226
rect 128698 310170 128766 310226
rect 128822 310170 128918 310226
rect 128298 310102 128918 310170
rect 128298 310046 128394 310102
rect 128450 310046 128518 310102
rect 128574 310046 128642 310102
rect 128698 310046 128766 310102
rect 128822 310046 128918 310102
rect 128298 309978 128918 310046
rect 128298 309922 128394 309978
rect 128450 309922 128518 309978
rect 128574 309922 128642 309978
rect 128698 309922 128766 309978
rect 128822 309922 128918 309978
rect 128298 292350 128918 309922
rect 128298 292294 128394 292350
rect 128450 292294 128518 292350
rect 128574 292294 128642 292350
rect 128698 292294 128766 292350
rect 128822 292294 128918 292350
rect 128298 292226 128918 292294
rect 128298 292170 128394 292226
rect 128450 292170 128518 292226
rect 128574 292170 128642 292226
rect 128698 292170 128766 292226
rect 128822 292170 128918 292226
rect 128298 292102 128918 292170
rect 128298 292046 128394 292102
rect 128450 292046 128518 292102
rect 128574 292046 128642 292102
rect 128698 292046 128766 292102
rect 128822 292046 128918 292102
rect 128298 291978 128918 292046
rect 128298 291922 128394 291978
rect 128450 291922 128518 291978
rect 128574 291922 128642 291978
rect 128698 291922 128766 291978
rect 128822 291922 128918 291978
rect 128298 274350 128918 291922
rect 128298 274294 128394 274350
rect 128450 274294 128518 274350
rect 128574 274294 128642 274350
rect 128698 274294 128766 274350
rect 128822 274294 128918 274350
rect 128298 274226 128918 274294
rect 128298 274170 128394 274226
rect 128450 274170 128518 274226
rect 128574 274170 128642 274226
rect 128698 274170 128766 274226
rect 128822 274170 128918 274226
rect 128298 274102 128918 274170
rect 128298 274046 128394 274102
rect 128450 274046 128518 274102
rect 128574 274046 128642 274102
rect 128698 274046 128766 274102
rect 128822 274046 128918 274102
rect 128298 273978 128918 274046
rect 128298 273922 128394 273978
rect 128450 273922 128518 273978
rect 128574 273922 128642 273978
rect 128698 273922 128766 273978
rect 128822 273922 128918 273978
rect 128298 256350 128918 273922
rect 128298 256294 128394 256350
rect 128450 256294 128518 256350
rect 128574 256294 128642 256350
rect 128698 256294 128766 256350
rect 128822 256294 128918 256350
rect 128298 256226 128918 256294
rect 128298 256170 128394 256226
rect 128450 256170 128518 256226
rect 128574 256170 128642 256226
rect 128698 256170 128766 256226
rect 128822 256170 128918 256226
rect 128298 256102 128918 256170
rect 128298 256046 128394 256102
rect 128450 256046 128518 256102
rect 128574 256046 128642 256102
rect 128698 256046 128766 256102
rect 128822 256046 128918 256102
rect 128298 255978 128918 256046
rect 128298 255922 128394 255978
rect 128450 255922 128518 255978
rect 128574 255922 128642 255978
rect 128698 255922 128766 255978
rect 128822 255922 128918 255978
rect 128298 238350 128918 255922
rect 128298 238294 128394 238350
rect 128450 238294 128518 238350
rect 128574 238294 128642 238350
rect 128698 238294 128766 238350
rect 128822 238294 128918 238350
rect 128298 238226 128918 238294
rect 128298 238170 128394 238226
rect 128450 238170 128518 238226
rect 128574 238170 128642 238226
rect 128698 238170 128766 238226
rect 128822 238170 128918 238226
rect 128298 238102 128918 238170
rect 128298 238046 128394 238102
rect 128450 238046 128518 238102
rect 128574 238046 128642 238102
rect 128698 238046 128766 238102
rect 128822 238046 128918 238102
rect 128298 237978 128918 238046
rect 128298 237922 128394 237978
rect 128450 237922 128518 237978
rect 128574 237922 128642 237978
rect 128698 237922 128766 237978
rect 128822 237922 128918 237978
rect 101298 226294 101394 226350
rect 101450 226294 101518 226350
rect 101574 226294 101642 226350
rect 101698 226294 101766 226350
rect 101822 226294 101918 226350
rect 101298 226226 101918 226294
rect 101298 226170 101394 226226
rect 101450 226170 101518 226226
rect 101574 226170 101642 226226
rect 101698 226170 101766 226226
rect 101822 226170 101918 226226
rect 101298 226102 101918 226170
rect 101298 226046 101394 226102
rect 101450 226046 101518 226102
rect 101574 226046 101642 226102
rect 101698 226046 101766 226102
rect 101822 226046 101918 226102
rect 101298 225978 101918 226046
rect 101298 225922 101394 225978
rect 101450 225922 101518 225978
rect 101574 225922 101642 225978
rect 101698 225922 101766 225978
rect 101822 225922 101918 225978
rect 101298 210462 101918 225922
rect 128298 220350 128918 237922
rect 128298 220294 128394 220350
rect 128450 220294 128518 220350
rect 128574 220294 128642 220350
rect 128698 220294 128766 220350
rect 128822 220294 128918 220350
rect 128298 220226 128918 220294
rect 128298 220170 128394 220226
rect 128450 220170 128518 220226
rect 128574 220170 128642 220226
rect 128698 220170 128766 220226
rect 128822 220170 128918 220226
rect 128298 220102 128918 220170
rect 128298 220046 128394 220102
rect 128450 220046 128518 220102
rect 128574 220046 128642 220102
rect 128698 220046 128766 220102
rect 128822 220046 128918 220102
rect 128298 219978 128918 220046
rect 128298 219922 128394 219978
rect 128450 219922 128518 219978
rect 128574 219922 128642 219978
rect 128698 219922 128766 219978
rect 128822 219922 128918 219978
rect 128298 210462 128918 219922
rect 132018 496350 132638 500388
rect 132018 496294 132114 496350
rect 132170 496294 132238 496350
rect 132294 496294 132362 496350
rect 132418 496294 132486 496350
rect 132542 496294 132638 496350
rect 132018 496226 132638 496294
rect 132018 496170 132114 496226
rect 132170 496170 132238 496226
rect 132294 496170 132362 496226
rect 132418 496170 132486 496226
rect 132542 496170 132638 496226
rect 132018 496102 132638 496170
rect 132018 496046 132114 496102
rect 132170 496046 132238 496102
rect 132294 496046 132362 496102
rect 132418 496046 132486 496102
rect 132542 496046 132638 496102
rect 132018 495978 132638 496046
rect 132018 495922 132114 495978
rect 132170 495922 132238 495978
rect 132294 495922 132362 495978
rect 132418 495922 132486 495978
rect 132542 495922 132638 495978
rect 132018 478350 132638 495922
rect 132018 478294 132114 478350
rect 132170 478294 132238 478350
rect 132294 478294 132362 478350
rect 132418 478294 132486 478350
rect 132542 478294 132638 478350
rect 132018 478226 132638 478294
rect 132018 478170 132114 478226
rect 132170 478170 132238 478226
rect 132294 478170 132362 478226
rect 132418 478170 132486 478226
rect 132542 478170 132638 478226
rect 132018 478102 132638 478170
rect 132018 478046 132114 478102
rect 132170 478046 132238 478102
rect 132294 478046 132362 478102
rect 132418 478046 132486 478102
rect 132542 478046 132638 478102
rect 132018 477978 132638 478046
rect 132018 477922 132114 477978
rect 132170 477922 132238 477978
rect 132294 477922 132362 477978
rect 132418 477922 132486 477978
rect 132542 477922 132638 477978
rect 132018 460350 132638 477922
rect 159018 490350 159638 507922
rect 159018 490294 159114 490350
rect 159170 490294 159238 490350
rect 159294 490294 159362 490350
rect 159418 490294 159486 490350
rect 159542 490294 159638 490350
rect 159018 490226 159638 490294
rect 159018 490170 159114 490226
rect 159170 490170 159238 490226
rect 159294 490170 159362 490226
rect 159418 490170 159486 490226
rect 159542 490170 159638 490226
rect 159018 490102 159638 490170
rect 159018 490046 159114 490102
rect 159170 490046 159238 490102
rect 159294 490046 159362 490102
rect 159418 490046 159486 490102
rect 159542 490046 159638 490102
rect 159018 489978 159638 490046
rect 159018 489922 159114 489978
rect 159170 489922 159238 489978
rect 159294 489922 159362 489978
rect 159418 489922 159486 489978
rect 159542 489922 159638 489978
rect 146972 476308 147028 476318
rect 132018 460294 132114 460350
rect 132170 460294 132238 460350
rect 132294 460294 132362 460350
rect 132418 460294 132486 460350
rect 132542 460294 132638 460350
rect 132018 460226 132638 460294
rect 132018 460170 132114 460226
rect 132170 460170 132238 460226
rect 132294 460170 132362 460226
rect 132418 460170 132486 460226
rect 132542 460170 132638 460226
rect 132018 460102 132638 460170
rect 132018 460046 132114 460102
rect 132170 460046 132238 460102
rect 132294 460046 132362 460102
rect 132418 460046 132486 460102
rect 132542 460046 132638 460102
rect 132018 459978 132638 460046
rect 132018 459922 132114 459978
rect 132170 459922 132238 459978
rect 132294 459922 132362 459978
rect 132418 459922 132486 459978
rect 132542 459922 132638 459978
rect 132018 442350 132638 459922
rect 132018 442294 132114 442350
rect 132170 442294 132238 442350
rect 132294 442294 132362 442350
rect 132418 442294 132486 442350
rect 132542 442294 132638 442350
rect 132018 442226 132638 442294
rect 132018 442170 132114 442226
rect 132170 442170 132238 442226
rect 132294 442170 132362 442226
rect 132418 442170 132486 442226
rect 132542 442170 132638 442226
rect 132018 442102 132638 442170
rect 132018 442046 132114 442102
rect 132170 442046 132238 442102
rect 132294 442046 132362 442102
rect 132418 442046 132486 442102
rect 132542 442046 132638 442102
rect 132018 441978 132638 442046
rect 132018 441922 132114 441978
rect 132170 441922 132238 441978
rect 132294 441922 132362 441978
rect 132418 441922 132486 441978
rect 132542 441922 132638 441978
rect 132018 424350 132638 441922
rect 141932 474292 141988 474302
rect 132018 424294 132114 424350
rect 132170 424294 132238 424350
rect 132294 424294 132362 424350
rect 132418 424294 132486 424350
rect 132542 424294 132638 424350
rect 132018 424226 132638 424294
rect 132018 424170 132114 424226
rect 132170 424170 132238 424226
rect 132294 424170 132362 424226
rect 132418 424170 132486 424226
rect 132542 424170 132638 424226
rect 132018 424102 132638 424170
rect 132018 424046 132114 424102
rect 132170 424046 132238 424102
rect 132294 424046 132362 424102
rect 132418 424046 132486 424102
rect 132542 424046 132638 424102
rect 132018 423978 132638 424046
rect 132018 423922 132114 423978
rect 132170 423922 132238 423978
rect 132294 423922 132362 423978
rect 132418 423922 132486 423978
rect 132542 423922 132638 423978
rect 132018 406350 132638 423922
rect 132018 406294 132114 406350
rect 132170 406294 132238 406350
rect 132294 406294 132362 406350
rect 132418 406294 132486 406350
rect 132542 406294 132638 406350
rect 132018 406226 132638 406294
rect 132018 406170 132114 406226
rect 132170 406170 132238 406226
rect 132294 406170 132362 406226
rect 132418 406170 132486 406226
rect 132542 406170 132638 406226
rect 132018 406102 132638 406170
rect 132018 406046 132114 406102
rect 132170 406046 132238 406102
rect 132294 406046 132362 406102
rect 132418 406046 132486 406102
rect 132542 406046 132638 406102
rect 132018 405978 132638 406046
rect 132018 405922 132114 405978
rect 132170 405922 132238 405978
rect 132294 405922 132362 405978
rect 132418 405922 132486 405978
rect 132542 405922 132638 405978
rect 132018 388350 132638 405922
rect 132018 388294 132114 388350
rect 132170 388294 132238 388350
rect 132294 388294 132362 388350
rect 132418 388294 132486 388350
rect 132542 388294 132638 388350
rect 132018 388226 132638 388294
rect 132018 388170 132114 388226
rect 132170 388170 132238 388226
rect 132294 388170 132362 388226
rect 132418 388170 132486 388226
rect 132542 388170 132638 388226
rect 132018 388102 132638 388170
rect 132018 388046 132114 388102
rect 132170 388046 132238 388102
rect 132294 388046 132362 388102
rect 132418 388046 132486 388102
rect 132542 388046 132638 388102
rect 132018 387978 132638 388046
rect 132018 387922 132114 387978
rect 132170 387922 132238 387978
rect 132294 387922 132362 387978
rect 132418 387922 132486 387978
rect 132542 387922 132638 387978
rect 132018 370350 132638 387922
rect 132018 370294 132114 370350
rect 132170 370294 132238 370350
rect 132294 370294 132362 370350
rect 132418 370294 132486 370350
rect 132542 370294 132638 370350
rect 132018 370226 132638 370294
rect 132018 370170 132114 370226
rect 132170 370170 132238 370226
rect 132294 370170 132362 370226
rect 132418 370170 132486 370226
rect 132542 370170 132638 370226
rect 132018 370102 132638 370170
rect 132018 370046 132114 370102
rect 132170 370046 132238 370102
rect 132294 370046 132362 370102
rect 132418 370046 132486 370102
rect 132542 370046 132638 370102
rect 132018 369978 132638 370046
rect 132018 369922 132114 369978
rect 132170 369922 132238 369978
rect 132294 369922 132362 369978
rect 132418 369922 132486 369978
rect 132542 369922 132638 369978
rect 132018 352350 132638 369922
rect 132018 352294 132114 352350
rect 132170 352294 132238 352350
rect 132294 352294 132362 352350
rect 132418 352294 132486 352350
rect 132542 352294 132638 352350
rect 132018 352226 132638 352294
rect 132018 352170 132114 352226
rect 132170 352170 132238 352226
rect 132294 352170 132362 352226
rect 132418 352170 132486 352226
rect 132542 352170 132638 352226
rect 132018 352102 132638 352170
rect 132018 352046 132114 352102
rect 132170 352046 132238 352102
rect 132294 352046 132362 352102
rect 132418 352046 132486 352102
rect 132542 352046 132638 352102
rect 132018 351978 132638 352046
rect 132018 351922 132114 351978
rect 132170 351922 132238 351978
rect 132294 351922 132362 351978
rect 132418 351922 132486 351978
rect 132542 351922 132638 351978
rect 132018 334350 132638 351922
rect 140252 431956 140308 431966
rect 132018 334294 132114 334350
rect 132170 334294 132238 334350
rect 132294 334294 132362 334350
rect 132418 334294 132486 334350
rect 132542 334294 132638 334350
rect 132018 334226 132638 334294
rect 132018 334170 132114 334226
rect 132170 334170 132238 334226
rect 132294 334170 132362 334226
rect 132418 334170 132486 334226
rect 132542 334170 132638 334226
rect 132018 334102 132638 334170
rect 132018 334046 132114 334102
rect 132170 334046 132238 334102
rect 132294 334046 132362 334102
rect 132418 334046 132486 334102
rect 132542 334046 132638 334102
rect 132018 333978 132638 334046
rect 132018 333922 132114 333978
rect 132170 333922 132238 333978
rect 132294 333922 132362 333978
rect 132418 333922 132486 333978
rect 132542 333922 132638 333978
rect 132018 316350 132638 333922
rect 132018 316294 132114 316350
rect 132170 316294 132238 316350
rect 132294 316294 132362 316350
rect 132418 316294 132486 316350
rect 132542 316294 132638 316350
rect 132018 316226 132638 316294
rect 132018 316170 132114 316226
rect 132170 316170 132238 316226
rect 132294 316170 132362 316226
rect 132418 316170 132486 316226
rect 132542 316170 132638 316226
rect 132018 316102 132638 316170
rect 132018 316046 132114 316102
rect 132170 316046 132238 316102
rect 132294 316046 132362 316102
rect 132418 316046 132486 316102
rect 132542 316046 132638 316102
rect 132018 315978 132638 316046
rect 132018 315922 132114 315978
rect 132170 315922 132238 315978
rect 132294 315922 132362 315978
rect 132418 315922 132486 315978
rect 132542 315922 132638 315978
rect 132018 298350 132638 315922
rect 132018 298294 132114 298350
rect 132170 298294 132238 298350
rect 132294 298294 132362 298350
rect 132418 298294 132486 298350
rect 132542 298294 132638 298350
rect 132018 298226 132638 298294
rect 132018 298170 132114 298226
rect 132170 298170 132238 298226
rect 132294 298170 132362 298226
rect 132418 298170 132486 298226
rect 132542 298170 132638 298226
rect 132018 298102 132638 298170
rect 132018 298046 132114 298102
rect 132170 298046 132238 298102
rect 132294 298046 132362 298102
rect 132418 298046 132486 298102
rect 132542 298046 132638 298102
rect 132018 297978 132638 298046
rect 132018 297922 132114 297978
rect 132170 297922 132238 297978
rect 132294 297922 132362 297978
rect 132418 297922 132486 297978
rect 132542 297922 132638 297978
rect 132018 280350 132638 297922
rect 138572 345268 138628 345278
rect 138572 296884 138628 345212
rect 138572 296818 138628 296828
rect 140252 294644 140308 431900
rect 140252 294578 140308 294588
rect 141932 293524 141988 474236
rect 141932 293458 141988 293468
rect 145292 469588 145348 469598
rect 145292 292404 145348 469532
rect 145292 292338 145348 292348
rect 146972 291284 147028 476252
rect 159018 472350 159638 489922
rect 159018 472294 159114 472350
rect 159170 472294 159238 472350
rect 159294 472294 159362 472350
rect 159418 472294 159486 472350
rect 159542 472294 159638 472350
rect 159018 472226 159638 472294
rect 159018 472170 159114 472226
rect 159170 472170 159238 472226
rect 159294 472170 159362 472226
rect 159418 472170 159486 472226
rect 159542 472170 159638 472226
rect 159018 472102 159638 472170
rect 159018 472046 159114 472102
rect 159170 472046 159238 472102
rect 159294 472046 159362 472102
rect 159418 472046 159486 472102
rect 159542 472046 159638 472102
rect 159018 471978 159638 472046
rect 159018 471922 159114 471978
rect 159170 471922 159238 471978
rect 159294 471922 159362 471978
rect 159418 471922 159486 471978
rect 159542 471922 159638 471978
rect 159018 454350 159638 471922
rect 162738 598172 163358 598268
rect 162738 598116 162834 598172
rect 162890 598116 162958 598172
rect 163014 598116 163082 598172
rect 163138 598116 163206 598172
rect 163262 598116 163358 598172
rect 162738 598048 163358 598116
rect 162738 597992 162834 598048
rect 162890 597992 162958 598048
rect 163014 597992 163082 598048
rect 163138 597992 163206 598048
rect 163262 597992 163358 598048
rect 162738 597924 163358 597992
rect 162738 597868 162834 597924
rect 162890 597868 162958 597924
rect 163014 597868 163082 597924
rect 163138 597868 163206 597924
rect 163262 597868 163358 597924
rect 162738 597800 163358 597868
rect 162738 597744 162834 597800
rect 162890 597744 162958 597800
rect 163014 597744 163082 597800
rect 163138 597744 163206 597800
rect 163262 597744 163358 597800
rect 162738 586350 163358 597744
rect 162738 586294 162834 586350
rect 162890 586294 162958 586350
rect 163014 586294 163082 586350
rect 163138 586294 163206 586350
rect 163262 586294 163358 586350
rect 162738 586226 163358 586294
rect 162738 586170 162834 586226
rect 162890 586170 162958 586226
rect 163014 586170 163082 586226
rect 163138 586170 163206 586226
rect 163262 586170 163358 586226
rect 162738 586102 163358 586170
rect 162738 586046 162834 586102
rect 162890 586046 162958 586102
rect 163014 586046 163082 586102
rect 163138 586046 163206 586102
rect 163262 586046 163358 586102
rect 162738 585978 163358 586046
rect 162738 585922 162834 585978
rect 162890 585922 162958 585978
rect 163014 585922 163082 585978
rect 163138 585922 163206 585978
rect 163262 585922 163358 585978
rect 162738 568350 163358 585922
rect 162738 568294 162834 568350
rect 162890 568294 162958 568350
rect 163014 568294 163082 568350
rect 163138 568294 163206 568350
rect 163262 568294 163358 568350
rect 162738 568226 163358 568294
rect 162738 568170 162834 568226
rect 162890 568170 162958 568226
rect 163014 568170 163082 568226
rect 163138 568170 163206 568226
rect 163262 568170 163358 568226
rect 162738 568102 163358 568170
rect 162738 568046 162834 568102
rect 162890 568046 162958 568102
rect 163014 568046 163082 568102
rect 163138 568046 163206 568102
rect 163262 568046 163358 568102
rect 162738 567978 163358 568046
rect 162738 567922 162834 567978
rect 162890 567922 162958 567978
rect 163014 567922 163082 567978
rect 163138 567922 163206 567978
rect 163262 567922 163358 567978
rect 162738 550350 163358 567922
rect 189738 597212 190358 598268
rect 189738 597156 189834 597212
rect 189890 597156 189958 597212
rect 190014 597156 190082 597212
rect 190138 597156 190206 597212
rect 190262 597156 190358 597212
rect 189738 597088 190358 597156
rect 189738 597032 189834 597088
rect 189890 597032 189958 597088
rect 190014 597032 190082 597088
rect 190138 597032 190206 597088
rect 190262 597032 190358 597088
rect 189738 596964 190358 597032
rect 189738 596908 189834 596964
rect 189890 596908 189958 596964
rect 190014 596908 190082 596964
rect 190138 596908 190206 596964
rect 190262 596908 190358 596964
rect 189738 596840 190358 596908
rect 189738 596784 189834 596840
rect 189890 596784 189958 596840
rect 190014 596784 190082 596840
rect 190138 596784 190206 596840
rect 190262 596784 190358 596840
rect 189738 580350 190358 596784
rect 193458 598172 194078 598268
rect 193458 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 194078 598172
rect 193458 598048 194078 598116
rect 193458 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 194078 598048
rect 193458 597924 194078 597992
rect 193458 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 194078 597924
rect 193458 597800 194078 597868
rect 193458 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 194078 597800
rect 189738 580294 189834 580350
rect 189890 580294 189958 580350
rect 190014 580294 190082 580350
rect 190138 580294 190206 580350
rect 190262 580294 190358 580350
rect 189738 580226 190358 580294
rect 189738 580170 189834 580226
rect 189890 580170 189958 580226
rect 190014 580170 190082 580226
rect 190138 580170 190206 580226
rect 190262 580170 190358 580226
rect 189738 580102 190358 580170
rect 189738 580046 189834 580102
rect 189890 580046 189958 580102
rect 190014 580046 190082 580102
rect 190138 580046 190206 580102
rect 190262 580046 190358 580102
rect 189738 579978 190358 580046
rect 189738 579922 189834 579978
rect 189890 579922 189958 579978
rect 190014 579922 190082 579978
rect 190138 579922 190206 579978
rect 190262 579922 190358 579978
rect 162738 550294 162834 550350
rect 162890 550294 162958 550350
rect 163014 550294 163082 550350
rect 163138 550294 163206 550350
rect 163262 550294 163358 550350
rect 162738 550226 163358 550294
rect 162738 550170 162834 550226
rect 162890 550170 162958 550226
rect 163014 550170 163082 550226
rect 163138 550170 163206 550226
rect 163262 550170 163358 550226
rect 162738 550102 163358 550170
rect 162738 550046 162834 550102
rect 162890 550046 162958 550102
rect 163014 550046 163082 550102
rect 163138 550046 163206 550102
rect 163262 550046 163358 550102
rect 162738 549978 163358 550046
rect 162738 549922 162834 549978
rect 162890 549922 162958 549978
rect 163014 549922 163082 549978
rect 163138 549922 163206 549978
rect 163262 549922 163358 549978
rect 162738 532350 163358 549922
rect 162738 532294 162834 532350
rect 162890 532294 162958 532350
rect 163014 532294 163082 532350
rect 163138 532294 163206 532350
rect 163262 532294 163358 532350
rect 162738 532226 163358 532294
rect 162738 532170 162834 532226
rect 162890 532170 162958 532226
rect 163014 532170 163082 532226
rect 163138 532170 163206 532226
rect 163262 532170 163358 532226
rect 162738 532102 163358 532170
rect 162738 532046 162834 532102
rect 162890 532046 162958 532102
rect 163014 532046 163082 532102
rect 163138 532046 163206 532102
rect 163262 532046 163358 532102
rect 162738 531978 163358 532046
rect 162738 531922 162834 531978
rect 162890 531922 162958 531978
rect 163014 531922 163082 531978
rect 163138 531922 163206 531978
rect 163262 531922 163358 531978
rect 162738 514350 163358 531922
rect 162738 514294 162834 514350
rect 162890 514294 162958 514350
rect 163014 514294 163082 514350
rect 163138 514294 163206 514350
rect 163262 514294 163358 514350
rect 162738 514226 163358 514294
rect 162738 514170 162834 514226
rect 162890 514170 162958 514226
rect 163014 514170 163082 514226
rect 163138 514170 163206 514226
rect 163262 514170 163358 514226
rect 162738 514102 163358 514170
rect 162738 514046 162834 514102
rect 162890 514046 162958 514102
rect 163014 514046 163082 514102
rect 163138 514046 163206 514102
rect 163262 514046 163358 514102
rect 162738 513978 163358 514046
rect 162738 513922 162834 513978
rect 162890 513922 162958 513978
rect 163014 513922 163082 513978
rect 163138 513922 163206 513978
rect 163262 513922 163358 513978
rect 162738 496350 163358 513922
rect 184716 565124 184772 565134
rect 162738 496294 162834 496350
rect 162890 496294 162958 496350
rect 163014 496294 163082 496350
rect 163138 496294 163206 496350
rect 163262 496294 163358 496350
rect 162738 496226 163358 496294
rect 162738 496170 162834 496226
rect 162890 496170 162958 496226
rect 163014 496170 163082 496226
rect 163138 496170 163206 496226
rect 163262 496170 163358 496226
rect 162738 496102 163358 496170
rect 162738 496046 162834 496102
rect 162890 496046 162958 496102
rect 163014 496046 163082 496102
rect 163138 496046 163206 496102
rect 163262 496046 163358 496102
rect 162738 495978 163358 496046
rect 162738 495922 162834 495978
rect 162890 495922 162958 495978
rect 163014 495922 163082 495978
rect 163138 495922 163206 495978
rect 163262 495922 163358 495978
rect 162738 478350 163358 495922
rect 162738 478294 162834 478350
rect 162890 478294 162958 478350
rect 163014 478294 163082 478350
rect 163138 478294 163206 478350
rect 163262 478294 163358 478350
rect 162738 478226 163358 478294
rect 162738 478170 162834 478226
rect 162890 478170 162958 478226
rect 163014 478170 163082 478226
rect 163138 478170 163206 478226
rect 163262 478170 163358 478226
rect 162738 478102 163358 478170
rect 162738 478046 162834 478102
rect 162890 478046 162958 478102
rect 163014 478046 163082 478102
rect 163138 478046 163206 478102
rect 163262 478046 163358 478102
rect 162738 477978 163358 478046
rect 162738 477922 162834 477978
rect 162890 477922 162958 477978
rect 163014 477922 163082 477978
rect 163138 477922 163206 477978
rect 163262 477922 163358 477978
rect 159018 454294 159114 454350
rect 159170 454294 159238 454350
rect 159294 454294 159362 454350
rect 159418 454294 159486 454350
rect 159542 454294 159638 454350
rect 159018 454226 159638 454294
rect 159018 454170 159114 454226
rect 159170 454170 159238 454226
rect 159294 454170 159362 454226
rect 159418 454170 159486 454226
rect 159542 454170 159638 454226
rect 159018 454102 159638 454170
rect 159018 454046 159114 454102
rect 159170 454046 159238 454102
rect 159294 454046 159362 454102
rect 159418 454046 159486 454102
rect 159542 454046 159638 454102
rect 159018 453978 159638 454046
rect 159018 453922 159114 453978
rect 159170 453922 159238 453978
rect 159294 453922 159362 453978
rect 159418 453922 159486 453978
rect 159542 453922 159638 453978
rect 159018 436350 159638 453922
rect 159018 436294 159114 436350
rect 159170 436294 159238 436350
rect 159294 436294 159362 436350
rect 159418 436294 159486 436350
rect 159542 436294 159638 436350
rect 159018 436226 159638 436294
rect 159018 436170 159114 436226
rect 159170 436170 159238 436226
rect 159294 436170 159362 436226
rect 159418 436170 159486 436226
rect 159542 436170 159638 436226
rect 159018 436102 159638 436170
rect 159018 436046 159114 436102
rect 159170 436046 159238 436102
rect 159294 436046 159362 436102
rect 159418 436046 159486 436102
rect 159542 436046 159638 436102
rect 159018 435978 159638 436046
rect 159018 435922 159114 435978
rect 159170 435922 159238 435978
rect 159294 435922 159362 435978
rect 159418 435922 159486 435978
rect 159542 435922 159638 435978
rect 159018 418350 159638 435922
rect 159018 418294 159114 418350
rect 159170 418294 159238 418350
rect 159294 418294 159362 418350
rect 159418 418294 159486 418350
rect 159542 418294 159638 418350
rect 159018 418226 159638 418294
rect 159018 418170 159114 418226
rect 159170 418170 159238 418226
rect 159294 418170 159362 418226
rect 159418 418170 159486 418226
rect 159542 418170 159638 418226
rect 159018 418102 159638 418170
rect 159018 418046 159114 418102
rect 159170 418046 159238 418102
rect 159294 418046 159362 418102
rect 159418 418046 159486 418102
rect 159542 418046 159638 418102
rect 159018 417978 159638 418046
rect 159018 417922 159114 417978
rect 159170 417922 159238 417978
rect 159294 417922 159362 417978
rect 159418 417922 159486 417978
rect 159542 417922 159638 417978
rect 159018 400350 159638 417922
rect 159018 400294 159114 400350
rect 159170 400294 159238 400350
rect 159294 400294 159362 400350
rect 159418 400294 159486 400350
rect 159542 400294 159638 400350
rect 159018 400226 159638 400294
rect 159018 400170 159114 400226
rect 159170 400170 159238 400226
rect 159294 400170 159362 400226
rect 159418 400170 159486 400226
rect 159542 400170 159638 400226
rect 159018 400102 159638 400170
rect 159018 400046 159114 400102
rect 159170 400046 159238 400102
rect 159294 400046 159362 400102
rect 159418 400046 159486 400102
rect 159542 400046 159638 400102
rect 159018 399978 159638 400046
rect 159018 399922 159114 399978
rect 159170 399922 159238 399978
rect 159294 399922 159362 399978
rect 159418 399922 159486 399978
rect 159542 399922 159638 399978
rect 159018 382350 159638 399922
rect 159018 382294 159114 382350
rect 159170 382294 159238 382350
rect 159294 382294 159362 382350
rect 159418 382294 159486 382350
rect 159542 382294 159638 382350
rect 159018 382226 159638 382294
rect 159018 382170 159114 382226
rect 159170 382170 159238 382226
rect 159294 382170 159362 382226
rect 159418 382170 159486 382226
rect 159542 382170 159638 382226
rect 159018 382102 159638 382170
rect 159018 382046 159114 382102
rect 159170 382046 159238 382102
rect 159294 382046 159362 382102
rect 159418 382046 159486 382102
rect 159542 382046 159638 382102
rect 159018 381978 159638 382046
rect 159018 381922 159114 381978
rect 159170 381922 159238 381978
rect 159294 381922 159362 381978
rect 159418 381922 159486 381978
rect 159542 381922 159638 381978
rect 159018 364350 159638 381922
rect 159018 364294 159114 364350
rect 159170 364294 159238 364350
rect 159294 364294 159362 364350
rect 159418 364294 159486 364350
rect 159542 364294 159638 364350
rect 159018 364226 159638 364294
rect 159018 364170 159114 364226
rect 159170 364170 159238 364226
rect 159294 364170 159362 364226
rect 159418 364170 159486 364226
rect 159542 364170 159638 364226
rect 159018 364102 159638 364170
rect 159018 364046 159114 364102
rect 159170 364046 159238 364102
rect 159294 364046 159362 364102
rect 159418 364046 159486 364102
rect 159542 364046 159638 364102
rect 159018 363978 159638 364046
rect 159018 363922 159114 363978
rect 159170 363922 159238 363978
rect 159294 363922 159362 363978
rect 159418 363922 159486 363978
rect 159542 363922 159638 363978
rect 154448 346350 154768 346384
rect 154448 346294 154518 346350
rect 154574 346294 154642 346350
rect 154698 346294 154768 346350
rect 154448 346226 154768 346294
rect 154448 346170 154518 346226
rect 154574 346170 154642 346226
rect 154698 346170 154768 346226
rect 154448 346102 154768 346170
rect 154448 346046 154518 346102
rect 154574 346046 154642 346102
rect 154698 346046 154768 346102
rect 154448 345978 154768 346046
rect 154448 345922 154518 345978
rect 154574 345922 154642 345978
rect 154698 345922 154768 345978
rect 154448 345888 154768 345922
rect 159018 346350 159638 363922
rect 159018 346294 159114 346350
rect 159170 346294 159238 346350
rect 159294 346294 159362 346350
rect 159418 346294 159486 346350
rect 159542 346294 159638 346350
rect 159018 346226 159638 346294
rect 159018 346170 159114 346226
rect 159170 346170 159238 346226
rect 159294 346170 159362 346226
rect 159418 346170 159486 346226
rect 159542 346170 159638 346226
rect 159018 346102 159638 346170
rect 159018 346046 159114 346102
rect 159170 346046 159238 346102
rect 159294 346046 159362 346102
rect 159418 346046 159486 346102
rect 159542 346046 159638 346102
rect 159018 345978 159638 346046
rect 159018 345922 159114 345978
rect 159170 345922 159238 345978
rect 159294 345922 159362 345978
rect 159418 345922 159486 345978
rect 159542 345922 159638 345978
rect 154448 328350 154768 328384
rect 154448 328294 154518 328350
rect 154574 328294 154642 328350
rect 154698 328294 154768 328350
rect 154448 328226 154768 328294
rect 154448 328170 154518 328226
rect 154574 328170 154642 328226
rect 154698 328170 154768 328226
rect 154448 328102 154768 328170
rect 154448 328046 154518 328102
rect 154574 328046 154642 328102
rect 154698 328046 154768 328102
rect 154448 327978 154768 328046
rect 154448 327922 154518 327978
rect 154574 327922 154642 327978
rect 154698 327922 154768 327978
rect 154448 327888 154768 327922
rect 159018 328350 159638 345922
rect 159018 328294 159114 328350
rect 159170 328294 159238 328350
rect 159294 328294 159362 328350
rect 159418 328294 159486 328350
rect 159542 328294 159638 328350
rect 159018 328226 159638 328294
rect 159018 328170 159114 328226
rect 159170 328170 159238 328226
rect 159294 328170 159362 328226
rect 159418 328170 159486 328226
rect 159542 328170 159638 328226
rect 159018 328102 159638 328170
rect 159018 328046 159114 328102
rect 159170 328046 159238 328102
rect 159294 328046 159362 328102
rect 159418 328046 159486 328102
rect 159542 328046 159638 328102
rect 159018 327978 159638 328046
rect 159018 327922 159114 327978
rect 159170 327922 159238 327978
rect 159294 327922 159362 327978
rect 159418 327922 159486 327978
rect 159542 327922 159638 327978
rect 146972 291218 147028 291228
rect 159018 310350 159638 327922
rect 159018 310294 159114 310350
rect 159170 310294 159238 310350
rect 159294 310294 159362 310350
rect 159418 310294 159486 310350
rect 159542 310294 159638 310350
rect 159018 310226 159638 310294
rect 159018 310170 159114 310226
rect 159170 310170 159238 310226
rect 159294 310170 159362 310226
rect 159418 310170 159486 310226
rect 159542 310170 159638 310226
rect 159018 310102 159638 310170
rect 159018 310046 159114 310102
rect 159170 310046 159238 310102
rect 159294 310046 159362 310102
rect 159418 310046 159486 310102
rect 159542 310046 159638 310102
rect 159018 309978 159638 310046
rect 159018 309922 159114 309978
rect 159170 309922 159238 309978
rect 159294 309922 159362 309978
rect 159418 309922 159486 309978
rect 159542 309922 159638 309978
rect 159018 292350 159638 309922
rect 159018 292294 159114 292350
rect 159170 292294 159238 292350
rect 159294 292294 159362 292350
rect 159418 292294 159486 292350
rect 159542 292294 159638 292350
rect 159018 292226 159638 292294
rect 159018 292170 159114 292226
rect 159170 292170 159238 292226
rect 159294 292170 159362 292226
rect 159418 292170 159486 292226
rect 159542 292170 159638 292226
rect 159018 292102 159638 292170
rect 159018 292046 159114 292102
rect 159170 292046 159238 292102
rect 159294 292046 159362 292102
rect 159418 292046 159486 292102
rect 159542 292046 159638 292102
rect 159018 291978 159638 292046
rect 159018 291922 159114 291978
rect 159170 291922 159238 291978
rect 159294 291922 159362 291978
rect 159418 291922 159486 291978
rect 159542 291922 159638 291978
rect 132018 280294 132114 280350
rect 132170 280294 132238 280350
rect 132294 280294 132362 280350
rect 132418 280294 132486 280350
rect 132542 280294 132638 280350
rect 132018 280226 132638 280294
rect 132018 280170 132114 280226
rect 132170 280170 132238 280226
rect 132294 280170 132362 280226
rect 132418 280170 132486 280226
rect 132542 280170 132638 280226
rect 132018 280102 132638 280170
rect 132018 280046 132114 280102
rect 132170 280046 132238 280102
rect 132294 280046 132362 280102
rect 132418 280046 132486 280102
rect 132542 280046 132638 280102
rect 132018 279978 132638 280046
rect 132018 279922 132114 279978
rect 132170 279922 132238 279978
rect 132294 279922 132362 279978
rect 132418 279922 132486 279978
rect 132542 279922 132638 279978
rect 132018 262350 132638 279922
rect 132018 262294 132114 262350
rect 132170 262294 132238 262350
rect 132294 262294 132362 262350
rect 132418 262294 132486 262350
rect 132542 262294 132638 262350
rect 132018 262226 132638 262294
rect 132018 262170 132114 262226
rect 132170 262170 132238 262226
rect 132294 262170 132362 262226
rect 132418 262170 132486 262226
rect 132542 262170 132638 262226
rect 132018 262102 132638 262170
rect 132018 262046 132114 262102
rect 132170 262046 132238 262102
rect 132294 262046 132362 262102
rect 132418 262046 132486 262102
rect 132542 262046 132638 262102
rect 132018 261978 132638 262046
rect 132018 261922 132114 261978
rect 132170 261922 132238 261978
rect 132294 261922 132362 261978
rect 132418 261922 132486 261978
rect 132542 261922 132638 261978
rect 132018 244350 132638 261922
rect 132018 244294 132114 244350
rect 132170 244294 132238 244350
rect 132294 244294 132362 244350
rect 132418 244294 132486 244350
rect 132542 244294 132638 244350
rect 132018 244226 132638 244294
rect 132018 244170 132114 244226
rect 132170 244170 132238 244226
rect 132294 244170 132362 244226
rect 132418 244170 132486 244226
rect 132542 244170 132638 244226
rect 132018 244102 132638 244170
rect 132018 244046 132114 244102
rect 132170 244046 132238 244102
rect 132294 244046 132362 244102
rect 132418 244046 132486 244102
rect 132542 244046 132638 244102
rect 132018 243978 132638 244046
rect 132018 243922 132114 243978
rect 132170 243922 132238 243978
rect 132294 243922 132362 243978
rect 132418 243922 132486 243978
rect 132542 243922 132638 243978
rect 132018 226350 132638 243922
rect 132018 226294 132114 226350
rect 132170 226294 132238 226350
rect 132294 226294 132362 226350
rect 132418 226294 132486 226350
rect 132542 226294 132638 226350
rect 132018 226226 132638 226294
rect 132018 226170 132114 226226
rect 132170 226170 132238 226226
rect 132294 226170 132362 226226
rect 132418 226170 132486 226226
rect 132542 226170 132638 226226
rect 132018 226102 132638 226170
rect 132018 226046 132114 226102
rect 132170 226046 132238 226102
rect 132294 226046 132362 226102
rect 132418 226046 132486 226102
rect 132542 226046 132638 226102
rect 132018 225978 132638 226046
rect 132018 225922 132114 225978
rect 132170 225922 132238 225978
rect 132294 225922 132362 225978
rect 132418 225922 132486 225978
rect 132542 225922 132638 225978
rect 132018 210462 132638 225922
rect 159018 274350 159638 291922
rect 162540 464772 162596 464782
rect 162540 286580 162596 464716
rect 162540 286514 162596 286524
rect 162738 460350 163358 477922
rect 162738 460294 162834 460350
rect 162890 460294 162958 460350
rect 163014 460294 163082 460350
rect 163138 460294 163206 460350
rect 163262 460294 163358 460350
rect 162738 460226 163358 460294
rect 162738 460170 162834 460226
rect 162890 460170 162958 460226
rect 163014 460170 163082 460226
rect 163138 460170 163206 460226
rect 163262 460170 163358 460226
rect 162738 460102 163358 460170
rect 162738 460046 162834 460102
rect 162890 460046 162958 460102
rect 163014 460046 163082 460102
rect 163138 460046 163206 460102
rect 163262 460046 163358 460102
rect 162738 459978 163358 460046
rect 162738 459922 162834 459978
rect 162890 459922 162958 459978
rect 163014 459922 163082 459978
rect 163138 459922 163206 459978
rect 163262 459922 163358 459978
rect 162738 442350 163358 459922
rect 166236 506548 166292 506558
rect 162738 442294 162834 442350
rect 162890 442294 162958 442350
rect 163014 442294 163082 442350
rect 163138 442294 163206 442350
rect 163262 442294 163358 442350
rect 162738 442226 163358 442294
rect 162738 442170 162834 442226
rect 162890 442170 162958 442226
rect 163014 442170 163082 442226
rect 163138 442170 163206 442226
rect 163262 442170 163358 442226
rect 162738 442102 163358 442170
rect 162738 442046 162834 442102
rect 162890 442046 162958 442102
rect 163014 442046 163082 442102
rect 163138 442046 163206 442102
rect 163262 442046 163358 442102
rect 162738 441978 163358 442046
rect 162738 441922 162834 441978
rect 162890 441922 162958 441978
rect 163014 441922 163082 441978
rect 163138 441922 163206 441978
rect 163262 441922 163358 441978
rect 162738 424350 163358 441922
rect 162738 424294 162834 424350
rect 162890 424294 162958 424350
rect 163014 424294 163082 424350
rect 163138 424294 163206 424350
rect 163262 424294 163358 424350
rect 162738 424226 163358 424294
rect 162738 424170 162834 424226
rect 162890 424170 162958 424226
rect 163014 424170 163082 424226
rect 163138 424170 163206 424226
rect 163262 424170 163358 424226
rect 162738 424102 163358 424170
rect 162738 424046 162834 424102
rect 162890 424046 162958 424102
rect 163014 424046 163082 424102
rect 163138 424046 163206 424102
rect 163262 424046 163358 424102
rect 162738 423978 163358 424046
rect 162738 423922 162834 423978
rect 162890 423922 162958 423978
rect 163014 423922 163082 423978
rect 163138 423922 163206 423978
rect 163262 423922 163358 423978
rect 162738 406350 163358 423922
rect 162738 406294 162834 406350
rect 162890 406294 162958 406350
rect 163014 406294 163082 406350
rect 163138 406294 163206 406350
rect 163262 406294 163358 406350
rect 162738 406226 163358 406294
rect 162738 406170 162834 406226
rect 162890 406170 162958 406226
rect 163014 406170 163082 406226
rect 163138 406170 163206 406226
rect 163262 406170 163358 406226
rect 162738 406102 163358 406170
rect 162738 406046 162834 406102
rect 162890 406046 162958 406102
rect 163014 406046 163082 406102
rect 163138 406046 163206 406102
rect 163262 406046 163358 406102
rect 162738 405978 163358 406046
rect 162738 405922 162834 405978
rect 162890 405922 162958 405978
rect 163014 405922 163082 405978
rect 163138 405922 163206 405978
rect 163262 405922 163358 405978
rect 162738 388350 163358 405922
rect 162738 388294 162834 388350
rect 162890 388294 162958 388350
rect 163014 388294 163082 388350
rect 163138 388294 163206 388350
rect 163262 388294 163358 388350
rect 162738 388226 163358 388294
rect 162738 388170 162834 388226
rect 162890 388170 162958 388226
rect 163014 388170 163082 388226
rect 163138 388170 163206 388226
rect 163262 388170 163358 388226
rect 162738 388102 163358 388170
rect 162738 388046 162834 388102
rect 162890 388046 162958 388102
rect 163014 388046 163082 388102
rect 163138 388046 163206 388102
rect 163262 388046 163358 388102
rect 162738 387978 163358 388046
rect 162738 387922 162834 387978
rect 162890 387922 162958 387978
rect 163014 387922 163082 387978
rect 163138 387922 163206 387978
rect 163262 387922 163358 387978
rect 162738 370350 163358 387922
rect 162738 370294 162834 370350
rect 162890 370294 162958 370350
rect 163014 370294 163082 370350
rect 163138 370294 163206 370350
rect 163262 370294 163358 370350
rect 162738 370226 163358 370294
rect 162738 370170 162834 370226
rect 162890 370170 162958 370226
rect 163014 370170 163082 370226
rect 163138 370170 163206 370226
rect 163262 370170 163358 370226
rect 162738 370102 163358 370170
rect 162738 370046 162834 370102
rect 162890 370046 162958 370102
rect 163014 370046 163082 370102
rect 163138 370046 163206 370102
rect 163262 370046 163358 370102
rect 162738 369978 163358 370046
rect 162738 369922 162834 369978
rect 162890 369922 162958 369978
rect 163014 369922 163082 369978
rect 163138 369922 163206 369978
rect 163262 369922 163358 369978
rect 162738 352350 163358 369922
rect 162738 352294 162834 352350
rect 162890 352294 162958 352350
rect 163014 352294 163082 352350
rect 163138 352294 163206 352350
rect 163262 352294 163358 352350
rect 162738 352226 163358 352294
rect 162738 352170 162834 352226
rect 162890 352170 162958 352226
rect 163014 352170 163082 352226
rect 163138 352170 163206 352226
rect 163262 352170 163358 352226
rect 162738 352102 163358 352170
rect 162738 352046 162834 352102
rect 162890 352046 162958 352102
rect 163014 352046 163082 352102
rect 163138 352046 163206 352102
rect 163262 352046 163358 352102
rect 162738 351978 163358 352046
rect 162738 351922 162834 351978
rect 162890 351922 162958 351978
rect 163014 351922 163082 351978
rect 163138 351922 163206 351978
rect 163262 351922 163358 351978
rect 162738 334350 163358 351922
rect 162738 334294 162834 334350
rect 162890 334294 162958 334350
rect 163014 334294 163082 334350
rect 163138 334294 163206 334350
rect 163262 334294 163358 334350
rect 162738 334226 163358 334294
rect 162738 334170 162834 334226
rect 162890 334170 162958 334226
rect 163014 334170 163082 334226
rect 163138 334170 163206 334226
rect 163262 334170 163358 334226
rect 162738 334102 163358 334170
rect 162738 334046 162834 334102
rect 162890 334046 162958 334102
rect 163014 334046 163082 334102
rect 163138 334046 163206 334102
rect 163262 334046 163358 334102
rect 162738 333978 163358 334046
rect 162738 333922 162834 333978
rect 162890 333922 162958 333978
rect 163014 333922 163082 333978
rect 163138 333922 163206 333978
rect 163262 333922 163358 333978
rect 162738 316350 163358 333922
rect 162738 316294 162834 316350
rect 162890 316294 162958 316350
rect 163014 316294 163082 316350
rect 163138 316294 163206 316350
rect 163262 316294 163358 316350
rect 162738 316226 163358 316294
rect 162738 316170 162834 316226
rect 162890 316170 162958 316226
rect 163014 316170 163082 316226
rect 163138 316170 163206 316226
rect 163262 316170 163358 316226
rect 162738 316102 163358 316170
rect 162738 316046 162834 316102
rect 162890 316046 162958 316102
rect 163014 316046 163082 316102
rect 163138 316046 163206 316102
rect 163262 316046 163358 316102
rect 162738 315978 163358 316046
rect 162738 315922 162834 315978
rect 162890 315922 162958 315978
rect 163014 315922 163082 315978
rect 163138 315922 163206 315978
rect 163262 315922 163358 315978
rect 162738 298350 163358 315922
rect 162738 298294 162834 298350
rect 162890 298294 162958 298350
rect 163014 298294 163082 298350
rect 163138 298294 163206 298350
rect 163262 298294 163358 298350
rect 162738 298226 163358 298294
rect 162738 298170 162834 298226
rect 162890 298170 162958 298226
rect 163014 298170 163082 298226
rect 163138 298170 163206 298226
rect 163262 298170 163358 298226
rect 162738 298102 163358 298170
rect 162738 298046 162834 298102
rect 162890 298046 162958 298102
rect 163014 298046 163082 298102
rect 163138 298046 163206 298102
rect 163262 298046 163358 298102
rect 162738 297978 163358 298046
rect 162738 297922 162834 297978
rect 162890 297922 162958 297978
rect 163014 297922 163082 297978
rect 163138 297922 163206 297978
rect 163262 297922 163358 297978
rect 159018 274294 159114 274350
rect 159170 274294 159238 274350
rect 159294 274294 159362 274350
rect 159418 274294 159486 274350
rect 159542 274294 159638 274350
rect 159018 274226 159638 274294
rect 159018 274170 159114 274226
rect 159170 274170 159238 274226
rect 159294 274170 159362 274226
rect 159418 274170 159486 274226
rect 159542 274170 159638 274226
rect 159018 274102 159638 274170
rect 159018 274046 159114 274102
rect 159170 274046 159238 274102
rect 159294 274046 159362 274102
rect 159418 274046 159486 274102
rect 159542 274046 159638 274102
rect 159018 273978 159638 274046
rect 159018 273922 159114 273978
rect 159170 273922 159238 273978
rect 159294 273922 159362 273978
rect 159418 273922 159486 273978
rect 159542 273922 159638 273978
rect 159018 256350 159638 273922
rect 159018 256294 159114 256350
rect 159170 256294 159238 256350
rect 159294 256294 159362 256350
rect 159418 256294 159486 256350
rect 159542 256294 159638 256350
rect 159018 256226 159638 256294
rect 159018 256170 159114 256226
rect 159170 256170 159238 256226
rect 159294 256170 159362 256226
rect 159418 256170 159486 256226
rect 159542 256170 159638 256226
rect 159018 256102 159638 256170
rect 159018 256046 159114 256102
rect 159170 256046 159238 256102
rect 159294 256046 159362 256102
rect 159418 256046 159486 256102
rect 159542 256046 159638 256102
rect 159018 255978 159638 256046
rect 159018 255922 159114 255978
rect 159170 255922 159238 255978
rect 159294 255922 159362 255978
rect 159418 255922 159486 255978
rect 159542 255922 159638 255978
rect 159018 238350 159638 255922
rect 159018 238294 159114 238350
rect 159170 238294 159238 238350
rect 159294 238294 159362 238350
rect 159418 238294 159486 238350
rect 159542 238294 159638 238350
rect 159018 238226 159638 238294
rect 159018 238170 159114 238226
rect 159170 238170 159238 238226
rect 159294 238170 159362 238226
rect 159418 238170 159486 238226
rect 159542 238170 159638 238226
rect 159018 238102 159638 238170
rect 159018 238046 159114 238102
rect 159170 238046 159238 238102
rect 159294 238046 159362 238102
rect 159418 238046 159486 238102
rect 159542 238046 159638 238102
rect 159018 237978 159638 238046
rect 159018 237922 159114 237978
rect 159170 237922 159238 237978
rect 159294 237922 159362 237978
rect 159418 237922 159486 237978
rect 159542 237922 159638 237978
rect 159018 220350 159638 237922
rect 159018 220294 159114 220350
rect 159170 220294 159238 220350
rect 159294 220294 159362 220350
rect 159418 220294 159486 220350
rect 159542 220294 159638 220350
rect 159018 220226 159638 220294
rect 159018 220170 159114 220226
rect 159170 220170 159238 220226
rect 159294 220170 159362 220226
rect 159418 220170 159486 220226
rect 159542 220170 159638 220226
rect 159018 220102 159638 220170
rect 159018 220046 159114 220102
rect 159170 220046 159238 220102
rect 159294 220046 159362 220102
rect 159418 220046 159486 220102
rect 159542 220046 159638 220102
rect 159018 219978 159638 220046
rect 159018 219922 159114 219978
rect 159170 219922 159238 219978
rect 159294 219922 159362 219978
rect 159418 219922 159486 219978
rect 159542 219922 159638 219978
rect 159018 210462 159638 219922
rect 162738 280350 163358 297922
rect 166124 450436 166180 450446
rect 166124 285460 166180 450380
rect 166124 285394 166180 285404
rect 166236 284228 166292 506492
rect 167916 500612 167972 500622
rect 167804 443268 167860 443278
rect 167804 286692 167860 443212
rect 167804 286626 167860 286636
rect 167916 285572 167972 500556
rect 184716 397908 184772 565068
rect 189738 562350 190358 579922
rect 189738 562294 189834 562350
rect 189890 562294 189958 562350
rect 190014 562294 190082 562350
rect 190138 562294 190206 562350
rect 190262 562294 190358 562350
rect 189738 562226 190358 562294
rect 189738 562170 189834 562226
rect 189890 562170 189958 562226
rect 190014 562170 190082 562226
rect 190138 562170 190206 562226
rect 190262 562170 190358 562226
rect 189738 562102 190358 562170
rect 189738 562046 189834 562102
rect 189890 562046 189958 562102
rect 190014 562046 190082 562102
rect 190138 562046 190206 562102
rect 190262 562046 190358 562102
rect 189738 561978 190358 562046
rect 189738 561922 189834 561978
rect 189890 561922 189958 561978
rect 190014 561922 190082 561978
rect 190138 561922 190206 561978
rect 190262 561922 190358 561978
rect 187852 557956 187908 557966
rect 186396 550788 186452 550798
rect 186284 536452 186340 536462
rect 184716 397842 184772 397852
rect 186172 514948 186228 514958
rect 186172 396228 186228 514892
rect 186284 405972 186340 536396
rect 186284 405906 186340 405916
rect 186396 399364 186452 550732
rect 187516 543620 187572 543630
rect 187404 507780 187460 507790
rect 187404 506548 187460 507724
rect 187404 506482 187460 506492
rect 186396 399298 186452 399308
rect 187292 436100 187348 436110
rect 186172 396162 186228 396172
rect 169808 352350 170128 352384
rect 169808 352294 169878 352350
rect 169934 352294 170002 352350
rect 170058 352294 170128 352350
rect 169808 352226 170128 352294
rect 169808 352170 169878 352226
rect 169934 352170 170002 352226
rect 170058 352170 170128 352226
rect 169808 352102 170128 352170
rect 169808 352046 169878 352102
rect 169934 352046 170002 352102
rect 170058 352046 170128 352102
rect 169808 351978 170128 352046
rect 169808 351922 169878 351978
rect 169934 351922 170002 351978
rect 170058 351922 170128 351978
rect 169808 351888 170128 351922
rect 185168 346350 185488 346384
rect 185168 346294 185238 346350
rect 185294 346294 185362 346350
rect 185418 346294 185488 346350
rect 185168 346226 185488 346294
rect 185168 346170 185238 346226
rect 185294 346170 185362 346226
rect 185418 346170 185488 346226
rect 185168 346102 185488 346170
rect 185168 346046 185238 346102
rect 185294 346046 185362 346102
rect 185418 346046 185488 346102
rect 185168 345978 185488 346046
rect 185168 345922 185238 345978
rect 185294 345922 185362 345978
rect 185418 345922 185488 345978
rect 185168 345888 185488 345922
rect 169808 334350 170128 334384
rect 169808 334294 169878 334350
rect 169934 334294 170002 334350
rect 170058 334294 170128 334350
rect 169808 334226 170128 334294
rect 169808 334170 169878 334226
rect 169934 334170 170002 334226
rect 170058 334170 170128 334226
rect 169808 334102 170128 334170
rect 169808 334046 169878 334102
rect 169934 334046 170002 334102
rect 170058 334046 170128 334102
rect 169808 333978 170128 334046
rect 169808 333922 169878 333978
rect 169934 333922 170002 333978
rect 170058 333922 170128 333978
rect 169808 333888 170128 333922
rect 185168 328350 185488 328384
rect 185168 328294 185238 328350
rect 185294 328294 185362 328350
rect 185418 328294 185488 328350
rect 185168 328226 185488 328294
rect 185168 328170 185238 328226
rect 185294 328170 185362 328226
rect 185418 328170 185488 328226
rect 185168 328102 185488 328170
rect 185168 328046 185238 328102
rect 185294 328046 185362 328102
rect 185418 328046 185488 328102
rect 185168 327978 185488 328046
rect 185168 327922 185238 327978
rect 185294 327922 185362 327978
rect 185418 327922 185488 327978
rect 185168 327888 185488 327922
rect 167916 285506 167972 285516
rect 186508 296100 186564 296110
rect 166236 284162 166292 284172
rect 162738 280294 162834 280350
rect 162890 280294 162958 280350
rect 163014 280294 163082 280350
rect 163138 280294 163206 280350
rect 163262 280294 163358 280350
rect 162738 280226 163358 280294
rect 162738 280170 162834 280226
rect 162890 280170 162958 280226
rect 163014 280170 163082 280226
rect 163138 280170 163206 280226
rect 163262 280170 163358 280226
rect 162738 280102 163358 280170
rect 162738 280046 162834 280102
rect 162890 280046 162958 280102
rect 163014 280046 163082 280102
rect 163138 280046 163206 280102
rect 163262 280046 163358 280102
rect 162738 279978 163358 280046
rect 162738 279922 162834 279978
rect 162890 279922 162958 279978
rect 163014 279922 163082 279978
rect 163138 279922 163206 279978
rect 163262 279922 163358 279978
rect 162738 262350 163358 279922
rect 167008 280350 167328 280384
rect 167008 280294 167078 280350
rect 167134 280294 167202 280350
rect 167258 280294 167328 280350
rect 167008 280226 167328 280294
rect 167008 280170 167078 280226
rect 167134 280170 167202 280226
rect 167258 280170 167328 280226
rect 167008 280102 167328 280170
rect 167008 280046 167078 280102
rect 167134 280046 167202 280102
rect 167258 280046 167328 280102
rect 167008 279978 167328 280046
rect 167008 279922 167078 279978
rect 167134 279922 167202 279978
rect 167258 279922 167328 279978
rect 167008 279888 167328 279922
rect 172832 280350 173152 280384
rect 172832 280294 172902 280350
rect 172958 280294 173026 280350
rect 173082 280294 173152 280350
rect 172832 280226 173152 280294
rect 172832 280170 172902 280226
rect 172958 280170 173026 280226
rect 173082 280170 173152 280226
rect 172832 280102 173152 280170
rect 172832 280046 172902 280102
rect 172958 280046 173026 280102
rect 173082 280046 173152 280102
rect 172832 279978 173152 280046
rect 172832 279922 172902 279978
rect 172958 279922 173026 279978
rect 173082 279922 173152 279978
rect 172832 279888 173152 279922
rect 178656 280350 178976 280384
rect 178656 280294 178726 280350
rect 178782 280294 178850 280350
rect 178906 280294 178976 280350
rect 178656 280226 178976 280294
rect 178656 280170 178726 280226
rect 178782 280170 178850 280226
rect 178906 280170 178976 280226
rect 178656 280102 178976 280170
rect 178656 280046 178726 280102
rect 178782 280046 178850 280102
rect 178906 280046 178976 280102
rect 178656 279978 178976 280046
rect 178656 279922 178726 279978
rect 178782 279922 178850 279978
rect 178906 279922 178976 279978
rect 178656 279888 178976 279922
rect 184480 280350 184800 280384
rect 184480 280294 184550 280350
rect 184606 280294 184674 280350
rect 184730 280294 184800 280350
rect 184480 280226 184800 280294
rect 184480 280170 184550 280226
rect 184606 280170 184674 280226
rect 184730 280170 184800 280226
rect 184480 280102 184800 280170
rect 184480 280046 184550 280102
rect 184606 280046 184674 280102
rect 184730 280046 184800 280102
rect 184480 279978 184800 280046
rect 184480 279922 184550 279978
rect 184606 279922 184674 279978
rect 184730 279922 184800 279978
rect 184480 279888 184800 279922
rect 164096 274350 164416 274384
rect 164096 274294 164166 274350
rect 164222 274294 164290 274350
rect 164346 274294 164416 274350
rect 164096 274226 164416 274294
rect 164096 274170 164166 274226
rect 164222 274170 164290 274226
rect 164346 274170 164416 274226
rect 164096 274102 164416 274170
rect 164096 274046 164166 274102
rect 164222 274046 164290 274102
rect 164346 274046 164416 274102
rect 164096 273978 164416 274046
rect 164096 273922 164166 273978
rect 164222 273922 164290 273978
rect 164346 273922 164416 273978
rect 164096 273888 164416 273922
rect 169920 274350 170240 274384
rect 169920 274294 169990 274350
rect 170046 274294 170114 274350
rect 170170 274294 170240 274350
rect 169920 274226 170240 274294
rect 169920 274170 169990 274226
rect 170046 274170 170114 274226
rect 170170 274170 170240 274226
rect 169920 274102 170240 274170
rect 169920 274046 169990 274102
rect 170046 274046 170114 274102
rect 170170 274046 170240 274102
rect 169920 273978 170240 274046
rect 169920 273922 169990 273978
rect 170046 273922 170114 273978
rect 170170 273922 170240 273978
rect 169920 273888 170240 273922
rect 175744 274350 176064 274384
rect 175744 274294 175814 274350
rect 175870 274294 175938 274350
rect 175994 274294 176064 274350
rect 175744 274226 176064 274294
rect 175744 274170 175814 274226
rect 175870 274170 175938 274226
rect 175994 274170 176064 274226
rect 175744 274102 176064 274170
rect 175744 274046 175814 274102
rect 175870 274046 175938 274102
rect 175994 274046 176064 274102
rect 175744 273978 176064 274046
rect 175744 273922 175814 273978
rect 175870 273922 175938 273978
rect 175994 273922 176064 273978
rect 175744 273888 176064 273922
rect 181568 274350 181888 274384
rect 181568 274294 181638 274350
rect 181694 274294 181762 274350
rect 181818 274294 181888 274350
rect 181568 274226 181888 274294
rect 181568 274170 181638 274226
rect 181694 274170 181762 274226
rect 181818 274170 181888 274226
rect 181568 274102 181888 274170
rect 181568 274046 181638 274102
rect 181694 274046 181762 274102
rect 181818 274046 181888 274102
rect 181568 273978 181888 274046
rect 181568 273922 181638 273978
rect 181694 273922 181762 273978
rect 181818 273922 181888 273978
rect 181568 273888 181888 273922
rect 186508 264628 186564 296044
rect 187292 296100 187348 436044
rect 187292 296034 187348 296044
rect 187404 428932 187460 428942
rect 187404 290276 187460 428876
rect 187516 404292 187572 543564
rect 187740 529284 187796 529294
rect 187628 522116 187684 522126
rect 187628 408996 187684 522060
rect 187628 408930 187684 408940
rect 187516 404226 187572 404236
rect 187740 396340 187796 529228
rect 187852 402836 187908 557900
rect 189738 544350 190358 561922
rect 189738 544294 189834 544350
rect 189890 544294 189958 544350
rect 190014 544294 190082 544350
rect 190138 544294 190206 544350
rect 190262 544294 190358 544350
rect 189738 544226 190358 544294
rect 189738 544170 189834 544226
rect 189890 544170 189958 544226
rect 190014 544170 190082 544226
rect 190138 544170 190206 544226
rect 190262 544170 190358 544226
rect 189738 544102 190358 544170
rect 189738 544046 189834 544102
rect 189890 544046 189958 544102
rect 190014 544046 190082 544102
rect 190138 544046 190206 544102
rect 190262 544046 190358 544102
rect 189738 543978 190358 544046
rect 189738 543922 189834 543978
rect 189890 543922 189958 543978
rect 190014 543922 190082 543978
rect 190138 543922 190206 543978
rect 190262 543922 190358 543978
rect 189738 526350 190358 543922
rect 189738 526294 189834 526350
rect 189890 526294 189958 526350
rect 190014 526294 190082 526350
rect 190138 526294 190206 526350
rect 190262 526294 190358 526350
rect 189738 526226 190358 526294
rect 189738 526170 189834 526226
rect 189890 526170 189958 526226
rect 190014 526170 190082 526226
rect 190138 526170 190206 526226
rect 190262 526170 190358 526226
rect 189738 526102 190358 526170
rect 189738 526046 189834 526102
rect 189890 526046 189958 526102
rect 190014 526046 190082 526102
rect 190138 526046 190206 526102
rect 190262 526046 190358 526102
rect 189738 525978 190358 526046
rect 189738 525922 189834 525978
rect 189890 525922 189958 525978
rect 190014 525922 190082 525978
rect 190138 525922 190206 525978
rect 190262 525922 190358 525978
rect 189738 508350 190358 525922
rect 189738 508294 189834 508350
rect 189890 508294 189958 508350
rect 190014 508294 190082 508350
rect 190138 508294 190206 508350
rect 190262 508294 190358 508350
rect 189738 508226 190358 508294
rect 189738 508170 189834 508226
rect 189890 508170 189958 508226
rect 190014 508170 190082 508226
rect 190138 508170 190206 508226
rect 190262 508170 190358 508226
rect 189738 508102 190358 508170
rect 189738 508046 189834 508102
rect 189890 508046 189958 508102
rect 190014 508046 190082 508102
rect 190138 508046 190206 508102
rect 190262 508046 190358 508102
rect 189738 507978 190358 508046
rect 189738 507922 189834 507978
rect 189890 507922 189958 507978
rect 190014 507922 190082 507978
rect 190138 507922 190206 507978
rect 190262 507922 190358 507978
rect 188972 493444 189028 493454
rect 187964 471940 188020 471950
rect 187964 462178 188020 471884
rect 187964 462122 188244 462178
rect 187852 402770 187908 402780
rect 187964 457604 188020 457614
rect 187740 396274 187796 396284
rect 186508 264562 186564 264572
rect 186620 289044 186676 289054
rect 162738 262294 162834 262350
rect 162890 262294 162958 262350
rect 163014 262294 163082 262350
rect 163138 262294 163206 262350
rect 163262 262294 163358 262350
rect 162738 262226 163358 262294
rect 162738 262170 162834 262226
rect 162890 262170 162958 262226
rect 163014 262170 163082 262226
rect 163138 262170 163206 262226
rect 163262 262170 163358 262226
rect 162738 262102 163358 262170
rect 162738 262046 162834 262102
rect 162890 262046 162958 262102
rect 163014 262046 163082 262102
rect 163138 262046 163206 262102
rect 163262 262046 163358 262102
rect 162738 261978 163358 262046
rect 162738 261922 162834 261978
rect 162890 261922 162958 261978
rect 163014 261922 163082 261978
rect 163138 261922 163206 261978
rect 163262 261922 163358 261978
rect 162738 244350 163358 261922
rect 186620 261828 186676 288988
rect 187404 289044 187460 290220
rect 187404 288978 187460 288988
rect 187964 269892 188020 457548
rect 188188 455308 188244 462122
rect 188188 455252 188692 455308
rect 188076 414596 188132 414606
rect 188076 290612 188132 414540
rect 188076 289044 188132 290556
rect 188076 288978 188132 288988
rect 188300 286692 188356 286702
rect 188188 285572 188244 285582
rect 188188 281428 188244 285516
rect 188188 281362 188244 281372
rect 187964 269826 188020 269836
rect 188300 266308 188356 286636
rect 188524 286580 188580 286590
rect 188412 285460 188468 285470
rect 188412 267988 188468 285404
rect 188524 271348 188580 286524
rect 188636 273924 188692 455252
rect 188636 273858 188692 273868
rect 188972 279972 189028 493388
rect 189738 490350 190358 507922
rect 189738 490294 189834 490350
rect 189890 490294 189958 490350
rect 190014 490294 190082 490350
rect 190138 490294 190206 490350
rect 190262 490294 190358 490350
rect 189738 490226 190358 490294
rect 189738 490170 189834 490226
rect 189890 490170 189958 490226
rect 190014 490170 190082 490226
rect 190138 490170 190206 490226
rect 190262 490170 190358 490226
rect 189738 490102 190358 490170
rect 189738 490046 189834 490102
rect 189890 490046 189958 490102
rect 190014 490046 190082 490102
rect 190138 490046 190206 490102
rect 190262 490046 190358 490102
rect 189738 489978 190358 490046
rect 189738 489922 189834 489978
rect 189890 489922 189958 489978
rect 190014 489922 190082 489978
rect 190138 489922 190206 489978
rect 190262 489922 190358 489978
rect 189532 486276 189588 486286
rect 189420 479108 189476 479118
rect 189308 421764 189364 421774
rect 189308 396452 189364 421708
rect 189308 396386 189364 396396
rect 188524 271282 188580 271292
rect 188412 267922 188468 267932
rect 188300 266242 188356 266252
rect 186620 261762 186676 261772
rect 188972 246820 189028 279916
rect 189420 276388 189476 479052
rect 189532 278068 189588 486220
rect 189532 278002 189588 278012
rect 189738 472350 190358 489922
rect 189738 472294 189834 472350
rect 189890 472294 189958 472350
rect 190014 472294 190082 472350
rect 190138 472294 190206 472350
rect 190262 472294 190358 472350
rect 189738 472226 190358 472294
rect 189738 472170 189834 472226
rect 189890 472170 189958 472226
rect 190014 472170 190082 472226
rect 190138 472170 190206 472226
rect 190262 472170 190358 472226
rect 189738 472102 190358 472170
rect 189738 472046 189834 472102
rect 189890 472046 189958 472102
rect 190014 472046 190082 472102
rect 190138 472046 190206 472102
rect 190262 472046 190358 472102
rect 189738 471978 190358 472046
rect 189738 471922 189834 471978
rect 189890 471922 189958 471978
rect 190014 471922 190082 471978
rect 190138 471922 190206 471978
rect 190262 471922 190358 471978
rect 189738 454350 190358 471922
rect 189738 454294 189834 454350
rect 189890 454294 189958 454350
rect 190014 454294 190082 454350
rect 190138 454294 190206 454350
rect 190262 454294 190358 454350
rect 189738 454226 190358 454294
rect 189738 454170 189834 454226
rect 189890 454170 189958 454226
rect 190014 454170 190082 454226
rect 190138 454170 190206 454226
rect 190262 454170 190358 454226
rect 189738 454102 190358 454170
rect 189738 454046 189834 454102
rect 189890 454046 189958 454102
rect 190014 454046 190082 454102
rect 190138 454046 190206 454102
rect 190262 454046 190358 454102
rect 189738 453978 190358 454046
rect 189738 453922 189834 453978
rect 189890 453922 189958 453978
rect 190014 453922 190082 453978
rect 190138 453922 190206 453978
rect 190262 453922 190358 453978
rect 189738 436350 190358 453922
rect 189738 436294 189834 436350
rect 189890 436294 189958 436350
rect 190014 436294 190082 436350
rect 190138 436294 190206 436350
rect 190262 436294 190358 436350
rect 189738 436226 190358 436294
rect 189738 436170 189834 436226
rect 189890 436170 189958 436226
rect 190014 436170 190082 436226
rect 190138 436170 190206 436226
rect 190262 436170 190358 436226
rect 189738 436102 190358 436170
rect 189738 436046 189834 436102
rect 189890 436046 189958 436102
rect 190014 436046 190082 436102
rect 190138 436046 190206 436102
rect 190262 436046 190358 436102
rect 189738 435978 190358 436046
rect 189738 435922 189834 435978
rect 189890 435922 189958 435978
rect 190014 435922 190082 435978
rect 190138 435922 190206 435978
rect 190262 435922 190358 435978
rect 189738 418350 190358 435922
rect 189738 418294 189834 418350
rect 189890 418294 189958 418350
rect 190014 418294 190082 418350
rect 190138 418294 190206 418350
rect 190262 418294 190358 418350
rect 189738 418226 190358 418294
rect 189738 418170 189834 418226
rect 189890 418170 189958 418226
rect 190014 418170 190082 418226
rect 190138 418170 190206 418226
rect 190262 418170 190358 418226
rect 189738 418102 190358 418170
rect 189738 418046 189834 418102
rect 189890 418046 189958 418102
rect 190014 418046 190082 418102
rect 190138 418046 190206 418102
rect 190262 418046 190358 418102
rect 189738 417978 190358 418046
rect 189738 417922 189834 417978
rect 189890 417922 189958 417978
rect 190014 417922 190082 417978
rect 190138 417922 190206 417978
rect 190262 417922 190358 417978
rect 189738 400350 190358 417922
rect 190428 591332 190484 591342
rect 190428 404068 190484 591276
rect 192780 591108 192836 591118
rect 190540 590660 190596 590670
rect 190540 406532 190596 590604
rect 192668 590548 192724 590558
rect 190540 406466 190596 406476
rect 190652 589978 190708 589988
rect 190428 404002 190484 404012
rect 189738 400294 189834 400350
rect 189890 400294 189958 400350
rect 190014 400294 190082 400350
rect 190138 400294 190206 400350
rect 190262 400294 190358 400350
rect 189738 400226 190358 400294
rect 189738 400170 189834 400226
rect 189890 400170 189958 400226
rect 190014 400170 190082 400226
rect 190138 400170 190206 400226
rect 190262 400170 190358 400226
rect 189738 400102 190358 400170
rect 189738 400046 189834 400102
rect 189890 400046 189958 400102
rect 190014 400046 190082 400102
rect 190138 400046 190206 400102
rect 190262 400046 190358 400102
rect 189738 399978 190358 400046
rect 189738 399922 189834 399978
rect 189890 399922 189958 399978
rect 190014 399922 190082 399978
rect 190138 399922 190206 399978
rect 190262 399922 190358 399978
rect 189738 382350 190358 399922
rect 189738 382294 189834 382350
rect 189890 382294 189958 382350
rect 190014 382294 190082 382350
rect 190138 382294 190206 382350
rect 190262 382294 190358 382350
rect 189738 382226 190358 382294
rect 189738 382170 189834 382226
rect 189890 382170 189958 382226
rect 190014 382170 190082 382226
rect 190138 382170 190206 382226
rect 190262 382170 190358 382226
rect 189738 382102 190358 382170
rect 189738 382046 189834 382102
rect 189890 382046 189958 382102
rect 190014 382046 190082 382102
rect 190138 382046 190206 382102
rect 190262 382046 190358 382102
rect 189738 381978 190358 382046
rect 189738 381922 189834 381978
rect 189890 381922 189958 381978
rect 190014 381922 190082 381978
rect 190138 381922 190206 381978
rect 190262 381922 190358 381978
rect 189738 364350 190358 381922
rect 189738 364294 189834 364350
rect 189890 364294 189958 364350
rect 190014 364294 190082 364350
rect 190138 364294 190206 364350
rect 190262 364294 190358 364350
rect 189738 364226 190358 364294
rect 189738 364170 189834 364226
rect 189890 364170 189958 364226
rect 190014 364170 190082 364226
rect 190138 364170 190206 364226
rect 190262 364170 190358 364226
rect 189738 364102 190358 364170
rect 189738 364046 189834 364102
rect 189890 364046 189958 364102
rect 190014 364046 190082 364102
rect 190138 364046 190206 364102
rect 190262 364046 190358 364102
rect 189738 363978 190358 364046
rect 189738 363922 189834 363978
rect 189890 363922 189958 363978
rect 190014 363922 190082 363978
rect 190138 363922 190206 363978
rect 190262 363922 190358 363978
rect 189738 346350 190358 363922
rect 189738 346294 189834 346350
rect 189890 346294 189958 346350
rect 190014 346294 190082 346350
rect 190138 346294 190206 346350
rect 190262 346294 190358 346350
rect 189738 346226 190358 346294
rect 189738 346170 189834 346226
rect 189890 346170 189958 346226
rect 190014 346170 190082 346226
rect 190138 346170 190206 346226
rect 190262 346170 190358 346226
rect 189738 346102 190358 346170
rect 189738 346046 189834 346102
rect 189890 346046 189958 346102
rect 190014 346046 190082 346102
rect 190138 346046 190206 346102
rect 190262 346046 190358 346102
rect 189738 345978 190358 346046
rect 189738 345922 189834 345978
rect 189890 345922 189958 345978
rect 190014 345922 190082 345978
rect 190138 345922 190206 345978
rect 190262 345922 190358 345978
rect 189738 328350 190358 345922
rect 189738 328294 189834 328350
rect 189890 328294 189958 328350
rect 190014 328294 190082 328350
rect 190138 328294 190206 328350
rect 190262 328294 190358 328350
rect 189738 328226 190358 328294
rect 189738 328170 189834 328226
rect 189890 328170 189958 328226
rect 190014 328170 190082 328226
rect 190138 328170 190206 328226
rect 190262 328170 190358 328226
rect 189738 328102 190358 328170
rect 189738 328046 189834 328102
rect 189890 328046 189958 328102
rect 190014 328046 190082 328102
rect 190138 328046 190206 328102
rect 190262 328046 190358 328102
rect 189738 327978 190358 328046
rect 189738 327922 189834 327978
rect 189890 327922 189958 327978
rect 190014 327922 190082 327978
rect 190138 327922 190206 327978
rect 190262 327922 190358 327978
rect 189738 310350 190358 327922
rect 189738 310294 189834 310350
rect 189890 310294 189958 310350
rect 190014 310294 190082 310350
rect 190138 310294 190206 310350
rect 190262 310294 190358 310350
rect 189738 310226 190358 310294
rect 189738 310170 189834 310226
rect 189890 310170 189958 310226
rect 190014 310170 190082 310226
rect 190138 310170 190206 310226
rect 190262 310170 190358 310226
rect 189738 310102 190358 310170
rect 189738 310046 189834 310102
rect 189890 310046 189958 310102
rect 190014 310046 190082 310102
rect 190138 310046 190206 310102
rect 190262 310046 190358 310102
rect 189738 309978 190358 310046
rect 189738 309922 189834 309978
rect 189890 309922 189958 309978
rect 190014 309922 190082 309978
rect 190138 309922 190206 309978
rect 190262 309922 190358 309978
rect 189738 292350 190358 309922
rect 189738 292294 189834 292350
rect 189890 292294 189958 292350
rect 190014 292294 190082 292350
rect 190138 292294 190206 292350
rect 190262 292294 190358 292350
rect 189738 292226 190358 292294
rect 189738 292170 189834 292226
rect 189890 292170 189958 292226
rect 190014 292170 190082 292226
rect 190138 292170 190206 292226
rect 190262 292170 190358 292226
rect 189738 292102 190358 292170
rect 189738 292046 189834 292102
rect 189890 292046 189958 292102
rect 190014 292046 190082 292102
rect 190138 292046 190206 292102
rect 190262 292046 190358 292102
rect 189738 291978 190358 292046
rect 189738 291922 189834 291978
rect 189890 291922 189958 291978
rect 190014 291922 190082 291978
rect 190138 291922 190206 291978
rect 190262 291922 190358 291978
rect 189420 276322 189476 276332
rect 189738 274350 190358 291922
rect 190652 283444 190708 589922
rect 192668 409444 192724 590492
rect 192668 409378 192724 409388
rect 192780 409332 192836 591052
rect 193004 590884 193060 590894
rect 192780 409266 192836 409276
rect 192892 590436 192948 590446
rect 192892 286804 192948 590380
rect 192892 286738 192948 286748
rect 193004 284564 193060 590828
rect 193004 284498 193060 284508
rect 193116 589798 193172 589808
rect 190652 283378 190708 283388
rect 193116 282324 193172 589742
rect 193458 586350 194078 597744
rect 193458 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 194078 586350
rect 193458 586226 194078 586294
rect 193458 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 194078 586226
rect 193458 586102 194078 586170
rect 193458 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 194078 586102
rect 193458 585978 194078 586046
rect 193458 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 194078 585978
rect 193458 569342 194078 585922
rect 220458 597212 221078 598268
rect 220458 597156 220554 597212
rect 220610 597156 220678 597212
rect 220734 597156 220802 597212
rect 220858 597156 220926 597212
rect 220982 597156 221078 597212
rect 220458 597088 221078 597156
rect 220458 597032 220554 597088
rect 220610 597032 220678 597088
rect 220734 597032 220802 597088
rect 220858 597032 220926 597088
rect 220982 597032 221078 597088
rect 220458 596964 221078 597032
rect 220458 596908 220554 596964
rect 220610 596908 220678 596964
rect 220734 596908 220802 596964
rect 220858 596908 220926 596964
rect 220982 596908 221078 596964
rect 220458 596840 221078 596908
rect 220458 596784 220554 596840
rect 220610 596784 220678 596840
rect 220734 596784 220802 596840
rect 220858 596784 220926 596840
rect 220982 596784 221078 596840
rect 220458 580350 221078 596784
rect 220458 580294 220554 580350
rect 220610 580294 220678 580350
rect 220734 580294 220802 580350
rect 220858 580294 220926 580350
rect 220982 580294 221078 580350
rect 220458 580226 221078 580294
rect 220458 580170 220554 580226
rect 220610 580170 220678 580226
rect 220734 580170 220802 580226
rect 220858 580170 220926 580226
rect 220982 580170 221078 580226
rect 220458 580102 221078 580170
rect 220458 580046 220554 580102
rect 220610 580046 220678 580102
rect 220734 580046 220802 580102
rect 220858 580046 220926 580102
rect 220982 580046 221078 580102
rect 220458 579978 221078 580046
rect 220458 579922 220554 579978
rect 220610 579922 220678 579978
rect 220734 579922 220802 579978
rect 220858 579922 220926 579978
rect 220982 579922 221078 579978
rect 220458 569342 221078 579922
rect 224178 598172 224798 598268
rect 224178 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 224798 598172
rect 224178 598048 224798 598116
rect 224178 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 224798 598048
rect 224178 597924 224798 597992
rect 224178 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 224798 597924
rect 224178 597800 224798 597868
rect 224178 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 224798 597800
rect 224178 586350 224798 597744
rect 224178 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 224798 586350
rect 224178 586226 224798 586294
rect 224178 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 224798 586226
rect 224178 586102 224798 586170
rect 224178 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 224798 586102
rect 224178 585978 224798 586046
rect 224178 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 224798 585978
rect 224178 569342 224798 585922
rect 251178 597212 251798 598268
rect 251178 597156 251274 597212
rect 251330 597156 251398 597212
rect 251454 597156 251522 597212
rect 251578 597156 251646 597212
rect 251702 597156 251798 597212
rect 251178 597088 251798 597156
rect 251178 597032 251274 597088
rect 251330 597032 251398 597088
rect 251454 597032 251522 597088
rect 251578 597032 251646 597088
rect 251702 597032 251798 597088
rect 251178 596964 251798 597032
rect 251178 596908 251274 596964
rect 251330 596908 251398 596964
rect 251454 596908 251522 596964
rect 251578 596908 251646 596964
rect 251702 596908 251798 596964
rect 251178 596840 251798 596908
rect 251178 596784 251274 596840
rect 251330 596784 251398 596840
rect 251454 596784 251522 596840
rect 251578 596784 251646 596840
rect 251702 596784 251798 596840
rect 251178 580350 251798 596784
rect 251178 580294 251274 580350
rect 251330 580294 251398 580350
rect 251454 580294 251522 580350
rect 251578 580294 251646 580350
rect 251702 580294 251798 580350
rect 251178 580226 251798 580294
rect 251178 580170 251274 580226
rect 251330 580170 251398 580226
rect 251454 580170 251522 580226
rect 251578 580170 251646 580226
rect 251702 580170 251798 580226
rect 251178 580102 251798 580170
rect 251178 580046 251274 580102
rect 251330 580046 251398 580102
rect 251454 580046 251522 580102
rect 251578 580046 251646 580102
rect 251702 580046 251798 580102
rect 251178 579978 251798 580046
rect 251178 579922 251274 579978
rect 251330 579922 251398 579978
rect 251454 579922 251522 579978
rect 251578 579922 251646 579978
rect 251702 579922 251798 579978
rect 251178 569342 251798 579922
rect 254898 598172 255518 598268
rect 254898 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 255518 598172
rect 254898 598048 255518 598116
rect 254898 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 255518 598048
rect 254898 597924 255518 597992
rect 254898 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 255518 597924
rect 254898 597800 255518 597868
rect 254898 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 255518 597800
rect 254898 586350 255518 597744
rect 254898 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 255518 586350
rect 254898 586226 255518 586294
rect 254898 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 255518 586226
rect 254898 586102 255518 586170
rect 254898 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 255518 586102
rect 254898 585978 255518 586046
rect 254898 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 255518 585978
rect 254898 569342 255518 585922
rect 281898 597212 282518 598268
rect 281898 597156 281994 597212
rect 282050 597156 282118 597212
rect 282174 597156 282242 597212
rect 282298 597156 282366 597212
rect 282422 597156 282518 597212
rect 281898 597088 282518 597156
rect 281898 597032 281994 597088
rect 282050 597032 282118 597088
rect 282174 597032 282242 597088
rect 282298 597032 282366 597088
rect 282422 597032 282518 597088
rect 281898 596964 282518 597032
rect 281898 596908 281994 596964
rect 282050 596908 282118 596964
rect 282174 596908 282242 596964
rect 282298 596908 282366 596964
rect 282422 596908 282518 596964
rect 281898 596840 282518 596908
rect 281898 596784 281994 596840
rect 282050 596784 282118 596840
rect 282174 596784 282242 596840
rect 282298 596784 282366 596840
rect 282422 596784 282518 596840
rect 281898 580350 282518 596784
rect 281898 580294 281994 580350
rect 282050 580294 282118 580350
rect 282174 580294 282242 580350
rect 282298 580294 282366 580350
rect 282422 580294 282518 580350
rect 281898 580226 282518 580294
rect 281898 580170 281994 580226
rect 282050 580170 282118 580226
rect 282174 580170 282242 580226
rect 282298 580170 282366 580226
rect 282422 580170 282518 580226
rect 281898 580102 282518 580170
rect 281898 580046 281994 580102
rect 282050 580046 282118 580102
rect 282174 580046 282242 580102
rect 282298 580046 282366 580102
rect 282422 580046 282518 580102
rect 281898 579978 282518 580046
rect 281898 579922 281994 579978
rect 282050 579922 282118 579978
rect 282174 579922 282242 579978
rect 282298 579922 282366 579978
rect 282422 579922 282518 579978
rect 281898 569342 282518 579922
rect 285618 598172 286238 598268
rect 285618 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 286238 598172
rect 285618 598048 286238 598116
rect 285618 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 286238 598048
rect 285618 597924 286238 597992
rect 285618 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 286238 597924
rect 285618 597800 286238 597868
rect 285618 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 286238 597800
rect 285618 586350 286238 597744
rect 285618 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 286238 586350
rect 285618 586226 286238 586294
rect 285618 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 286238 586226
rect 285618 586102 286238 586170
rect 285618 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 286238 586102
rect 285618 585978 286238 586046
rect 285618 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 286238 585978
rect 285618 569342 286238 585922
rect 312618 597212 313238 598268
rect 312618 597156 312714 597212
rect 312770 597156 312838 597212
rect 312894 597156 312962 597212
rect 313018 597156 313086 597212
rect 313142 597156 313238 597212
rect 312618 597088 313238 597156
rect 312618 597032 312714 597088
rect 312770 597032 312838 597088
rect 312894 597032 312962 597088
rect 313018 597032 313086 597088
rect 313142 597032 313238 597088
rect 312618 596964 313238 597032
rect 312618 596908 312714 596964
rect 312770 596908 312838 596964
rect 312894 596908 312962 596964
rect 313018 596908 313086 596964
rect 313142 596908 313238 596964
rect 312618 596840 313238 596908
rect 312618 596784 312714 596840
rect 312770 596784 312838 596840
rect 312894 596784 312962 596840
rect 313018 596784 313086 596840
rect 313142 596784 313238 596840
rect 312618 580350 313238 596784
rect 312618 580294 312714 580350
rect 312770 580294 312838 580350
rect 312894 580294 312962 580350
rect 313018 580294 313086 580350
rect 313142 580294 313238 580350
rect 312618 580226 313238 580294
rect 312618 580170 312714 580226
rect 312770 580170 312838 580226
rect 312894 580170 312962 580226
rect 313018 580170 313086 580226
rect 313142 580170 313238 580226
rect 312618 580102 313238 580170
rect 312618 580046 312714 580102
rect 312770 580046 312838 580102
rect 312894 580046 312962 580102
rect 313018 580046 313086 580102
rect 313142 580046 313238 580102
rect 312618 579978 313238 580046
rect 312618 579922 312714 579978
rect 312770 579922 312838 579978
rect 312894 579922 312962 579978
rect 313018 579922 313086 579978
rect 313142 579922 313238 579978
rect 312618 569342 313238 579922
rect 316338 598172 316958 598268
rect 316338 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 316958 598172
rect 316338 598048 316958 598116
rect 316338 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 316958 598048
rect 316338 597924 316958 597992
rect 316338 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 316958 597924
rect 316338 597800 316958 597868
rect 316338 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 316958 597800
rect 316338 586350 316958 597744
rect 316338 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 316958 586350
rect 316338 586226 316958 586294
rect 316338 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 316958 586226
rect 316338 586102 316958 586170
rect 316338 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 316958 586102
rect 316338 585978 316958 586046
rect 316338 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 316958 585978
rect 316338 569342 316958 585922
rect 343338 597212 343958 598268
rect 343338 597156 343434 597212
rect 343490 597156 343558 597212
rect 343614 597156 343682 597212
rect 343738 597156 343806 597212
rect 343862 597156 343958 597212
rect 343338 597088 343958 597156
rect 343338 597032 343434 597088
rect 343490 597032 343558 597088
rect 343614 597032 343682 597088
rect 343738 597032 343806 597088
rect 343862 597032 343958 597088
rect 343338 596964 343958 597032
rect 343338 596908 343434 596964
rect 343490 596908 343558 596964
rect 343614 596908 343682 596964
rect 343738 596908 343806 596964
rect 343862 596908 343958 596964
rect 343338 596840 343958 596908
rect 343338 596784 343434 596840
rect 343490 596784 343558 596840
rect 343614 596784 343682 596840
rect 343738 596784 343806 596840
rect 343862 596784 343958 596840
rect 343338 580350 343958 596784
rect 343338 580294 343434 580350
rect 343490 580294 343558 580350
rect 343614 580294 343682 580350
rect 343738 580294 343806 580350
rect 343862 580294 343958 580350
rect 343338 580226 343958 580294
rect 343338 580170 343434 580226
rect 343490 580170 343558 580226
rect 343614 580170 343682 580226
rect 343738 580170 343806 580226
rect 343862 580170 343958 580226
rect 343338 580102 343958 580170
rect 343338 580046 343434 580102
rect 343490 580046 343558 580102
rect 343614 580046 343682 580102
rect 343738 580046 343806 580102
rect 343862 580046 343958 580102
rect 343338 579978 343958 580046
rect 343338 579922 343434 579978
rect 343490 579922 343558 579978
rect 343614 579922 343682 579978
rect 343738 579922 343806 579978
rect 343862 579922 343958 579978
rect 343338 569342 343958 579922
rect 347058 598172 347678 598268
rect 347058 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 347678 598172
rect 347058 598048 347678 598116
rect 347058 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 347678 598048
rect 347058 597924 347678 597992
rect 347058 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 347678 597924
rect 347058 597800 347678 597868
rect 347058 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 347678 597800
rect 347058 586350 347678 597744
rect 347058 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 347678 586350
rect 347058 586226 347678 586294
rect 347058 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 347678 586226
rect 347058 586102 347678 586170
rect 347058 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 347678 586102
rect 347058 585978 347678 586046
rect 347058 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 347678 585978
rect 347058 569342 347678 585922
rect 374058 597212 374678 598268
rect 374058 597156 374154 597212
rect 374210 597156 374278 597212
rect 374334 597156 374402 597212
rect 374458 597156 374526 597212
rect 374582 597156 374678 597212
rect 374058 597088 374678 597156
rect 374058 597032 374154 597088
rect 374210 597032 374278 597088
rect 374334 597032 374402 597088
rect 374458 597032 374526 597088
rect 374582 597032 374678 597088
rect 374058 596964 374678 597032
rect 374058 596908 374154 596964
rect 374210 596908 374278 596964
rect 374334 596908 374402 596964
rect 374458 596908 374526 596964
rect 374582 596908 374678 596964
rect 374058 596840 374678 596908
rect 374058 596784 374154 596840
rect 374210 596784 374278 596840
rect 374334 596784 374402 596840
rect 374458 596784 374526 596840
rect 374582 596784 374678 596840
rect 374058 580350 374678 596784
rect 374058 580294 374154 580350
rect 374210 580294 374278 580350
rect 374334 580294 374402 580350
rect 374458 580294 374526 580350
rect 374582 580294 374678 580350
rect 374058 580226 374678 580294
rect 374058 580170 374154 580226
rect 374210 580170 374278 580226
rect 374334 580170 374402 580226
rect 374458 580170 374526 580226
rect 374582 580170 374678 580226
rect 374058 580102 374678 580170
rect 374058 580046 374154 580102
rect 374210 580046 374278 580102
rect 374334 580046 374402 580102
rect 374458 580046 374526 580102
rect 374582 580046 374678 580102
rect 374058 579978 374678 580046
rect 374058 579922 374154 579978
rect 374210 579922 374278 579978
rect 374334 579922 374402 579978
rect 374458 579922 374526 579978
rect 374582 579922 374678 579978
rect 374058 569342 374678 579922
rect 377778 598172 378398 598268
rect 377778 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 378398 598172
rect 377778 598048 378398 598116
rect 377778 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 378398 598048
rect 377778 597924 378398 597992
rect 377778 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 378398 597924
rect 377778 597800 378398 597868
rect 377778 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 378398 597800
rect 377778 586350 378398 597744
rect 377778 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 378398 586350
rect 377778 586226 378398 586294
rect 377778 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 378398 586226
rect 377778 586102 378398 586170
rect 377778 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 378398 586102
rect 377778 585978 378398 586046
rect 377778 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 378398 585978
rect 377778 569342 378398 585922
rect 404778 597212 405398 598268
rect 404778 597156 404874 597212
rect 404930 597156 404998 597212
rect 405054 597156 405122 597212
rect 405178 597156 405246 597212
rect 405302 597156 405398 597212
rect 404778 597088 405398 597156
rect 404778 597032 404874 597088
rect 404930 597032 404998 597088
rect 405054 597032 405122 597088
rect 405178 597032 405246 597088
rect 405302 597032 405398 597088
rect 404778 596964 405398 597032
rect 404778 596908 404874 596964
rect 404930 596908 404998 596964
rect 405054 596908 405122 596964
rect 405178 596908 405246 596964
rect 405302 596908 405398 596964
rect 404778 596840 405398 596908
rect 404778 596784 404874 596840
rect 404930 596784 404998 596840
rect 405054 596784 405122 596840
rect 405178 596784 405246 596840
rect 405302 596784 405398 596840
rect 404778 580350 405398 596784
rect 408498 598172 409118 598268
rect 408498 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 409118 598172
rect 408498 598048 409118 598116
rect 408498 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 409118 598048
rect 408498 597924 409118 597992
rect 408498 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 409118 597924
rect 408498 597800 409118 597868
rect 408498 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 409118 597800
rect 408268 591332 408324 591342
rect 408268 589978 408324 591276
rect 408268 589912 408324 589922
rect 404778 580294 404874 580350
rect 404930 580294 404998 580350
rect 405054 580294 405122 580350
rect 405178 580294 405246 580350
rect 405302 580294 405398 580350
rect 404778 580226 405398 580294
rect 404778 580170 404874 580226
rect 404930 580170 404998 580226
rect 405054 580170 405122 580226
rect 405178 580170 405246 580226
rect 405302 580170 405398 580226
rect 404778 580102 405398 580170
rect 404778 580046 404874 580102
rect 404930 580046 404998 580102
rect 405054 580046 405122 580102
rect 405178 580046 405246 580102
rect 405302 580046 405398 580102
rect 404778 579978 405398 580046
rect 404778 579922 404874 579978
rect 404930 579922 404998 579978
rect 405054 579922 405122 579978
rect 405178 579922 405246 579978
rect 405302 579922 405398 579978
rect 404778 569342 405398 579922
rect 408498 586350 409118 597744
rect 408498 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 409118 586350
rect 408498 586226 409118 586294
rect 408498 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 409118 586226
rect 408498 586102 409118 586170
rect 408498 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 409118 586102
rect 408498 585978 409118 586046
rect 408498 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 409118 585978
rect 408498 569342 409118 585922
rect 435498 597212 436118 598268
rect 435498 597156 435594 597212
rect 435650 597156 435718 597212
rect 435774 597156 435842 597212
rect 435898 597156 435966 597212
rect 436022 597156 436118 597212
rect 435498 597088 436118 597156
rect 435498 597032 435594 597088
rect 435650 597032 435718 597088
rect 435774 597032 435842 597088
rect 435898 597032 435966 597088
rect 436022 597032 436118 597088
rect 435498 596964 436118 597032
rect 435498 596908 435594 596964
rect 435650 596908 435718 596964
rect 435774 596908 435842 596964
rect 435898 596908 435966 596964
rect 436022 596908 436118 596964
rect 435498 596840 436118 596908
rect 435498 596784 435594 596840
rect 435650 596784 435718 596840
rect 435774 596784 435842 596840
rect 435898 596784 435966 596840
rect 436022 596784 436118 596840
rect 435498 580350 436118 596784
rect 435498 580294 435594 580350
rect 435650 580294 435718 580350
rect 435774 580294 435842 580350
rect 435898 580294 435966 580350
rect 436022 580294 436118 580350
rect 435498 580226 436118 580294
rect 435498 580170 435594 580226
rect 435650 580170 435718 580226
rect 435774 580170 435842 580226
rect 435898 580170 435966 580226
rect 436022 580170 436118 580226
rect 435498 580102 436118 580170
rect 435498 580046 435594 580102
rect 435650 580046 435718 580102
rect 435774 580046 435842 580102
rect 435898 580046 435966 580102
rect 436022 580046 436118 580102
rect 435498 579978 436118 580046
rect 435498 579922 435594 579978
rect 435650 579922 435718 579978
rect 435774 579922 435842 579978
rect 435898 579922 435966 579978
rect 436022 579922 436118 579978
rect 435498 569342 436118 579922
rect 439218 598172 439838 598268
rect 439218 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 439838 598172
rect 439218 598048 439838 598116
rect 439218 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 439838 598048
rect 439218 597924 439838 597992
rect 439218 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 439838 597924
rect 439218 597800 439838 597868
rect 439218 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 439838 597800
rect 439218 586350 439838 597744
rect 439218 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 439838 586350
rect 439218 586226 439838 586294
rect 439218 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 439838 586226
rect 439218 586102 439838 586170
rect 439218 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 439838 586102
rect 439218 585978 439838 586046
rect 439218 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 439838 585978
rect 439218 569342 439838 585922
rect 466218 597212 466838 598268
rect 466218 597156 466314 597212
rect 466370 597156 466438 597212
rect 466494 597156 466562 597212
rect 466618 597156 466686 597212
rect 466742 597156 466838 597212
rect 466218 597088 466838 597156
rect 466218 597032 466314 597088
rect 466370 597032 466438 597088
rect 466494 597032 466562 597088
rect 466618 597032 466686 597088
rect 466742 597032 466838 597088
rect 466218 596964 466838 597032
rect 466218 596908 466314 596964
rect 466370 596908 466438 596964
rect 466494 596908 466562 596964
rect 466618 596908 466686 596964
rect 466742 596908 466838 596964
rect 466218 596840 466838 596908
rect 466218 596784 466314 596840
rect 466370 596784 466438 596840
rect 466494 596784 466562 596840
rect 466618 596784 466686 596840
rect 466742 596784 466838 596840
rect 466218 580350 466838 596784
rect 466218 580294 466314 580350
rect 466370 580294 466438 580350
rect 466494 580294 466562 580350
rect 466618 580294 466686 580350
rect 466742 580294 466838 580350
rect 466218 580226 466838 580294
rect 466218 580170 466314 580226
rect 466370 580170 466438 580226
rect 466494 580170 466562 580226
rect 466618 580170 466686 580226
rect 466742 580170 466838 580226
rect 466218 580102 466838 580170
rect 466218 580046 466314 580102
rect 466370 580046 466438 580102
rect 466494 580046 466562 580102
rect 466618 580046 466686 580102
rect 466742 580046 466838 580102
rect 466218 579978 466838 580046
rect 466218 579922 466314 579978
rect 466370 579922 466438 579978
rect 466494 579922 466562 579978
rect 466618 579922 466686 579978
rect 466742 579922 466838 579978
rect 466218 569342 466838 579922
rect 469938 598172 470558 598268
rect 469938 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 470558 598172
rect 469938 598048 470558 598116
rect 469938 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 470558 598048
rect 469938 597924 470558 597992
rect 469938 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 470558 597924
rect 469938 597800 470558 597868
rect 469938 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 470558 597800
rect 469938 586350 470558 597744
rect 496938 597212 497558 598268
rect 496938 597156 497034 597212
rect 497090 597156 497158 597212
rect 497214 597156 497282 597212
rect 497338 597156 497406 597212
rect 497462 597156 497558 597212
rect 496938 597088 497558 597156
rect 496938 597032 497034 597088
rect 497090 597032 497158 597088
rect 497214 597032 497282 597088
rect 497338 597032 497406 597088
rect 497462 597032 497558 597088
rect 496938 596964 497558 597032
rect 496938 596908 497034 596964
rect 497090 596908 497158 596964
rect 497214 596908 497282 596964
rect 497338 596908 497406 596964
rect 497462 596908 497558 596964
rect 496938 596840 497558 596908
rect 496938 596784 497034 596840
rect 497090 596784 497158 596840
rect 497214 596784 497282 596840
rect 497338 596784 497406 596840
rect 497462 596784 497558 596840
rect 474348 591332 474404 591342
rect 474348 589798 474404 591276
rect 474348 589732 474404 589742
rect 469938 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 470558 586350
rect 469938 586226 470558 586294
rect 469938 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 470558 586226
rect 469938 586102 470558 586170
rect 469938 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 470558 586102
rect 469938 585978 470558 586046
rect 469938 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 470558 585978
rect 469938 569342 470558 585922
rect 496938 580350 497558 596784
rect 496938 580294 497034 580350
rect 497090 580294 497158 580350
rect 497214 580294 497282 580350
rect 497338 580294 497406 580350
rect 497462 580294 497558 580350
rect 496938 580226 497558 580294
rect 496938 580170 497034 580226
rect 497090 580170 497158 580226
rect 497214 580170 497282 580226
rect 497338 580170 497406 580226
rect 497462 580170 497558 580226
rect 496938 580102 497558 580170
rect 496938 580046 497034 580102
rect 497090 580046 497158 580102
rect 497214 580046 497282 580102
rect 497338 580046 497406 580102
rect 497462 580046 497558 580102
rect 496938 579978 497558 580046
rect 496938 579922 497034 579978
rect 497090 579922 497158 579978
rect 497214 579922 497282 579978
rect 497338 579922 497406 579978
rect 497462 579922 497558 579978
rect 496938 569342 497558 579922
rect 500658 598172 501278 598268
rect 500658 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 501278 598172
rect 500658 598048 501278 598116
rect 500658 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 501278 598048
rect 500658 597924 501278 597992
rect 500658 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 501278 597924
rect 500658 597800 501278 597868
rect 500658 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 501278 597800
rect 500658 586350 501278 597744
rect 500658 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 501278 586350
rect 500658 586226 501278 586294
rect 500658 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 501278 586226
rect 500658 586102 501278 586170
rect 500658 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 501278 586102
rect 500658 585978 501278 586046
rect 500658 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 501278 585978
rect 500658 569342 501278 585922
rect 527658 597212 528278 598268
rect 527658 597156 527754 597212
rect 527810 597156 527878 597212
rect 527934 597156 528002 597212
rect 528058 597156 528126 597212
rect 528182 597156 528278 597212
rect 527658 597088 528278 597156
rect 527658 597032 527754 597088
rect 527810 597032 527878 597088
rect 527934 597032 528002 597088
rect 528058 597032 528126 597088
rect 528182 597032 528278 597088
rect 527658 596964 528278 597032
rect 527658 596908 527754 596964
rect 527810 596908 527878 596964
rect 527934 596908 528002 596964
rect 528058 596908 528126 596964
rect 528182 596908 528278 596964
rect 527658 596840 528278 596908
rect 527658 596784 527754 596840
rect 527810 596784 527878 596840
rect 527934 596784 528002 596840
rect 528058 596784 528126 596840
rect 528182 596784 528278 596840
rect 527658 580350 528278 596784
rect 527658 580294 527754 580350
rect 527810 580294 527878 580350
rect 527934 580294 528002 580350
rect 528058 580294 528126 580350
rect 528182 580294 528278 580350
rect 527658 580226 528278 580294
rect 527658 580170 527754 580226
rect 527810 580170 527878 580226
rect 527934 580170 528002 580226
rect 528058 580170 528126 580226
rect 528182 580170 528278 580226
rect 527658 580102 528278 580170
rect 527658 580046 527754 580102
rect 527810 580046 527878 580102
rect 527934 580046 528002 580102
rect 528058 580046 528126 580102
rect 528182 580046 528278 580102
rect 527658 579978 528278 580046
rect 527658 579922 527754 579978
rect 527810 579922 527878 579978
rect 527934 579922 528002 579978
rect 528058 579922 528126 579978
rect 528182 579922 528278 579978
rect 527658 569342 528278 579922
rect 531378 598172 531998 598268
rect 531378 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 531998 598172
rect 531378 598048 531998 598116
rect 531378 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 531998 598048
rect 531378 597924 531998 597992
rect 531378 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 531998 597924
rect 531378 597800 531998 597868
rect 531378 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 531998 597800
rect 531378 586350 531998 597744
rect 558378 597212 558998 598268
rect 558378 597156 558474 597212
rect 558530 597156 558598 597212
rect 558654 597156 558722 597212
rect 558778 597156 558846 597212
rect 558902 597156 558998 597212
rect 558378 597088 558998 597156
rect 558378 597032 558474 597088
rect 558530 597032 558598 597088
rect 558654 597032 558722 597088
rect 558778 597032 558846 597088
rect 558902 597032 558998 597088
rect 558378 596964 558998 597032
rect 558378 596908 558474 596964
rect 558530 596908 558598 596964
rect 558654 596908 558722 596964
rect 558778 596908 558846 596964
rect 558902 596908 558998 596964
rect 558378 596840 558998 596908
rect 558378 596784 558474 596840
rect 558530 596784 558598 596840
rect 558654 596784 558722 596840
rect 558778 596784 558846 596840
rect 558902 596784 558998 596840
rect 546028 590660 546084 590670
rect 531378 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 531998 586350
rect 531378 586226 531998 586294
rect 531378 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 531998 586226
rect 531378 586102 531998 586170
rect 531378 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 531998 586102
rect 531378 585978 531998 586046
rect 531378 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 531998 585978
rect 531378 569342 531998 585922
rect 545580 590548 545636 590558
rect 194448 562350 194768 562384
rect 194448 562294 194518 562350
rect 194574 562294 194642 562350
rect 194698 562294 194768 562350
rect 194448 562226 194768 562294
rect 194448 562170 194518 562226
rect 194574 562170 194642 562226
rect 194698 562170 194768 562226
rect 194448 562102 194768 562170
rect 194448 562046 194518 562102
rect 194574 562046 194642 562102
rect 194698 562046 194768 562102
rect 194448 561978 194768 562046
rect 194448 561922 194518 561978
rect 194574 561922 194642 561978
rect 194698 561922 194768 561978
rect 194448 561888 194768 561922
rect 225168 562350 225488 562384
rect 225168 562294 225238 562350
rect 225294 562294 225362 562350
rect 225418 562294 225488 562350
rect 225168 562226 225488 562294
rect 225168 562170 225238 562226
rect 225294 562170 225362 562226
rect 225418 562170 225488 562226
rect 225168 562102 225488 562170
rect 225168 562046 225238 562102
rect 225294 562046 225362 562102
rect 225418 562046 225488 562102
rect 225168 561978 225488 562046
rect 225168 561922 225238 561978
rect 225294 561922 225362 561978
rect 225418 561922 225488 561978
rect 225168 561888 225488 561922
rect 255888 562350 256208 562384
rect 255888 562294 255958 562350
rect 256014 562294 256082 562350
rect 256138 562294 256208 562350
rect 255888 562226 256208 562294
rect 255888 562170 255958 562226
rect 256014 562170 256082 562226
rect 256138 562170 256208 562226
rect 255888 562102 256208 562170
rect 255888 562046 255958 562102
rect 256014 562046 256082 562102
rect 256138 562046 256208 562102
rect 255888 561978 256208 562046
rect 255888 561922 255958 561978
rect 256014 561922 256082 561978
rect 256138 561922 256208 561978
rect 255888 561888 256208 561922
rect 286608 562350 286928 562384
rect 286608 562294 286678 562350
rect 286734 562294 286802 562350
rect 286858 562294 286928 562350
rect 286608 562226 286928 562294
rect 286608 562170 286678 562226
rect 286734 562170 286802 562226
rect 286858 562170 286928 562226
rect 286608 562102 286928 562170
rect 286608 562046 286678 562102
rect 286734 562046 286802 562102
rect 286858 562046 286928 562102
rect 286608 561978 286928 562046
rect 286608 561922 286678 561978
rect 286734 561922 286802 561978
rect 286858 561922 286928 561978
rect 286608 561888 286928 561922
rect 317328 562350 317648 562384
rect 317328 562294 317398 562350
rect 317454 562294 317522 562350
rect 317578 562294 317648 562350
rect 317328 562226 317648 562294
rect 317328 562170 317398 562226
rect 317454 562170 317522 562226
rect 317578 562170 317648 562226
rect 317328 562102 317648 562170
rect 317328 562046 317398 562102
rect 317454 562046 317522 562102
rect 317578 562046 317648 562102
rect 317328 561978 317648 562046
rect 317328 561922 317398 561978
rect 317454 561922 317522 561978
rect 317578 561922 317648 561978
rect 317328 561888 317648 561922
rect 348048 562350 348368 562384
rect 348048 562294 348118 562350
rect 348174 562294 348242 562350
rect 348298 562294 348368 562350
rect 348048 562226 348368 562294
rect 348048 562170 348118 562226
rect 348174 562170 348242 562226
rect 348298 562170 348368 562226
rect 348048 562102 348368 562170
rect 348048 562046 348118 562102
rect 348174 562046 348242 562102
rect 348298 562046 348368 562102
rect 348048 561978 348368 562046
rect 348048 561922 348118 561978
rect 348174 561922 348242 561978
rect 348298 561922 348368 561978
rect 348048 561888 348368 561922
rect 378768 562350 379088 562384
rect 378768 562294 378838 562350
rect 378894 562294 378962 562350
rect 379018 562294 379088 562350
rect 378768 562226 379088 562294
rect 378768 562170 378838 562226
rect 378894 562170 378962 562226
rect 379018 562170 379088 562226
rect 378768 562102 379088 562170
rect 378768 562046 378838 562102
rect 378894 562046 378962 562102
rect 379018 562046 379088 562102
rect 378768 561978 379088 562046
rect 378768 561922 378838 561978
rect 378894 561922 378962 561978
rect 379018 561922 379088 561978
rect 378768 561888 379088 561922
rect 409488 562350 409808 562384
rect 409488 562294 409558 562350
rect 409614 562294 409682 562350
rect 409738 562294 409808 562350
rect 409488 562226 409808 562294
rect 409488 562170 409558 562226
rect 409614 562170 409682 562226
rect 409738 562170 409808 562226
rect 409488 562102 409808 562170
rect 409488 562046 409558 562102
rect 409614 562046 409682 562102
rect 409738 562046 409808 562102
rect 409488 561978 409808 562046
rect 409488 561922 409558 561978
rect 409614 561922 409682 561978
rect 409738 561922 409808 561978
rect 409488 561888 409808 561922
rect 440208 562350 440528 562384
rect 440208 562294 440278 562350
rect 440334 562294 440402 562350
rect 440458 562294 440528 562350
rect 440208 562226 440528 562294
rect 440208 562170 440278 562226
rect 440334 562170 440402 562226
rect 440458 562170 440528 562226
rect 440208 562102 440528 562170
rect 440208 562046 440278 562102
rect 440334 562046 440402 562102
rect 440458 562046 440528 562102
rect 440208 561978 440528 562046
rect 440208 561922 440278 561978
rect 440334 561922 440402 561978
rect 440458 561922 440528 561978
rect 440208 561888 440528 561922
rect 470928 562350 471248 562384
rect 470928 562294 470998 562350
rect 471054 562294 471122 562350
rect 471178 562294 471248 562350
rect 470928 562226 471248 562294
rect 470928 562170 470998 562226
rect 471054 562170 471122 562226
rect 471178 562170 471248 562226
rect 470928 562102 471248 562170
rect 470928 562046 470998 562102
rect 471054 562046 471122 562102
rect 471178 562046 471248 562102
rect 470928 561978 471248 562046
rect 470928 561922 470998 561978
rect 471054 561922 471122 561978
rect 471178 561922 471248 561978
rect 470928 561888 471248 561922
rect 501648 562350 501968 562384
rect 501648 562294 501718 562350
rect 501774 562294 501842 562350
rect 501898 562294 501968 562350
rect 501648 562226 501968 562294
rect 501648 562170 501718 562226
rect 501774 562170 501842 562226
rect 501898 562170 501968 562226
rect 501648 562102 501968 562170
rect 501648 562046 501718 562102
rect 501774 562046 501842 562102
rect 501898 562046 501968 562102
rect 501648 561978 501968 562046
rect 501648 561922 501718 561978
rect 501774 561922 501842 561978
rect 501898 561922 501968 561978
rect 501648 561888 501968 561922
rect 532368 562350 532688 562384
rect 532368 562294 532438 562350
rect 532494 562294 532562 562350
rect 532618 562294 532688 562350
rect 532368 562226 532688 562294
rect 532368 562170 532438 562226
rect 532494 562170 532562 562226
rect 532618 562170 532688 562226
rect 532368 562102 532688 562170
rect 532368 562046 532438 562102
rect 532494 562046 532562 562102
rect 532618 562046 532688 562102
rect 532368 561978 532688 562046
rect 532368 561922 532438 561978
rect 532494 561922 532562 561978
rect 532618 561922 532688 561978
rect 532368 561888 532688 561922
rect 209808 550350 210128 550384
rect 209808 550294 209878 550350
rect 209934 550294 210002 550350
rect 210058 550294 210128 550350
rect 209808 550226 210128 550294
rect 209808 550170 209878 550226
rect 209934 550170 210002 550226
rect 210058 550170 210128 550226
rect 209808 550102 210128 550170
rect 209808 550046 209878 550102
rect 209934 550046 210002 550102
rect 210058 550046 210128 550102
rect 209808 549978 210128 550046
rect 209808 549922 209878 549978
rect 209934 549922 210002 549978
rect 210058 549922 210128 549978
rect 209808 549888 210128 549922
rect 240528 550350 240848 550384
rect 240528 550294 240598 550350
rect 240654 550294 240722 550350
rect 240778 550294 240848 550350
rect 240528 550226 240848 550294
rect 240528 550170 240598 550226
rect 240654 550170 240722 550226
rect 240778 550170 240848 550226
rect 240528 550102 240848 550170
rect 240528 550046 240598 550102
rect 240654 550046 240722 550102
rect 240778 550046 240848 550102
rect 240528 549978 240848 550046
rect 240528 549922 240598 549978
rect 240654 549922 240722 549978
rect 240778 549922 240848 549978
rect 240528 549888 240848 549922
rect 271248 550350 271568 550384
rect 271248 550294 271318 550350
rect 271374 550294 271442 550350
rect 271498 550294 271568 550350
rect 271248 550226 271568 550294
rect 271248 550170 271318 550226
rect 271374 550170 271442 550226
rect 271498 550170 271568 550226
rect 271248 550102 271568 550170
rect 271248 550046 271318 550102
rect 271374 550046 271442 550102
rect 271498 550046 271568 550102
rect 271248 549978 271568 550046
rect 271248 549922 271318 549978
rect 271374 549922 271442 549978
rect 271498 549922 271568 549978
rect 271248 549888 271568 549922
rect 301968 550350 302288 550384
rect 301968 550294 302038 550350
rect 302094 550294 302162 550350
rect 302218 550294 302288 550350
rect 301968 550226 302288 550294
rect 301968 550170 302038 550226
rect 302094 550170 302162 550226
rect 302218 550170 302288 550226
rect 301968 550102 302288 550170
rect 301968 550046 302038 550102
rect 302094 550046 302162 550102
rect 302218 550046 302288 550102
rect 301968 549978 302288 550046
rect 301968 549922 302038 549978
rect 302094 549922 302162 549978
rect 302218 549922 302288 549978
rect 301968 549888 302288 549922
rect 332688 550350 333008 550384
rect 332688 550294 332758 550350
rect 332814 550294 332882 550350
rect 332938 550294 333008 550350
rect 332688 550226 333008 550294
rect 332688 550170 332758 550226
rect 332814 550170 332882 550226
rect 332938 550170 333008 550226
rect 332688 550102 333008 550170
rect 332688 550046 332758 550102
rect 332814 550046 332882 550102
rect 332938 550046 333008 550102
rect 332688 549978 333008 550046
rect 332688 549922 332758 549978
rect 332814 549922 332882 549978
rect 332938 549922 333008 549978
rect 332688 549888 333008 549922
rect 363408 550350 363728 550384
rect 363408 550294 363478 550350
rect 363534 550294 363602 550350
rect 363658 550294 363728 550350
rect 363408 550226 363728 550294
rect 363408 550170 363478 550226
rect 363534 550170 363602 550226
rect 363658 550170 363728 550226
rect 363408 550102 363728 550170
rect 363408 550046 363478 550102
rect 363534 550046 363602 550102
rect 363658 550046 363728 550102
rect 363408 549978 363728 550046
rect 363408 549922 363478 549978
rect 363534 549922 363602 549978
rect 363658 549922 363728 549978
rect 363408 549888 363728 549922
rect 394128 550350 394448 550384
rect 394128 550294 394198 550350
rect 394254 550294 394322 550350
rect 394378 550294 394448 550350
rect 394128 550226 394448 550294
rect 394128 550170 394198 550226
rect 394254 550170 394322 550226
rect 394378 550170 394448 550226
rect 394128 550102 394448 550170
rect 394128 550046 394198 550102
rect 394254 550046 394322 550102
rect 394378 550046 394448 550102
rect 394128 549978 394448 550046
rect 394128 549922 394198 549978
rect 394254 549922 394322 549978
rect 394378 549922 394448 549978
rect 394128 549888 394448 549922
rect 424848 550350 425168 550384
rect 424848 550294 424918 550350
rect 424974 550294 425042 550350
rect 425098 550294 425168 550350
rect 424848 550226 425168 550294
rect 424848 550170 424918 550226
rect 424974 550170 425042 550226
rect 425098 550170 425168 550226
rect 424848 550102 425168 550170
rect 424848 550046 424918 550102
rect 424974 550046 425042 550102
rect 425098 550046 425168 550102
rect 424848 549978 425168 550046
rect 424848 549922 424918 549978
rect 424974 549922 425042 549978
rect 425098 549922 425168 549978
rect 424848 549888 425168 549922
rect 455568 550350 455888 550384
rect 455568 550294 455638 550350
rect 455694 550294 455762 550350
rect 455818 550294 455888 550350
rect 455568 550226 455888 550294
rect 455568 550170 455638 550226
rect 455694 550170 455762 550226
rect 455818 550170 455888 550226
rect 455568 550102 455888 550170
rect 455568 550046 455638 550102
rect 455694 550046 455762 550102
rect 455818 550046 455888 550102
rect 455568 549978 455888 550046
rect 455568 549922 455638 549978
rect 455694 549922 455762 549978
rect 455818 549922 455888 549978
rect 455568 549888 455888 549922
rect 486288 550350 486608 550384
rect 486288 550294 486358 550350
rect 486414 550294 486482 550350
rect 486538 550294 486608 550350
rect 486288 550226 486608 550294
rect 486288 550170 486358 550226
rect 486414 550170 486482 550226
rect 486538 550170 486608 550226
rect 486288 550102 486608 550170
rect 486288 550046 486358 550102
rect 486414 550046 486482 550102
rect 486538 550046 486608 550102
rect 486288 549978 486608 550046
rect 486288 549922 486358 549978
rect 486414 549922 486482 549978
rect 486538 549922 486608 549978
rect 486288 549888 486608 549922
rect 517008 550350 517328 550384
rect 517008 550294 517078 550350
rect 517134 550294 517202 550350
rect 517258 550294 517328 550350
rect 517008 550226 517328 550294
rect 517008 550170 517078 550226
rect 517134 550170 517202 550226
rect 517258 550170 517328 550226
rect 517008 550102 517328 550170
rect 517008 550046 517078 550102
rect 517134 550046 517202 550102
rect 517258 550046 517328 550102
rect 517008 549978 517328 550046
rect 517008 549922 517078 549978
rect 517134 549922 517202 549978
rect 517258 549922 517328 549978
rect 517008 549888 517328 549922
rect 194448 544350 194768 544384
rect 194448 544294 194518 544350
rect 194574 544294 194642 544350
rect 194698 544294 194768 544350
rect 194448 544226 194768 544294
rect 194448 544170 194518 544226
rect 194574 544170 194642 544226
rect 194698 544170 194768 544226
rect 194448 544102 194768 544170
rect 194448 544046 194518 544102
rect 194574 544046 194642 544102
rect 194698 544046 194768 544102
rect 194448 543978 194768 544046
rect 194448 543922 194518 543978
rect 194574 543922 194642 543978
rect 194698 543922 194768 543978
rect 194448 543888 194768 543922
rect 225168 544350 225488 544384
rect 225168 544294 225238 544350
rect 225294 544294 225362 544350
rect 225418 544294 225488 544350
rect 225168 544226 225488 544294
rect 225168 544170 225238 544226
rect 225294 544170 225362 544226
rect 225418 544170 225488 544226
rect 225168 544102 225488 544170
rect 225168 544046 225238 544102
rect 225294 544046 225362 544102
rect 225418 544046 225488 544102
rect 225168 543978 225488 544046
rect 225168 543922 225238 543978
rect 225294 543922 225362 543978
rect 225418 543922 225488 543978
rect 225168 543888 225488 543922
rect 255888 544350 256208 544384
rect 255888 544294 255958 544350
rect 256014 544294 256082 544350
rect 256138 544294 256208 544350
rect 255888 544226 256208 544294
rect 255888 544170 255958 544226
rect 256014 544170 256082 544226
rect 256138 544170 256208 544226
rect 255888 544102 256208 544170
rect 255888 544046 255958 544102
rect 256014 544046 256082 544102
rect 256138 544046 256208 544102
rect 255888 543978 256208 544046
rect 255888 543922 255958 543978
rect 256014 543922 256082 543978
rect 256138 543922 256208 543978
rect 255888 543888 256208 543922
rect 286608 544350 286928 544384
rect 286608 544294 286678 544350
rect 286734 544294 286802 544350
rect 286858 544294 286928 544350
rect 286608 544226 286928 544294
rect 286608 544170 286678 544226
rect 286734 544170 286802 544226
rect 286858 544170 286928 544226
rect 286608 544102 286928 544170
rect 286608 544046 286678 544102
rect 286734 544046 286802 544102
rect 286858 544046 286928 544102
rect 286608 543978 286928 544046
rect 286608 543922 286678 543978
rect 286734 543922 286802 543978
rect 286858 543922 286928 543978
rect 286608 543888 286928 543922
rect 317328 544350 317648 544384
rect 317328 544294 317398 544350
rect 317454 544294 317522 544350
rect 317578 544294 317648 544350
rect 317328 544226 317648 544294
rect 317328 544170 317398 544226
rect 317454 544170 317522 544226
rect 317578 544170 317648 544226
rect 317328 544102 317648 544170
rect 317328 544046 317398 544102
rect 317454 544046 317522 544102
rect 317578 544046 317648 544102
rect 317328 543978 317648 544046
rect 317328 543922 317398 543978
rect 317454 543922 317522 543978
rect 317578 543922 317648 543978
rect 317328 543888 317648 543922
rect 348048 544350 348368 544384
rect 348048 544294 348118 544350
rect 348174 544294 348242 544350
rect 348298 544294 348368 544350
rect 348048 544226 348368 544294
rect 348048 544170 348118 544226
rect 348174 544170 348242 544226
rect 348298 544170 348368 544226
rect 348048 544102 348368 544170
rect 348048 544046 348118 544102
rect 348174 544046 348242 544102
rect 348298 544046 348368 544102
rect 348048 543978 348368 544046
rect 348048 543922 348118 543978
rect 348174 543922 348242 543978
rect 348298 543922 348368 543978
rect 348048 543888 348368 543922
rect 378768 544350 379088 544384
rect 378768 544294 378838 544350
rect 378894 544294 378962 544350
rect 379018 544294 379088 544350
rect 378768 544226 379088 544294
rect 378768 544170 378838 544226
rect 378894 544170 378962 544226
rect 379018 544170 379088 544226
rect 378768 544102 379088 544170
rect 378768 544046 378838 544102
rect 378894 544046 378962 544102
rect 379018 544046 379088 544102
rect 378768 543978 379088 544046
rect 378768 543922 378838 543978
rect 378894 543922 378962 543978
rect 379018 543922 379088 543978
rect 378768 543888 379088 543922
rect 409488 544350 409808 544384
rect 409488 544294 409558 544350
rect 409614 544294 409682 544350
rect 409738 544294 409808 544350
rect 409488 544226 409808 544294
rect 409488 544170 409558 544226
rect 409614 544170 409682 544226
rect 409738 544170 409808 544226
rect 409488 544102 409808 544170
rect 409488 544046 409558 544102
rect 409614 544046 409682 544102
rect 409738 544046 409808 544102
rect 409488 543978 409808 544046
rect 409488 543922 409558 543978
rect 409614 543922 409682 543978
rect 409738 543922 409808 543978
rect 409488 543888 409808 543922
rect 440208 544350 440528 544384
rect 440208 544294 440278 544350
rect 440334 544294 440402 544350
rect 440458 544294 440528 544350
rect 440208 544226 440528 544294
rect 440208 544170 440278 544226
rect 440334 544170 440402 544226
rect 440458 544170 440528 544226
rect 440208 544102 440528 544170
rect 440208 544046 440278 544102
rect 440334 544046 440402 544102
rect 440458 544046 440528 544102
rect 440208 543978 440528 544046
rect 440208 543922 440278 543978
rect 440334 543922 440402 543978
rect 440458 543922 440528 543978
rect 440208 543888 440528 543922
rect 470928 544350 471248 544384
rect 470928 544294 470998 544350
rect 471054 544294 471122 544350
rect 471178 544294 471248 544350
rect 470928 544226 471248 544294
rect 470928 544170 470998 544226
rect 471054 544170 471122 544226
rect 471178 544170 471248 544226
rect 470928 544102 471248 544170
rect 470928 544046 470998 544102
rect 471054 544046 471122 544102
rect 471178 544046 471248 544102
rect 470928 543978 471248 544046
rect 470928 543922 470998 543978
rect 471054 543922 471122 543978
rect 471178 543922 471248 543978
rect 470928 543888 471248 543922
rect 501648 544350 501968 544384
rect 501648 544294 501718 544350
rect 501774 544294 501842 544350
rect 501898 544294 501968 544350
rect 501648 544226 501968 544294
rect 501648 544170 501718 544226
rect 501774 544170 501842 544226
rect 501898 544170 501968 544226
rect 501648 544102 501968 544170
rect 501648 544046 501718 544102
rect 501774 544046 501842 544102
rect 501898 544046 501968 544102
rect 501648 543978 501968 544046
rect 501648 543922 501718 543978
rect 501774 543922 501842 543978
rect 501898 543922 501968 543978
rect 501648 543888 501968 543922
rect 532368 544350 532688 544384
rect 532368 544294 532438 544350
rect 532494 544294 532562 544350
rect 532618 544294 532688 544350
rect 532368 544226 532688 544294
rect 532368 544170 532438 544226
rect 532494 544170 532562 544226
rect 532618 544170 532688 544226
rect 532368 544102 532688 544170
rect 532368 544046 532438 544102
rect 532494 544046 532562 544102
rect 532618 544046 532688 544102
rect 532368 543978 532688 544046
rect 532368 543922 532438 543978
rect 532494 543922 532562 543978
rect 532618 543922 532688 543978
rect 532368 543888 532688 543922
rect 209808 532350 210128 532384
rect 209808 532294 209878 532350
rect 209934 532294 210002 532350
rect 210058 532294 210128 532350
rect 209808 532226 210128 532294
rect 209808 532170 209878 532226
rect 209934 532170 210002 532226
rect 210058 532170 210128 532226
rect 209808 532102 210128 532170
rect 209808 532046 209878 532102
rect 209934 532046 210002 532102
rect 210058 532046 210128 532102
rect 209808 531978 210128 532046
rect 209808 531922 209878 531978
rect 209934 531922 210002 531978
rect 210058 531922 210128 531978
rect 209808 531888 210128 531922
rect 240528 532350 240848 532384
rect 240528 532294 240598 532350
rect 240654 532294 240722 532350
rect 240778 532294 240848 532350
rect 240528 532226 240848 532294
rect 240528 532170 240598 532226
rect 240654 532170 240722 532226
rect 240778 532170 240848 532226
rect 240528 532102 240848 532170
rect 240528 532046 240598 532102
rect 240654 532046 240722 532102
rect 240778 532046 240848 532102
rect 240528 531978 240848 532046
rect 240528 531922 240598 531978
rect 240654 531922 240722 531978
rect 240778 531922 240848 531978
rect 240528 531888 240848 531922
rect 271248 532350 271568 532384
rect 271248 532294 271318 532350
rect 271374 532294 271442 532350
rect 271498 532294 271568 532350
rect 271248 532226 271568 532294
rect 271248 532170 271318 532226
rect 271374 532170 271442 532226
rect 271498 532170 271568 532226
rect 271248 532102 271568 532170
rect 271248 532046 271318 532102
rect 271374 532046 271442 532102
rect 271498 532046 271568 532102
rect 271248 531978 271568 532046
rect 271248 531922 271318 531978
rect 271374 531922 271442 531978
rect 271498 531922 271568 531978
rect 271248 531888 271568 531922
rect 301968 532350 302288 532384
rect 301968 532294 302038 532350
rect 302094 532294 302162 532350
rect 302218 532294 302288 532350
rect 301968 532226 302288 532294
rect 301968 532170 302038 532226
rect 302094 532170 302162 532226
rect 302218 532170 302288 532226
rect 301968 532102 302288 532170
rect 301968 532046 302038 532102
rect 302094 532046 302162 532102
rect 302218 532046 302288 532102
rect 301968 531978 302288 532046
rect 301968 531922 302038 531978
rect 302094 531922 302162 531978
rect 302218 531922 302288 531978
rect 301968 531888 302288 531922
rect 332688 532350 333008 532384
rect 332688 532294 332758 532350
rect 332814 532294 332882 532350
rect 332938 532294 333008 532350
rect 332688 532226 333008 532294
rect 332688 532170 332758 532226
rect 332814 532170 332882 532226
rect 332938 532170 333008 532226
rect 332688 532102 333008 532170
rect 332688 532046 332758 532102
rect 332814 532046 332882 532102
rect 332938 532046 333008 532102
rect 332688 531978 333008 532046
rect 332688 531922 332758 531978
rect 332814 531922 332882 531978
rect 332938 531922 333008 531978
rect 332688 531888 333008 531922
rect 363408 532350 363728 532384
rect 363408 532294 363478 532350
rect 363534 532294 363602 532350
rect 363658 532294 363728 532350
rect 363408 532226 363728 532294
rect 363408 532170 363478 532226
rect 363534 532170 363602 532226
rect 363658 532170 363728 532226
rect 363408 532102 363728 532170
rect 363408 532046 363478 532102
rect 363534 532046 363602 532102
rect 363658 532046 363728 532102
rect 363408 531978 363728 532046
rect 363408 531922 363478 531978
rect 363534 531922 363602 531978
rect 363658 531922 363728 531978
rect 363408 531888 363728 531922
rect 394128 532350 394448 532384
rect 394128 532294 394198 532350
rect 394254 532294 394322 532350
rect 394378 532294 394448 532350
rect 394128 532226 394448 532294
rect 394128 532170 394198 532226
rect 394254 532170 394322 532226
rect 394378 532170 394448 532226
rect 394128 532102 394448 532170
rect 394128 532046 394198 532102
rect 394254 532046 394322 532102
rect 394378 532046 394448 532102
rect 394128 531978 394448 532046
rect 394128 531922 394198 531978
rect 394254 531922 394322 531978
rect 394378 531922 394448 531978
rect 394128 531888 394448 531922
rect 424848 532350 425168 532384
rect 424848 532294 424918 532350
rect 424974 532294 425042 532350
rect 425098 532294 425168 532350
rect 424848 532226 425168 532294
rect 424848 532170 424918 532226
rect 424974 532170 425042 532226
rect 425098 532170 425168 532226
rect 424848 532102 425168 532170
rect 424848 532046 424918 532102
rect 424974 532046 425042 532102
rect 425098 532046 425168 532102
rect 424848 531978 425168 532046
rect 424848 531922 424918 531978
rect 424974 531922 425042 531978
rect 425098 531922 425168 531978
rect 424848 531888 425168 531922
rect 455568 532350 455888 532384
rect 455568 532294 455638 532350
rect 455694 532294 455762 532350
rect 455818 532294 455888 532350
rect 455568 532226 455888 532294
rect 455568 532170 455638 532226
rect 455694 532170 455762 532226
rect 455818 532170 455888 532226
rect 455568 532102 455888 532170
rect 455568 532046 455638 532102
rect 455694 532046 455762 532102
rect 455818 532046 455888 532102
rect 455568 531978 455888 532046
rect 455568 531922 455638 531978
rect 455694 531922 455762 531978
rect 455818 531922 455888 531978
rect 455568 531888 455888 531922
rect 486288 532350 486608 532384
rect 486288 532294 486358 532350
rect 486414 532294 486482 532350
rect 486538 532294 486608 532350
rect 486288 532226 486608 532294
rect 486288 532170 486358 532226
rect 486414 532170 486482 532226
rect 486538 532170 486608 532226
rect 486288 532102 486608 532170
rect 486288 532046 486358 532102
rect 486414 532046 486482 532102
rect 486538 532046 486608 532102
rect 486288 531978 486608 532046
rect 486288 531922 486358 531978
rect 486414 531922 486482 531978
rect 486538 531922 486608 531978
rect 486288 531888 486608 531922
rect 517008 532350 517328 532384
rect 517008 532294 517078 532350
rect 517134 532294 517202 532350
rect 517258 532294 517328 532350
rect 517008 532226 517328 532294
rect 517008 532170 517078 532226
rect 517134 532170 517202 532226
rect 517258 532170 517328 532226
rect 517008 532102 517328 532170
rect 517008 532046 517078 532102
rect 517134 532046 517202 532102
rect 517258 532046 517328 532102
rect 517008 531978 517328 532046
rect 517008 531922 517078 531978
rect 517134 531922 517202 531978
rect 517258 531922 517328 531978
rect 517008 531888 517328 531922
rect 194448 526350 194768 526384
rect 194448 526294 194518 526350
rect 194574 526294 194642 526350
rect 194698 526294 194768 526350
rect 194448 526226 194768 526294
rect 194448 526170 194518 526226
rect 194574 526170 194642 526226
rect 194698 526170 194768 526226
rect 194448 526102 194768 526170
rect 194448 526046 194518 526102
rect 194574 526046 194642 526102
rect 194698 526046 194768 526102
rect 194448 525978 194768 526046
rect 194448 525922 194518 525978
rect 194574 525922 194642 525978
rect 194698 525922 194768 525978
rect 194448 525888 194768 525922
rect 225168 526350 225488 526384
rect 225168 526294 225238 526350
rect 225294 526294 225362 526350
rect 225418 526294 225488 526350
rect 225168 526226 225488 526294
rect 225168 526170 225238 526226
rect 225294 526170 225362 526226
rect 225418 526170 225488 526226
rect 225168 526102 225488 526170
rect 225168 526046 225238 526102
rect 225294 526046 225362 526102
rect 225418 526046 225488 526102
rect 225168 525978 225488 526046
rect 225168 525922 225238 525978
rect 225294 525922 225362 525978
rect 225418 525922 225488 525978
rect 225168 525888 225488 525922
rect 255888 526350 256208 526384
rect 255888 526294 255958 526350
rect 256014 526294 256082 526350
rect 256138 526294 256208 526350
rect 255888 526226 256208 526294
rect 255888 526170 255958 526226
rect 256014 526170 256082 526226
rect 256138 526170 256208 526226
rect 255888 526102 256208 526170
rect 255888 526046 255958 526102
rect 256014 526046 256082 526102
rect 256138 526046 256208 526102
rect 255888 525978 256208 526046
rect 255888 525922 255958 525978
rect 256014 525922 256082 525978
rect 256138 525922 256208 525978
rect 255888 525888 256208 525922
rect 286608 526350 286928 526384
rect 286608 526294 286678 526350
rect 286734 526294 286802 526350
rect 286858 526294 286928 526350
rect 286608 526226 286928 526294
rect 286608 526170 286678 526226
rect 286734 526170 286802 526226
rect 286858 526170 286928 526226
rect 286608 526102 286928 526170
rect 286608 526046 286678 526102
rect 286734 526046 286802 526102
rect 286858 526046 286928 526102
rect 286608 525978 286928 526046
rect 286608 525922 286678 525978
rect 286734 525922 286802 525978
rect 286858 525922 286928 525978
rect 286608 525888 286928 525922
rect 317328 526350 317648 526384
rect 317328 526294 317398 526350
rect 317454 526294 317522 526350
rect 317578 526294 317648 526350
rect 317328 526226 317648 526294
rect 317328 526170 317398 526226
rect 317454 526170 317522 526226
rect 317578 526170 317648 526226
rect 317328 526102 317648 526170
rect 317328 526046 317398 526102
rect 317454 526046 317522 526102
rect 317578 526046 317648 526102
rect 317328 525978 317648 526046
rect 317328 525922 317398 525978
rect 317454 525922 317522 525978
rect 317578 525922 317648 525978
rect 317328 525888 317648 525922
rect 348048 526350 348368 526384
rect 348048 526294 348118 526350
rect 348174 526294 348242 526350
rect 348298 526294 348368 526350
rect 348048 526226 348368 526294
rect 348048 526170 348118 526226
rect 348174 526170 348242 526226
rect 348298 526170 348368 526226
rect 348048 526102 348368 526170
rect 348048 526046 348118 526102
rect 348174 526046 348242 526102
rect 348298 526046 348368 526102
rect 348048 525978 348368 526046
rect 348048 525922 348118 525978
rect 348174 525922 348242 525978
rect 348298 525922 348368 525978
rect 348048 525888 348368 525922
rect 378768 526350 379088 526384
rect 378768 526294 378838 526350
rect 378894 526294 378962 526350
rect 379018 526294 379088 526350
rect 378768 526226 379088 526294
rect 378768 526170 378838 526226
rect 378894 526170 378962 526226
rect 379018 526170 379088 526226
rect 378768 526102 379088 526170
rect 378768 526046 378838 526102
rect 378894 526046 378962 526102
rect 379018 526046 379088 526102
rect 378768 525978 379088 526046
rect 378768 525922 378838 525978
rect 378894 525922 378962 525978
rect 379018 525922 379088 525978
rect 378768 525888 379088 525922
rect 409488 526350 409808 526384
rect 409488 526294 409558 526350
rect 409614 526294 409682 526350
rect 409738 526294 409808 526350
rect 409488 526226 409808 526294
rect 409488 526170 409558 526226
rect 409614 526170 409682 526226
rect 409738 526170 409808 526226
rect 409488 526102 409808 526170
rect 409488 526046 409558 526102
rect 409614 526046 409682 526102
rect 409738 526046 409808 526102
rect 409488 525978 409808 526046
rect 409488 525922 409558 525978
rect 409614 525922 409682 525978
rect 409738 525922 409808 525978
rect 409488 525888 409808 525922
rect 440208 526350 440528 526384
rect 440208 526294 440278 526350
rect 440334 526294 440402 526350
rect 440458 526294 440528 526350
rect 440208 526226 440528 526294
rect 440208 526170 440278 526226
rect 440334 526170 440402 526226
rect 440458 526170 440528 526226
rect 440208 526102 440528 526170
rect 440208 526046 440278 526102
rect 440334 526046 440402 526102
rect 440458 526046 440528 526102
rect 440208 525978 440528 526046
rect 440208 525922 440278 525978
rect 440334 525922 440402 525978
rect 440458 525922 440528 525978
rect 440208 525888 440528 525922
rect 470928 526350 471248 526384
rect 470928 526294 470998 526350
rect 471054 526294 471122 526350
rect 471178 526294 471248 526350
rect 470928 526226 471248 526294
rect 470928 526170 470998 526226
rect 471054 526170 471122 526226
rect 471178 526170 471248 526226
rect 470928 526102 471248 526170
rect 470928 526046 470998 526102
rect 471054 526046 471122 526102
rect 471178 526046 471248 526102
rect 470928 525978 471248 526046
rect 470928 525922 470998 525978
rect 471054 525922 471122 525978
rect 471178 525922 471248 525978
rect 470928 525888 471248 525922
rect 501648 526350 501968 526384
rect 501648 526294 501718 526350
rect 501774 526294 501842 526350
rect 501898 526294 501968 526350
rect 501648 526226 501968 526294
rect 501648 526170 501718 526226
rect 501774 526170 501842 526226
rect 501898 526170 501968 526226
rect 501648 526102 501968 526170
rect 501648 526046 501718 526102
rect 501774 526046 501842 526102
rect 501898 526046 501968 526102
rect 501648 525978 501968 526046
rect 501648 525922 501718 525978
rect 501774 525922 501842 525978
rect 501898 525922 501968 525978
rect 501648 525888 501968 525922
rect 532368 526350 532688 526384
rect 532368 526294 532438 526350
rect 532494 526294 532562 526350
rect 532618 526294 532688 526350
rect 532368 526226 532688 526294
rect 532368 526170 532438 526226
rect 532494 526170 532562 526226
rect 532618 526170 532688 526226
rect 532368 526102 532688 526170
rect 532368 526046 532438 526102
rect 532494 526046 532562 526102
rect 532618 526046 532688 526102
rect 532368 525978 532688 526046
rect 532368 525922 532438 525978
rect 532494 525922 532562 525978
rect 532618 525922 532688 525978
rect 532368 525888 532688 525922
rect 209808 514350 210128 514384
rect 209808 514294 209878 514350
rect 209934 514294 210002 514350
rect 210058 514294 210128 514350
rect 209808 514226 210128 514294
rect 209808 514170 209878 514226
rect 209934 514170 210002 514226
rect 210058 514170 210128 514226
rect 209808 514102 210128 514170
rect 209808 514046 209878 514102
rect 209934 514046 210002 514102
rect 210058 514046 210128 514102
rect 209808 513978 210128 514046
rect 209808 513922 209878 513978
rect 209934 513922 210002 513978
rect 210058 513922 210128 513978
rect 209808 513888 210128 513922
rect 240528 514350 240848 514384
rect 240528 514294 240598 514350
rect 240654 514294 240722 514350
rect 240778 514294 240848 514350
rect 240528 514226 240848 514294
rect 240528 514170 240598 514226
rect 240654 514170 240722 514226
rect 240778 514170 240848 514226
rect 240528 514102 240848 514170
rect 240528 514046 240598 514102
rect 240654 514046 240722 514102
rect 240778 514046 240848 514102
rect 240528 513978 240848 514046
rect 240528 513922 240598 513978
rect 240654 513922 240722 513978
rect 240778 513922 240848 513978
rect 240528 513888 240848 513922
rect 271248 514350 271568 514384
rect 271248 514294 271318 514350
rect 271374 514294 271442 514350
rect 271498 514294 271568 514350
rect 271248 514226 271568 514294
rect 271248 514170 271318 514226
rect 271374 514170 271442 514226
rect 271498 514170 271568 514226
rect 271248 514102 271568 514170
rect 271248 514046 271318 514102
rect 271374 514046 271442 514102
rect 271498 514046 271568 514102
rect 271248 513978 271568 514046
rect 271248 513922 271318 513978
rect 271374 513922 271442 513978
rect 271498 513922 271568 513978
rect 271248 513888 271568 513922
rect 301968 514350 302288 514384
rect 301968 514294 302038 514350
rect 302094 514294 302162 514350
rect 302218 514294 302288 514350
rect 301968 514226 302288 514294
rect 301968 514170 302038 514226
rect 302094 514170 302162 514226
rect 302218 514170 302288 514226
rect 301968 514102 302288 514170
rect 301968 514046 302038 514102
rect 302094 514046 302162 514102
rect 302218 514046 302288 514102
rect 301968 513978 302288 514046
rect 301968 513922 302038 513978
rect 302094 513922 302162 513978
rect 302218 513922 302288 513978
rect 301968 513888 302288 513922
rect 332688 514350 333008 514384
rect 332688 514294 332758 514350
rect 332814 514294 332882 514350
rect 332938 514294 333008 514350
rect 332688 514226 333008 514294
rect 332688 514170 332758 514226
rect 332814 514170 332882 514226
rect 332938 514170 333008 514226
rect 332688 514102 333008 514170
rect 332688 514046 332758 514102
rect 332814 514046 332882 514102
rect 332938 514046 333008 514102
rect 332688 513978 333008 514046
rect 332688 513922 332758 513978
rect 332814 513922 332882 513978
rect 332938 513922 333008 513978
rect 332688 513888 333008 513922
rect 363408 514350 363728 514384
rect 363408 514294 363478 514350
rect 363534 514294 363602 514350
rect 363658 514294 363728 514350
rect 363408 514226 363728 514294
rect 363408 514170 363478 514226
rect 363534 514170 363602 514226
rect 363658 514170 363728 514226
rect 363408 514102 363728 514170
rect 363408 514046 363478 514102
rect 363534 514046 363602 514102
rect 363658 514046 363728 514102
rect 363408 513978 363728 514046
rect 363408 513922 363478 513978
rect 363534 513922 363602 513978
rect 363658 513922 363728 513978
rect 363408 513888 363728 513922
rect 394128 514350 394448 514384
rect 394128 514294 394198 514350
rect 394254 514294 394322 514350
rect 394378 514294 394448 514350
rect 394128 514226 394448 514294
rect 394128 514170 394198 514226
rect 394254 514170 394322 514226
rect 394378 514170 394448 514226
rect 394128 514102 394448 514170
rect 394128 514046 394198 514102
rect 394254 514046 394322 514102
rect 394378 514046 394448 514102
rect 394128 513978 394448 514046
rect 394128 513922 394198 513978
rect 394254 513922 394322 513978
rect 394378 513922 394448 513978
rect 394128 513888 394448 513922
rect 424848 514350 425168 514384
rect 424848 514294 424918 514350
rect 424974 514294 425042 514350
rect 425098 514294 425168 514350
rect 424848 514226 425168 514294
rect 424848 514170 424918 514226
rect 424974 514170 425042 514226
rect 425098 514170 425168 514226
rect 424848 514102 425168 514170
rect 424848 514046 424918 514102
rect 424974 514046 425042 514102
rect 425098 514046 425168 514102
rect 424848 513978 425168 514046
rect 424848 513922 424918 513978
rect 424974 513922 425042 513978
rect 425098 513922 425168 513978
rect 424848 513888 425168 513922
rect 455568 514350 455888 514384
rect 455568 514294 455638 514350
rect 455694 514294 455762 514350
rect 455818 514294 455888 514350
rect 455568 514226 455888 514294
rect 455568 514170 455638 514226
rect 455694 514170 455762 514226
rect 455818 514170 455888 514226
rect 455568 514102 455888 514170
rect 455568 514046 455638 514102
rect 455694 514046 455762 514102
rect 455818 514046 455888 514102
rect 455568 513978 455888 514046
rect 455568 513922 455638 513978
rect 455694 513922 455762 513978
rect 455818 513922 455888 513978
rect 455568 513888 455888 513922
rect 486288 514350 486608 514384
rect 486288 514294 486358 514350
rect 486414 514294 486482 514350
rect 486538 514294 486608 514350
rect 486288 514226 486608 514294
rect 486288 514170 486358 514226
rect 486414 514170 486482 514226
rect 486538 514170 486608 514226
rect 486288 514102 486608 514170
rect 486288 514046 486358 514102
rect 486414 514046 486482 514102
rect 486538 514046 486608 514102
rect 486288 513978 486608 514046
rect 486288 513922 486358 513978
rect 486414 513922 486482 513978
rect 486538 513922 486608 513978
rect 486288 513888 486608 513922
rect 517008 514350 517328 514384
rect 517008 514294 517078 514350
rect 517134 514294 517202 514350
rect 517258 514294 517328 514350
rect 517008 514226 517328 514294
rect 517008 514170 517078 514226
rect 517134 514170 517202 514226
rect 517258 514170 517328 514226
rect 517008 514102 517328 514170
rect 517008 514046 517078 514102
rect 517134 514046 517202 514102
rect 517258 514046 517328 514102
rect 517008 513978 517328 514046
rect 517008 513922 517078 513978
rect 517134 513922 517202 513978
rect 517258 513922 517328 513978
rect 517008 513888 517328 513922
rect 194448 508350 194768 508384
rect 194448 508294 194518 508350
rect 194574 508294 194642 508350
rect 194698 508294 194768 508350
rect 194448 508226 194768 508294
rect 194448 508170 194518 508226
rect 194574 508170 194642 508226
rect 194698 508170 194768 508226
rect 194448 508102 194768 508170
rect 194448 508046 194518 508102
rect 194574 508046 194642 508102
rect 194698 508046 194768 508102
rect 194448 507978 194768 508046
rect 194448 507922 194518 507978
rect 194574 507922 194642 507978
rect 194698 507922 194768 507978
rect 194448 507888 194768 507922
rect 225168 508350 225488 508384
rect 225168 508294 225238 508350
rect 225294 508294 225362 508350
rect 225418 508294 225488 508350
rect 225168 508226 225488 508294
rect 225168 508170 225238 508226
rect 225294 508170 225362 508226
rect 225418 508170 225488 508226
rect 225168 508102 225488 508170
rect 225168 508046 225238 508102
rect 225294 508046 225362 508102
rect 225418 508046 225488 508102
rect 225168 507978 225488 508046
rect 225168 507922 225238 507978
rect 225294 507922 225362 507978
rect 225418 507922 225488 507978
rect 225168 507888 225488 507922
rect 255888 508350 256208 508384
rect 255888 508294 255958 508350
rect 256014 508294 256082 508350
rect 256138 508294 256208 508350
rect 255888 508226 256208 508294
rect 255888 508170 255958 508226
rect 256014 508170 256082 508226
rect 256138 508170 256208 508226
rect 255888 508102 256208 508170
rect 255888 508046 255958 508102
rect 256014 508046 256082 508102
rect 256138 508046 256208 508102
rect 255888 507978 256208 508046
rect 255888 507922 255958 507978
rect 256014 507922 256082 507978
rect 256138 507922 256208 507978
rect 255888 507888 256208 507922
rect 286608 508350 286928 508384
rect 286608 508294 286678 508350
rect 286734 508294 286802 508350
rect 286858 508294 286928 508350
rect 286608 508226 286928 508294
rect 286608 508170 286678 508226
rect 286734 508170 286802 508226
rect 286858 508170 286928 508226
rect 286608 508102 286928 508170
rect 286608 508046 286678 508102
rect 286734 508046 286802 508102
rect 286858 508046 286928 508102
rect 286608 507978 286928 508046
rect 286608 507922 286678 507978
rect 286734 507922 286802 507978
rect 286858 507922 286928 507978
rect 286608 507888 286928 507922
rect 317328 508350 317648 508384
rect 317328 508294 317398 508350
rect 317454 508294 317522 508350
rect 317578 508294 317648 508350
rect 317328 508226 317648 508294
rect 317328 508170 317398 508226
rect 317454 508170 317522 508226
rect 317578 508170 317648 508226
rect 317328 508102 317648 508170
rect 317328 508046 317398 508102
rect 317454 508046 317522 508102
rect 317578 508046 317648 508102
rect 317328 507978 317648 508046
rect 317328 507922 317398 507978
rect 317454 507922 317522 507978
rect 317578 507922 317648 507978
rect 317328 507888 317648 507922
rect 348048 508350 348368 508384
rect 348048 508294 348118 508350
rect 348174 508294 348242 508350
rect 348298 508294 348368 508350
rect 348048 508226 348368 508294
rect 348048 508170 348118 508226
rect 348174 508170 348242 508226
rect 348298 508170 348368 508226
rect 348048 508102 348368 508170
rect 348048 508046 348118 508102
rect 348174 508046 348242 508102
rect 348298 508046 348368 508102
rect 348048 507978 348368 508046
rect 348048 507922 348118 507978
rect 348174 507922 348242 507978
rect 348298 507922 348368 507978
rect 348048 507888 348368 507922
rect 378768 508350 379088 508384
rect 378768 508294 378838 508350
rect 378894 508294 378962 508350
rect 379018 508294 379088 508350
rect 378768 508226 379088 508294
rect 378768 508170 378838 508226
rect 378894 508170 378962 508226
rect 379018 508170 379088 508226
rect 378768 508102 379088 508170
rect 378768 508046 378838 508102
rect 378894 508046 378962 508102
rect 379018 508046 379088 508102
rect 378768 507978 379088 508046
rect 378768 507922 378838 507978
rect 378894 507922 378962 507978
rect 379018 507922 379088 507978
rect 378768 507888 379088 507922
rect 409488 508350 409808 508384
rect 409488 508294 409558 508350
rect 409614 508294 409682 508350
rect 409738 508294 409808 508350
rect 409488 508226 409808 508294
rect 409488 508170 409558 508226
rect 409614 508170 409682 508226
rect 409738 508170 409808 508226
rect 409488 508102 409808 508170
rect 409488 508046 409558 508102
rect 409614 508046 409682 508102
rect 409738 508046 409808 508102
rect 409488 507978 409808 508046
rect 409488 507922 409558 507978
rect 409614 507922 409682 507978
rect 409738 507922 409808 507978
rect 409488 507888 409808 507922
rect 440208 508350 440528 508384
rect 440208 508294 440278 508350
rect 440334 508294 440402 508350
rect 440458 508294 440528 508350
rect 440208 508226 440528 508294
rect 440208 508170 440278 508226
rect 440334 508170 440402 508226
rect 440458 508170 440528 508226
rect 440208 508102 440528 508170
rect 440208 508046 440278 508102
rect 440334 508046 440402 508102
rect 440458 508046 440528 508102
rect 440208 507978 440528 508046
rect 440208 507922 440278 507978
rect 440334 507922 440402 507978
rect 440458 507922 440528 507978
rect 440208 507888 440528 507922
rect 470928 508350 471248 508384
rect 470928 508294 470998 508350
rect 471054 508294 471122 508350
rect 471178 508294 471248 508350
rect 470928 508226 471248 508294
rect 470928 508170 470998 508226
rect 471054 508170 471122 508226
rect 471178 508170 471248 508226
rect 470928 508102 471248 508170
rect 470928 508046 470998 508102
rect 471054 508046 471122 508102
rect 471178 508046 471248 508102
rect 470928 507978 471248 508046
rect 470928 507922 470998 507978
rect 471054 507922 471122 507978
rect 471178 507922 471248 507978
rect 470928 507888 471248 507922
rect 501648 508350 501968 508384
rect 501648 508294 501718 508350
rect 501774 508294 501842 508350
rect 501898 508294 501968 508350
rect 501648 508226 501968 508294
rect 501648 508170 501718 508226
rect 501774 508170 501842 508226
rect 501898 508170 501968 508226
rect 501648 508102 501968 508170
rect 501648 508046 501718 508102
rect 501774 508046 501842 508102
rect 501898 508046 501968 508102
rect 501648 507978 501968 508046
rect 501648 507922 501718 507978
rect 501774 507922 501842 507978
rect 501898 507922 501968 507978
rect 501648 507888 501968 507922
rect 532368 508350 532688 508384
rect 532368 508294 532438 508350
rect 532494 508294 532562 508350
rect 532618 508294 532688 508350
rect 532368 508226 532688 508294
rect 532368 508170 532438 508226
rect 532494 508170 532562 508226
rect 532618 508170 532688 508226
rect 532368 508102 532688 508170
rect 532368 508046 532438 508102
rect 532494 508046 532562 508102
rect 532618 508046 532688 508102
rect 532368 507978 532688 508046
rect 532368 507922 532438 507978
rect 532494 507922 532562 507978
rect 532618 507922 532688 507978
rect 532368 507888 532688 507922
rect 209808 496350 210128 496384
rect 209808 496294 209878 496350
rect 209934 496294 210002 496350
rect 210058 496294 210128 496350
rect 209808 496226 210128 496294
rect 209808 496170 209878 496226
rect 209934 496170 210002 496226
rect 210058 496170 210128 496226
rect 209808 496102 210128 496170
rect 209808 496046 209878 496102
rect 209934 496046 210002 496102
rect 210058 496046 210128 496102
rect 209808 495978 210128 496046
rect 209808 495922 209878 495978
rect 209934 495922 210002 495978
rect 210058 495922 210128 495978
rect 209808 495888 210128 495922
rect 240528 496350 240848 496384
rect 240528 496294 240598 496350
rect 240654 496294 240722 496350
rect 240778 496294 240848 496350
rect 240528 496226 240848 496294
rect 240528 496170 240598 496226
rect 240654 496170 240722 496226
rect 240778 496170 240848 496226
rect 240528 496102 240848 496170
rect 240528 496046 240598 496102
rect 240654 496046 240722 496102
rect 240778 496046 240848 496102
rect 240528 495978 240848 496046
rect 240528 495922 240598 495978
rect 240654 495922 240722 495978
rect 240778 495922 240848 495978
rect 240528 495888 240848 495922
rect 271248 496350 271568 496384
rect 271248 496294 271318 496350
rect 271374 496294 271442 496350
rect 271498 496294 271568 496350
rect 271248 496226 271568 496294
rect 271248 496170 271318 496226
rect 271374 496170 271442 496226
rect 271498 496170 271568 496226
rect 271248 496102 271568 496170
rect 271248 496046 271318 496102
rect 271374 496046 271442 496102
rect 271498 496046 271568 496102
rect 271248 495978 271568 496046
rect 271248 495922 271318 495978
rect 271374 495922 271442 495978
rect 271498 495922 271568 495978
rect 271248 495888 271568 495922
rect 301968 496350 302288 496384
rect 301968 496294 302038 496350
rect 302094 496294 302162 496350
rect 302218 496294 302288 496350
rect 301968 496226 302288 496294
rect 301968 496170 302038 496226
rect 302094 496170 302162 496226
rect 302218 496170 302288 496226
rect 301968 496102 302288 496170
rect 301968 496046 302038 496102
rect 302094 496046 302162 496102
rect 302218 496046 302288 496102
rect 301968 495978 302288 496046
rect 301968 495922 302038 495978
rect 302094 495922 302162 495978
rect 302218 495922 302288 495978
rect 301968 495888 302288 495922
rect 332688 496350 333008 496384
rect 332688 496294 332758 496350
rect 332814 496294 332882 496350
rect 332938 496294 333008 496350
rect 332688 496226 333008 496294
rect 332688 496170 332758 496226
rect 332814 496170 332882 496226
rect 332938 496170 333008 496226
rect 332688 496102 333008 496170
rect 332688 496046 332758 496102
rect 332814 496046 332882 496102
rect 332938 496046 333008 496102
rect 332688 495978 333008 496046
rect 332688 495922 332758 495978
rect 332814 495922 332882 495978
rect 332938 495922 333008 495978
rect 332688 495888 333008 495922
rect 363408 496350 363728 496384
rect 363408 496294 363478 496350
rect 363534 496294 363602 496350
rect 363658 496294 363728 496350
rect 363408 496226 363728 496294
rect 363408 496170 363478 496226
rect 363534 496170 363602 496226
rect 363658 496170 363728 496226
rect 363408 496102 363728 496170
rect 363408 496046 363478 496102
rect 363534 496046 363602 496102
rect 363658 496046 363728 496102
rect 363408 495978 363728 496046
rect 363408 495922 363478 495978
rect 363534 495922 363602 495978
rect 363658 495922 363728 495978
rect 363408 495888 363728 495922
rect 394128 496350 394448 496384
rect 394128 496294 394198 496350
rect 394254 496294 394322 496350
rect 394378 496294 394448 496350
rect 394128 496226 394448 496294
rect 394128 496170 394198 496226
rect 394254 496170 394322 496226
rect 394378 496170 394448 496226
rect 394128 496102 394448 496170
rect 394128 496046 394198 496102
rect 394254 496046 394322 496102
rect 394378 496046 394448 496102
rect 394128 495978 394448 496046
rect 394128 495922 394198 495978
rect 394254 495922 394322 495978
rect 394378 495922 394448 495978
rect 394128 495888 394448 495922
rect 424848 496350 425168 496384
rect 424848 496294 424918 496350
rect 424974 496294 425042 496350
rect 425098 496294 425168 496350
rect 424848 496226 425168 496294
rect 424848 496170 424918 496226
rect 424974 496170 425042 496226
rect 425098 496170 425168 496226
rect 424848 496102 425168 496170
rect 424848 496046 424918 496102
rect 424974 496046 425042 496102
rect 425098 496046 425168 496102
rect 424848 495978 425168 496046
rect 424848 495922 424918 495978
rect 424974 495922 425042 495978
rect 425098 495922 425168 495978
rect 424848 495888 425168 495922
rect 455568 496350 455888 496384
rect 455568 496294 455638 496350
rect 455694 496294 455762 496350
rect 455818 496294 455888 496350
rect 455568 496226 455888 496294
rect 455568 496170 455638 496226
rect 455694 496170 455762 496226
rect 455818 496170 455888 496226
rect 455568 496102 455888 496170
rect 455568 496046 455638 496102
rect 455694 496046 455762 496102
rect 455818 496046 455888 496102
rect 455568 495978 455888 496046
rect 455568 495922 455638 495978
rect 455694 495922 455762 495978
rect 455818 495922 455888 495978
rect 455568 495888 455888 495922
rect 486288 496350 486608 496384
rect 486288 496294 486358 496350
rect 486414 496294 486482 496350
rect 486538 496294 486608 496350
rect 486288 496226 486608 496294
rect 486288 496170 486358 496226
rect 486414 496170 486482 496226
rect 486538 496170 486608 496226
rect 486288 496102 486608 496170
rect 486288 496046 486358 496102
rect 486414 496046 486482 496102
rect 486538 496046 486608 496102
rect 486288 495978 486608 496046
rect 486288 495922 486358 495978
rect 486414 495922 486482 495978
rect 486538 495922 486608 495978
rect 486288 495888 486608 495922
rect 517008 496350 517328 496384
rect 517008 496294 517078 496350
rect 517134 496294 517202 496350
rect 517258 496294 517328 496350
rect 517008 496226 517328 496294
rect 517008 496170 517078 496226
rect 517134 496170 517202 496226
rect 517258 496170 517328 496226
rect 517008 496102 517328 496170
rect 517008 496046 517078 496102
rect 517134 496046 517202 496102
rect 517258 496046 517328 496102
rect 517008 495978 517328 496046
rect 517008 495922 517078 495978
rect 517134 495922 517202 495978
rect 517258 495922 517328 495978
rect 517008 495888 517328 495922
rect 194448 490350 194768 490384
rect 194448 490294 194518 490350
rect 194574 490294 194642 490350
rect 194698 490294 194768 490350
rect 194448 490226 194768 490294
rect 194448 490170 194518 490226
rect 194574 490170 194642 490226
rect 194698 490170 194768 490226
rect 194448 490102 194768 490170
rect 194448 490046 194518 490102
rect 194574 490046 194642 490102
rect 194698 490046 194768 490102
rect 194448 489978 194768 490046
rect 194448 489922 194518 489978
rect 194574 489922 194642 489978
rect 194698 489922 194768 489978
rect 194448 489888 194768 489922
rect 225168 490350 225488 490384
rect 225168 490294 225238 490350
rect 225294 490294 225362 490350
rect 225418 490294 225488 490350
rect 225168 490226 225488 490294
rect 225168 490170 225238 490226
rect 225294 490170 225362 490226
rect 225418 490170 225488 490226
rect 225168 490102 225488 490170
rect 225168 490046 225238 490102
rect 225294 490046 225362 490102
rect 225418 490046 225488 490102
rect 225168 489978 225488 490046
rect 225168 489922 225238 489978
rect 225294 489922 225362 489978
rect 225418 489922 225488 489978
rect 225168 489888 225488 489922
rect 255888 490350 256208 490384
rect 255888 490294 255958 490350
rect 256014 490294 256082 490350
rect 256138 490294 256208 490350
rect 255888 490226 256208 490294
rect 255888 490170 255958 490226
rect 256014 490170 256082 490226
rect 256138 490170 256208 490226
rect 255888 490102 256208 490170
rect 255888 490046 255958 490102
rect 256014 490046 256082 490102
rect 256138 490046 256208 490102
rect 255888 489978 256208 490046
rect 255888 489922 255958 489978
rect 256014 489922 256082 489978
rect 256138 489922 256208 489978
rect 255888 489888 256208 489922
rect 286608 490350 286928 490384
rect 286608 490294 286678 490350
rect 286734 490294 286802 490350
rect 286858 490294 286928 490350
rect 286608 490226 286928 490294
rect 286608 490170 286678 490226
rect 286734 490170 286802 490226
rect 286858 490170 286928 490226
rect 286608 490102 286928 490170
rect 286608 490046 286678 490102
rect 286734 490046 286802 490102
rect 286858 490046 286928 490102
rect 286608 489978 286928 490046
rect 286608 489922 286678 489978
rect 286734 489922 286802 489978
rect 286858 489922 286928 489978
rect 286608 489888 286928 489922
rect 317328 490350 317648 490384
rect 317328 490294 317398 490350
rect 317454 490294 317522 490350
rect 317578 490294 317648 490350
rect 317328 490226 317648 490294
rect 317328 490170 317398 490226
rect 317454 490170 317522 490226
rect 317578 490170 317648 490226
rect 317328 490102 317648 490170
rect 317328 490046 317398 490102
rect 317454 490046 317522 490102
rect 317578 490046 317648 490102
rect 317328 489978 317648 490046
rect 317328 489922 317398 489978
rect 317454 489922 317522 489978
rect 317578 489922 317648 489978
rect 317328 489888 317648 489922
rect 348048 490350 348368 490384
rect 348048 490294 348118 490350
rect 348174 490294 348242 490350
rect 348298 490294 348368 490350
rect 348048 490226 348368 490294
rect 348048 490170 348118 490226
rect 348174 490170 348242 490226
rect 348298 490170 348368 490226
rect 348048 490102 348368 490170
rect 348048 490046 348118 490102
rect 348174 490046 348242 490102
rect 348298 490046 348368 490102
rect 348048 489978 348368 490046
rect 348048 489922 348118 489978
rect 348174 489922 348242 489978
rect 348298 489922 348368 489978
rect 348048 489888 348368 489922
rect 378768 490350 379088 490384
rect 378768 490294 378838 490350
rect 378894 490294 378962 490350
rect 379018 490294 379088 490350
rect 378768 490226 379088 490294
rect 378768 490170 378838 490226
rect 378894 490170 378962 490226
rect 379018 490170 379088 490226
rect 378768 490102 379088 490170
rect 378768 490046 378838 490102
rect 378894 490046 378962 490102
rect 379018 490046 379088 490102
rect 378768 489978 379088 490046
rect 378768 489922 378838 489978
rect 378894 489922 378962 489978
rect 379018 489922 379088 489978
rect 378768 489888 379088 489922
rect 409488 490350 409808 490384
rect 409488 490294 409558 490350
rect 409614 490294 409682 490350
rect 409738 490294 409808 490350
rect 409488 490226 409808 490294
rect 409488 490170 409558 490226
rect 409614 490170 409682 490226
rect 409738 490170 409808 490226
rect 409488 490102 409808 490170
rect 409488 490046 409558 490102
rect 409614 490046 409682 490102
rect 409738 490046 409808 490102
rect 409488 489978 409808 490046
rect 409488 489922 409558 489978
rect 409614 489922 409682 489978
rect 409738 489922 409808 489978
rect 409488 489888 409808 489922
rect 440208 490350 440528 490384
rect 440208 490294 440278 490350
rect 440334 490294 440402 490350
rect 440458 490294 440528 490350
rect 440208 490226 440528 490294
rect 440208 490170 440278 490226
rect 440334 490170 440402 490226
rect 440458 490170 440528 490226
rect 440208 490102 440528 490170
rect 440208 490046 440278 490102
rect 440334 490046 440402 490102
rect 440458 490046 440528 490102
rect 440208 489978 440528 490046
rect 440208 489922 440278 489978
rect 440334 489922 440402 489978
rect 440458 489922 440528 489978
rect 440208 489888 440528 489922
rect 470928 490350 471248 490384
rect 470928 490294 470998 490350
rect 471054 490294 471122 490350
rect 471178 490294 471248 490350
rect 470928 490226 471248 490294
rect 470928 490170 470998 490226
rect 471054 490170 471122 490226
rect 471178 490170 471248 490226
rect 470928 490102 471248 490170
rect 470928 490046 470998 490102
rect 471054 490046 471122 490102
rect 471178 490046 471248 490102
rect 470928 489978 471248 490046
rect 470928 489922 470998 489978
rect 471054 489922 471122 489978
rect 471178 489922 471248 489978
rect 470928 489888 471248 489922
rect 501648 490350 501968 490384
rect 501648 490294 501718 490350
rect 501774 490294 501842 490350
rect 501898 490294 501968 490350
rect 501648 490226 501968 490294
rect 501648 490170 501718 490226
rect 501774 490170 501842 490226
rect 501898 490170 501968 490226
rect 501648 490102 501968 490170
rect 501648 490046 501718 490102
rect 501774 490046 501842 490102
rect 501898 490046 501968 490102
rect 501648 489978 501968 490046
rect 501648 489922 501718 489978
rect 501774 489922 501842 489978
rect 501898 489922 501968 489978
rect 501648 489888 501968 489922
rect 532368 490350 532688 490384
rect 532368 490294 532438 490350
rect 532494 490294 532562 490350
rect 532618 490294 532688 490350
rect 532368 490226 532688 490294
rect 532368 490170 532438 490226
rect 532494 490170 532562 490226
rect 532618 490170 532688 490226
rect 532368 490102 532688 490170
rect 532368 490046 532438 490102
rect 532494 490046 532562 490102
rect 532618 490046 532688 490102
rect 532368 489978 532688 490046
rect 532368 489922 532438 489978
rect 532494 489922 532562 489978
rect 532618 489922 532688 489978
rect 532368 489888 532688 489922
rect 209808 478350 210128 478384
rect 209808 478294 209878 478350
rect 209934 478294 210002 478350
rect 210058 478294 210128 478350
rect 209808 478226 210128 478294
rect 209808 478170 209878 478226
rect 209934 478170 210002 478226
rect 210058 478170 210128 478226
rect 209808 478102 210128 478170
rect 209808 478046 209878 478102
rect 209934 478046 210002 478102
rect 210058 478046 210128 478102
rect 209808 477978 210128 478046
rect 209808 477922 209878 477978
rect 209934 477922 210002 477978
rect 210058 477922 210128 477978
rect 209808 477888 210128 477922
rect 240528 478350 240848 478384
rect 240528 478294 240598 478350
rect 240654 478294 240722 478350
rect 240778 478294 240848 478350
rect 240528 478226 240848 478294
rect 240528 478170 240598 478226
rect 240654 478170 240722 478226
rect 240778 478170 240848 478226
rect 240528 478102 240848 478170
rect 240528 478046 240598 478102
rect 240654 478046 240722 478102
rect 240778 478046 240848 478102
rect 240528 477978 240848 478046
rect 240528 477922 240598 477978
rect 240654 477922 240722 477978
rect 240778 477922 240848 477978
rect 240528 477888 240848 477922
rect 271248 478350 271568 478384
rect 271248 478294 271318 478350
rect 271374 478294 271442 478350
rect 271498 478294 271568 478350
rect 271248 478226 271568 478294
rect 271248 478170 271318 478226
rect 271374 478170 271442 478226
rect 271498 478170 271568 478226
rect 271248 478102 271568 478170
rect 271248 478046 271318 478102
rect 271374 478046 271442 478102
rect 271498 478046 271568 478102
rect 271248 477978 271568 478046
rect 271248 477922 271318 477978
rect 271374 477922 271442 477978
rect 271498 477922 271568 477978
rect 271248 477888 271568 477922
rect 301968 478350 302288 478384
rect 301968 478294 302038 478350
rect 302094 478294 302162 478350
rect 302218 478294 302288 478350
rect 301968 478226 302288 478294
rect 301968 478170 302038 478226
rect 302094 478170 302162 478226
rect 302218 478170 302288 478226
rect 301968 478102 302288 478170
rect 301968 478046 302038 478102
rect 302094 478046 302162 478102
rect 302218 478046 302288 478102
rect 301968 477978 302288 478046
rect 301968 477922 302038 477978
rect 302094 477922 302162 477978
rect 302218 477922 302288 477978
rect 301968 477888 302288 477922
rect 332688 478350 333008 478384
rect 332688 478294 332758 478350
rect 332814 478294 332882 478350
rect 332938 478294 333008 478350
rect 332688 478226 333008 478294
rect 332688 478170 332758 478226
rect 332814 478170 332882 478226
rect 332938 478170 333008 478226
rect 332688 478102 333008 478170
rect 332688 478046 332758 478102
rect 332814 478046 332882 478102
rect 332938 478046 333008 478102
rect 332688 477978 333008 478046
rect 332688 477922 332758 477978
rect 332814 477922 332882 477978
rect 332938 477922 333008 477978
rect 332688 477888 333008 477922
rect 363408 478350 363728 478384
rect 363408 478294 363478 478350
rect 363534 478294 363602 478350
rect 363658 478294 363728 478350
rect 363408 478226 363728 478294
rect 363408 478170 363478 478226
rect 363534 478170 363602 478226
rect 363658 478170 363728 478226
rect 363408 478102 363728 478170
rect 363408 478046 363478 478102
rect 363534 478046 363602 478102
rect 363658 478046 363728 478102
rect 363408 477978 363728 478046
rect 363408 477922 363478 477978
rect 363534 477922 363602 477978
rect 363658 477922 363728 477978
rect 363408 477888 363728 477922
rect 394128 478350 394448 478384
rect 394128 478294 394198 478350
rect 394254 478294 394322 478350
rect 394378 478294 394448 478350
rect 394128 478226 394448 478294
rect 394128 478170 394198 478226
rect 394254 478170 394322 478226
rect 394378 478170 394448 478226
rect 394128 478102 394448 478170
rect 394128 478046 394198 478102
rect 394254 478046 394322 478102
rect 394378 478046 394448 478102
rect 394128 477978 394448 478046
rect 394128 477922 394198 477978
rect 394254 477922 394322 477978
rect 394378 477922 394448 477978
rect 394128 477888 394448 477922
rect 424848 478350 425168 478384
rect 424848 478294 424918 478350
rect 424974 478294 425042 478350
rect 425098 478294 425168 478350
rect 424848 478226 425168 478294
rect 424848 478170 424918 478226
rect 424974 478170 425042 478226
rect 425098 478170 425168 478226
rect 424848 478102 425168 478170
rect 424848 478046 424918 478102
rect 424974 478046 425042 478102
rect 425098 478046 425168 478102
rect 424848 477978 425168 478046
rect 424848 477922 424918 477978
rect 424974 477922 425042 477978
rect 425098 477922 425168 477978
rect 424848 477888 425168 477922
rect 455568 478350 455888 478384
rect 455568 478294 455638 478350
rect 455694 478294 455762 478350
rect 455818 478294 455888 478350
rect 455568 478226 455888 478294
rect 455568 478170 455638 478226
rect 455694 478170 455762 478226
rect 455818 478170 455888 478226
rect 455568 478102 455888 478170
rect 455568 478046 455638 478102
rect 455694 478046 455762 478102
rect 455818 478046 455888 478102
rect 455568 477978 455888 478046
rect 455568 477922 455638 477978
rect 455694 477922 455762 477978
rect 455818 477922 455888 477978
rect 455568 477888 455888 477922
rect 486288 478350 486608 478384
rect 486288 478294 486358 478350
rect 486414 478294 486482 478350
rect 486538 478294 486608 478350
rect 486288 478226 486608 478294
rect 486288 478170 486358 478226
rect 486414 478170 486482 478226
rect 486538 478170 486608 478226
rect 486288 478102 486608 478170
rect 486288 478046 486358 478102
rect 486414 478046 486482 478102
rect 486538 478046 486608 478102
rect 486288 477978 486608 478046
rect 486288 477922 486358 477978
rect 486414 477922 486482 477978
rect 486538 477922 486608 477978
rect 486288 477888 486608 477922
rect 517008 478350 517328 478384
rect 517008 478294 517078 478350
rect 517134 478294 517202 478350
rect 517258 478294 517328 478350
rect 517008 478226 517328 478294
rect 517008 478170 517078 478226
rect 517134 478170 517202 478226
rect 517258 478170 517328 478226
rect 517008 478102 517328 478170
rect 517008 478046 517078 478102
rect 517134 478046 517202 478102
rect 517258 478046 517328 478102
rect 517008 477978 517328 478046
rect 517008 477922 517078 477978
rect 517134 477922 517202 477978
rect 517258 477922 517328 477978
rect 517008 477888 517328 477922
rect 194448 472350 194768 472384
rect 194448 472294 194518 472350
rect 194574 472294 194642 472350
rect 194698 472294 194768 472350
rect 194448 472226 194768 472294
rect 194448 472170 194518 472226
rect 194574 472170 194642 472226
rect 194698 472170 194768 472226
rect 194448 472102 194768 472170
rect 194448 472046 194518 472102
rect 194574 472046 194642 472102
rect 194698 472046 194768 472102
rect 194448 471978 194768 472046
rect 194448 471922 194518 471978
rect 194574 471922 194642 471978
rect 194698 471922 194768 471978
rect 194448 471888 194768 471922
rect 225168 472350 225488 472384
rect 225168 472294 225238 472350
rect 225294 472294 225362 472350
rect 225418 472294 225488 472350
rect 225168 472226 225488 472294
rect 225168 472170 225238 472226
rect 225294 472170 225362 472226
rect 225418 472170 225488 472226
rect 225168 472102 225488 472170
rect 225168 472046 225238 472102
rect 225294 472046 225362 472102
rect 225418 472046 225488 472102
rect 225168 471978 225488 472046
rect 225168 471922 225238 471978
rect 225294 471922 225362 471978
rect 225418 471922 225488 471978
rect 225168 471888 225488 471922
rect 255888 472350 256208 472384
rect 255888 472294 255958 472350
rect 256014 472294 256082 472350
rect 256138 472294 256208 472350
rect 255888 472226 256208 472294
rect 255888 472170 255958 472226
rect 256014 472170 256082 472226
rect 256138 472170 256208 472226
rect 255888 472102 256208 472170
rect 255888 472046 255958 472102
rect 256014 472046 256082 472102
rect 256138 472046 256208 472102
rect 255888 471978 256208 472046
rect 255888 471922 255958 471978
rect 256014 471922 256082 471978
rect 256138 471922 256208 471978
rect 255888 471888 256208 471922
rect 286608 472350 286928 472384
rect 286608 472294 286678 472350
rect 286734 472294 286802 472350
rect 286858 472294 286928 472350
rect 286608 472226 286928 472294
rect 286608 472170 286678 472226
rect 286734 472170 286802 472226
rect 286858 472170 286928 472226
rect 286608 472102 286928 472170
rect 286608 472046 286678 472102
rect 286734 472046 286802 472102
rect 286858 472046 286928 472102
rect 286608 471978 286928 472046
rect 286608 471922 286678 471978
rect 286734 471922 286802 471978
rect 286858 471922 286928 471978
rect 286608 471888 286928 471922
rect 317328 472350 317648 472384
rect 317328 472294 317398 472350
rect 317454 472294 317522 472350
rect 317578 472294 317648 472350
rect 317328 472226 317648 472294
rect 317328 472170 317398 472226
rect 317454 472170 317522 472226
rect 317578 472170 317648 472226
rect 317328 472102 317648 472170
rect 317328 472046 317398 472102
rect 317454 472046 317522 472102
rect 317578 472046 317648 472102
rect 317328 471978 317648 472046
rect 317328 471922 317398 471978
rect 317454 471922 317522 471978
rect 317578 471922 317648 471978
rect 317328 471888 317648 471922
rect 348048 472350 348368 472384
rect 348048 472294 348118 472350
rect 348174 472294 348242 472350
rect 348298 472294 348368 472350
rect 348048 472226 348368 472294
rect 348048 472170 348118 472226
rect 348174 472170 348242 472226
rect 348298 472170 348368 472226
rect 348048 472102 348368 472170
rect 348048 472046 348118 472102
rect 348174 472046 348242 472102
rect 348298 472046 348368 472102
rect 348048 471978 348368 472046
rect 348048 471922 348118 471978
rect 348174 471922 348242 471978
rect 348298 471922 348368 471978
rect 348048 471888 348368 471922
rect 378768 472350 379088 472384
rect 378768 472294 378838 472350
rect 378894 472294 378962 472350
rect 379018 472294 379088 472350
rect 378768 472226 379088 472294
rect 378768 472170 378838 472226
rect 378894 472170 378962 472226
rect 379018 472170 379088 472226
rect 378768 472102 379088 472170
rect 378768 472046 378838 472102
rect 378894 472046 378962 472102
rect 379018 472046 379088 472102
rect 378768 471978 379088 472046
rect 378768 471922 378838 471978
rect 378894 471922 378962 471978
rect 379018 471922 379088 471978
rect 378768 471888 379088 471922
rect 409488 472350 409808 472384
rect 409488 472294 409558 472350
rect 409614 472294 409682 472350
rect 409738 472294 409808 472350
rect 409488 472226 409808 472294
rect 409488 472170 409558 472226
rect 409614 472170 409682 472226
rect 409738 472170 409808 472226
rect 409488 472102 409808 472170
rect 409488 472046 409558 472102
rect 409614 472046 409682 472102
rect 409738 472046 409808 472102
rect 409488 471978 409808 472046
rect 409488 471922 409558 471978
rect 409614 471922 409682 471978
rect 409738 471922 409808 471978
rect 409488 471888 409808 471922
rect 440208 472350 440528 472384
rect 440208 472294 440278 472350
rect 440334 472294 440402 472350
rect 440458 472294 440528 472350
rect 440208 472226 440528 472294
rect 440208 472170 440278 472226
rect 440334 472170 440402 472226
rect 440458 472170 440528 472226
rect 440208 472102 440528 472170
rect 440208 472046 440278 472102
rect 440334 472046 440402 472102
rect 440458 472046 440528 472102
rect 440208 471978 440528 472046
rect 440208 471922 440278 471978
rect 440334 471922 440402 471978
rect 440458 471922 440528 471978
rect 440208 471888 440528 471922
rect 470928 472350 471248 472384
rect 470928 472294 470998 472350
rect 471054 472294 471122 472350
rect 471178 472294 471248 472350
rect 470928 472226 471248 472294
rect 470928 472170 470998 472226
rect 471054 472170 471122 472226
rect 471178 472170 471248 472226
rect 470928 472102 471248 472170
rect 470928 472046 470998 472102
rect 471054 472046 471122 472102
rect 471178 472046 471248 472102
rect 470928 471978 471248 472046
rect 470928 471922 470998 471978
rect 471054 471922 471122 471978
rect 471178 471922 471248 471978
rect 470928 471888 471248 471922
rect 501648 472350 501968 472384
rect 501648 472294 501718 472350
rect 501774 472294 501842 472350
rect 501898 472294 501968 472350
rect 501648 472226 501968 472294
rect 501648 472170 501718 472226
rect 501774 472170 501842 472226
rect 501898 472170 501968 472226
rect 501648 472102 501968 472170
rect 501648 472046 501718 472102
rect 501774 472046 501842 472102
rect 501898 472046 501968 472102
rect 501648 471978 501968 472046
rect 501648 471922 501718 471978
rect 501774 471922 501842 471978
rect 501898 471922 501968 471978
rect 501648 471888 501968 471922
rect 532368 472350 532688 472384
rect 532368 472294 532438 472350
rect 532494 472294 532562 472350
rect 532618 472294 532688 472350
rect 532368 472226 532688 472294
rect 532368 472170 532438 472226
rect 532494 472170 532562 472226
rect 532618 472170 532688 472226
rect 532368 472102 532688 472170
rect 532368 472046 532438 472102
rect 532494 472046 532562 472102
rect 532618 472046 532688 472102
rect 532368 471978 532688 472046
rect 532368 471922 532438 471978
rect 532494 471922 532562 471978
rect 532618 471922 532688 471978
rect 532368 471888 532688 471922
rect 209808 460350 210128 460384
rect 209808 460294 209878 460350
rect 209934 460294 210002 460350
rect 210058 460294 210128 460350
rect 209808 460226 210128 460294
rect 209808 460170 209878 460226
rect 209934 460170 210002 460226
rect 210058 460170 210128 460226
rect 209808 460102 210128 460170
rect 209808 460046 209878 460102
rect 209934 460046 210002 460102
rect 210058 460046 210128 460102
rect 209808 459978 210128 460046
rect 209808 459922 209878 459978
rect 209934 459922 210002 459978
rect 210058 459922 210128 459978
rect 209808 459888 210128 459922
rect 240528 460350 240848 460384
rect 240528 460294 240598 460350
rect 240654 460294 240722 460350
rect 240778 460294 240848 460350
rect 240528 460226 240848 460294
rect 240528 460170 240598 460226
rect 240654 460170 240722 460226
rect 240778 460170 240848 460226
rect 240528 460102 240848 460170
rect 240528 460046 240598 460102
rect 240654 460046 240722 460102
rect 240778 460046 240848 460102
rect 240528 459978 240848 460046
rect 240528 459922 240598 459978
rect 240654 459922 240722 459978
rect 240778 459922 240848 459978
rect 240528 459888 240848 459922
rect 271248 460350 271568 460384
rect 271248 460294 271318 460350
rect 271374 460294 271442 460350
rect 271498 460294 271568 460350
rect 271248 460226 271568 460294
rect 271248 460170 271318 460226
rect 271374 460170 271442 460226
rect 271498 460170 271568 460226
rect 271248 460102 271568 460170
rect 271248 460046 271318 460102
rect 271374 460046 271442 460102
rect 271498 460046 271568 460102
rect 271248 459978 271568 460046
rect 271248 459922 271318 459978
rect 271374 459922 271442 459978
rect 271498 459922 271568 459978
rect 271248 459888 271568 459922
rect 301968 460350 302288 460384
rect 301968 460294 302038 460350
rect 302094 460294 302162 460350
rect 302218 460294 302288 460350
rect 301968 460226 302288 460294
rect 301968 460170 302038 460226
rect 302094 460170 302162 460226
rect 302218 460170 302288 460226
rect 301968 460102 302288 460170
rect 301968 460046 302038 460102
rect 302094 460046 302162 460102
rect 302218 460046 302288 460102
rect 301968 459978 302288 460046
rect 301968 459922 302038 459978
rect 302094 459922 302162 459978
rect 302218 459922 302288 459978
rect 301968 459888 302288 459922
rect 332688 460350 333008 460384
rect 332688 460294 332758 460350
rect 332814 460294 332882 460350
rect 332938 460294 333008 460350
rect 332688 460226 333008 460294
rect 332688 460170 332758 460226
rect 332814 460170 332882 460226
rect 332938 460170 333008 460226
rect 332688 460102 333008 460170
rect 332688 460046 332758 460102
rect 332814 460046 332882 460102
rect 332938 460046 333008 460102
rect 332688 459978 333008 460046
rect 332688 459922 332758 459978
rect 332814 459922 332882 459978
rect 332938 459922 333008 459978
rect 332688 459888 333008 459922
rect 363408 460350 363728 460384
rect 363408 460294 363478 460350
rect 363534 460294 363602 460350
rect 363658 460294 363728 460350
rect 363408 460226 363728 460294
rect 363408 460170 363478 460226
rect 363534 460170 363602 460226
rect 363658 460170 363728 460226
rect 363408 460102 363728 460170
rect 363408 460046 363478 460102
rect 363534 460046 363602 460102
rect 363658 460046 363728 460102
rect 363408 459978 363728 460046
rect 363408 459922 363478 459978
rect 363534 459922 363602 459978
rect 363658 459922 363728 459978
rect 363408 459888 363728 459922
rect 394128 460350 394448 460384
rect 394128 460294 394198 460350
rect 394254 460294 394322 460350
rect 394378 460294 394448 460350
rect 394128 460226 394448 460294
rect 394128 460170 394198 460226
rect 394254 460170 394322 460226
rect 394378 460170 394448 460226
rect 394128 460102 394448 460170
rect 394128 460046 394198 460102
rect 394254 460046 394322 460102
rect 394378 460046 394448 460102
rect 394128 459978 394448 460046
rect 394128 459922 394198 459978
rect 394254 459922 394322 459978
rect 394378 459922 394448 459978
rect 394128 459888 394448 459922
rect 424848 460350 425168 460384
rect 424848 460294 424918 460350
rect 424974 460294 425042 460350
rect 425098 460294 425168 460350
rect 424848 460226 425168 460294
rect 424848 460170 424918 460226
rect 424974 460170 425042 460226
rect 425098 460170 425168 460226
rect 424848 460102 425168 460170
rect 424848 460046 424918 460102
rect 424974 460046 425042 460102
rect 425098 460046 425168 460102
rect 424848 459978 425168 460046
rect 424848 459922 424918 459978
rect 424974 459922 425042 459978
rect 425098 459922 425168 459978
rect 424848 459888 425168 459922
rect 455568 460350 455888 460384
rect 455568 460294 455638 460350
rect 455694 460294 455762 460350
rect 455818 460294 455888 460350
rect 455568 460226 455888 460294
rect 455568 460170 455638 460226
rect 455694 460170 455762 460226
rect 455818 460170 455888 460226
rect 455568 460102 455888 460170
rect 455568 460046 455638 460102
rect 455694 460046 455762 460102
rect 455818 460046 455888 460102
rect 455568 459978 455888 460046
rect 455568 459922 455638 459978
rect 455694 459922 455762 459978
rect 455818 459922 455888 459978
rect 455568 459888 455888 459922
rect 486288 460350 486608 460384
rect 486288 460294 486358 460350
rect 486414 460294 486482 460350
rect 486538 460294 486608 460350
rect 486288 460226 486608 460294
rect 486288 460170 486358 460226
rect 486414 460170 486482 460226
rect 486538 460170 486608 460226
rect 486288 460102 486608 460170
rect 486288 460046 486358 460102
rect 486414 460046 486482 460102
rect 486538 460046 486608 460102
rect 486288 459978 486608 460046
rect 486288 459922 486358 459978
rect 486414 459922 486482 459978
rect 486538 459922 486608 459978
rect 486288 459888 486608 459922
rect 517008 460350 517328 460384
rect 517008 460294 517078 460350
rect 517134 460294 517202 460350
rect 517258 460294 517328 460350
rect 517008 460226 517328 460294
rect 517008 460170 517078 460226
rect 517134 460170 517202 460226
rect 517258 460170 517328 460226
rect 517008 460102 517328 460170
rect 517008 460046 517078 460102
rect 517134 460046 517202 460102
rect 517258 460046 517328 460102
rect 517008 459978 517328 460046
rect 517008 459922 517078 459978
rect 517134 459922 517202 459978
rect 517258 459922 517328 459978
rect 517008 459888 517328 459922
rect 194448 454350 194768 454384
rect 194448 454294 194518 454350
rect 194574 454294 194642 454350
rect 194698 454294 194768 454350
rect 194448 454226 194768 454294
rect 194448 454170 194518 454226
rect 194574 454170 194642 454226
rect 194698 454170 194768 454226
rect 194448 454102 194768 454170
rect 194448 454046 194518 454102
rect 194574 454046 194642 454102
rect 194698 454046 194768 454102
rect 194448 453978 194768 454046
rect 194448 453922 194518 453978
rect 194574 453922 194642 453978
rect 194698 453922 194768 453978
rect 194448 453888 194768 453922
rect 225168 454350 225488 454384
rect 225168 454294 225238 454350
rect 225294 454294 225362 454350
rect 225418 454294 225488 454350
rect 225168 454226 225488 454294
rect 225168 454170 225238 454226
rect 225294 454170 225362 454226
rect 225418 454170 225488 454226
rect 225168 454102 225488 454170
rect 225168 454046 225238 454102
rect 225294 454046 225362 454102
rect 225418 454046 225488 454102
rect 225168 453978 225488 454046
rect 225168 453922 225238 453978
rect 225294 453922 225362 453978
rect 225418 453922 225488 453978
rect 225168 453888 225488 453922
rect 255888 454350 256208 454384
rect 255888 454294 255958 454350
rect 256014 454294 256082 454350
rect 256138 454294 256208 454350
rect 255888 454226 256208 454294
rect 255888 454170 255958 454226
rect 256014 454170 256082 454226
rect 256138 454170 256208 454226
rect 255888 454102 256208 454170
rect 255888 454046 255958 454102
rect 256014 454046 256082 454102
rect 256138 454046 256208 454102
rect 255888 453978 256208 454046
rect 255888 453922 255958 453978
rect 256014 453922 256082 453978
rect 256138 453922 256208 453978
rect 255888 453888 256208 453922
rect 286608 454350 286928 454384
rect 286608 454294 286678 454350
rect 286734 454294 286802 454350
rect 286858 454294 286928 454350
rect 286608 454226 286928 454294
rect 286608 454170 286678 454226
rect 286734 454170 286802 454226
rect 286858 454170 286928 454226
rect 286608 454102 286928 454170
rect 286608 454046 286678 454102
rect 286734 454046 286802 454102
rect 286858 454046 286928 454102
rect 286608 453978 286928 454046
rect 286608 453922 286678 453978
rect 286734 453922 286802 453978
rect 286858 453922 286928 453978
rect 286608 453888 286928 453922
rect 317328 454350 317648 454384
rect 317328 454294 317398 454350
rect 317454 454294 317522 454350
rect 317578 454294 317648 454350
rect 317328 454226 317648 454294
rect 317328 454170 317398 454226
rect 317454 454170 317522 454226
rect 317578 454170 317648 454226
rect 317328 454102 317648 454170
rect 317328 454046 317398 454102
rect 317454 454046 317522 454102
rect 317578 454046 317648 454102
rect 317328 453978 317648 454046
rect 317328 453922 317398 453978
rect 317454 453922 317522 453978
rect 317578 453922 317648 453978
rect 317328 453888 317648 453922
rect 348048 454350 348368 454384
rect 348048 454294 348118 454350
rect 348174 454294 348242 454350
rect 348298 454294 348368 454350
rect 348048 454226 348368 454294
rect 348048 454170 348118 454226
rect 348174 454170 348242 454226
rect 348298 454170 348368 454226
rect 348048 454102 348368 454170
rect 348048 454046 348118 454102
rect 348174 454046 348242 454102
rect 348298 454046 348368 454102
rect 348048 453978 348368 454046
rect 348048 453922 348118 453978
rect 348174 453922 348242 453978
rect 348298 453922 348368 453978
rect 348048 453888 348368 453922
rect 378768 454350 379088 454384
rect 378768 454294 378838 454350
rect 378894 454294 378962 454350
rect 379018 454294 379088 454350
rect 378768 454226 379088 454294
rect 378768 454170 378838 454226
rect 378894 454170 378962 454226
rect 379018 454170 379088 454226
rect 378768 454102 379088 454170
rect 378768 454046 378838 454102
rect 378894 454046 378962 454102
rect 379018 454046 379088 454102
rect 378768 453978 379088 454046
rect 378768 453922 378838 453978
rect 378894 453922 378962 453978
rect 379018 453922 379088 453978
rect 378768 453888 379088 453922
rect 409488 454350 409808 454384
rect 409488 454294 409558 454350
rect 409614 454294 409682 454350
rect 409738 454294 409808 454350
rect 409488 454226 409808 454294
rect 409488 454170 409558 454226
rect 409614 454170 409682 454226
rect 409738 454170 409808 454226
rect 409488 454102 409808 454170
rect 409488 454046 409558 454102
rect 409614 454046 409682 454102
rect 409738 454046 409808 454102
rect 409488 453978 409808 454046
rect 409488 453922 409558 453978
rect 409614 453922 409682 453978
rect 409738 453922 409808 453978
rect 409488 453888 409808 453922
rect 440208 454350 440528 454384
rect 440208 454294 440278 454350
rect 440334 454294 440402 454350
rect 440458 454294 440528 454350
rect 440208 454226 440528 454294
rect 440208 454170 440278 454226
rect 440334 454170 440402 454226
rect 440458 454170 440528 454226
rect 440208 454102 440528 454170
rect 440208 454046 440278 454102
rect 440334 454046 440402 454102
rect 440458 454046 440528 454102
rect 440208 453978 440528 454046
rect 440208 453922 440278 453978
rect 440334 453922 440402 453978
rect 440458 453922 440528 453978
rect 440208 453888 440528 453922
rect 470928 454350 471248 454384
rect 470928 454294 470998 454350
rect 471054 454294 471122 454350
rect 471178 454294 471248 454350
rect 470928 454226 471248 454294
rect 470928 454170 470998 454226
rect 471054 454170 471122 454226
rect 471178 454170 471248 454226
rect 470928 454102 471248 454170
rect 470928 454046 470998 454102
rect 471054 454046 471122 454102
rect 471178 454046 471248 454102
rect 470928 453978 471248 454046
rect 470928 453922 470998 453978
rect 471054 453922 471122 453978
rect 471178 453922 471248 453978
rect 470928 453888 471248 453922
rect 501648 454350 501968 454384
rect 501648 454294 501718 454350
rect 501774 454294 501842 454350
rect 501898 454294 501968 454350
rect 501648 454226 501968 454294
rect 501648 454170 501718 454226
rect 501774 454170 501842 454226
rect 501898 454170 501968 454226
rect 501648 454102 501968 454170
rect 501648 454046 501718 454102
rect 501774 454046 501842 454102
rect 501898 454046 501968 454102
rect 501648 453978 501968 454046
rect 501648 453922 501718 453978
rect 501774 453922 501842 453978
rect 501898 453922 501968 453978
rect 501648 453888 501968 453922
rect 532368 454350 532688 454384
rect 532368 454294 532438 454350
rect 532494 454294 532562 454350
rect 532618 454294 532688 454350
rect 532368 454226 532688 454294
rect 532368 454170 532438 454226
rect 532494 454170 532562 454226
rect 532618 454170 532688 454226
rect 532368 454102 532688 454170
rect 532368 454046 532438 454102
rect 532494 454046 532562 454102
rect 532618 454046 532688 454102
rect 532368 453978 532688 454046
rect 532368 453922 532438 453978
rect 532494 453922 532562 453978
rect 532618 453922 532688 453978
rect 532368 453888 532688 453922
rect 209808 442350 210128 442384
rect 209808 442294 209878 442350
rect 209934 442294 210002 442350
rect 210058 442294 210128 442350
rect 209808 442226 210128 442294
rect 209808 442170 209878 442226
rect 209934 442170 210002 442226
rect 210058 442170 210128 442226
rect 209808 442102 210128 442170
rect 209808 442046 209878 442102
rect 209934 442046 210002 442102
rect 210058 442046 210128 442102
rect 209808 441978 210128 442046
rect 209808 441922 209878 441978
rect 209934 441922 210002 441978
rect 210058 441922 210128 441978
rect 209808 441888 210128 441922
rect 240528 442350 240848 442384
rect 240528 442294 240598 442350
rect 240654 442294 240722 442350
rect 240778 442294 240848 442350
rect 240528 442226 240848 442294
rect 240528 442170 240598 442226
rect 240654 442170 240722 442226
rect 240778 442170 240848 442226
rect 240528 442102 240848 442170
rect 240528 442046 240598 442102
rect 240654 442046 240722 442102
rect 240778 442046 240848 442102
rect 240528 441978 240848 442046
rect 240528 441922 240598 441978
rect 240654 441922 240722 441978
rect 240778 441922 240848 441978
rect 240528 441888 240848 441922
rect 271248 442350 271568 442384
rect 271248 442294 271318 442350
rect 271374 442294 271442 442350
rect 271498 442294 271568 442350
rect 271248 442226 271568 442294
rect 271248 442170 271318 442226
rect 271374 442170 271442 442226
rect 271498 442170 271568 442226
rect 271248 442102 271568 442170
rect 271248 442046 271318 442102
rect 271374 442046 271442 442102
rect 271498 442046 271568 442102
rect 271248 441978 271568 442046
rect 271248 441922 271318 441978
rect 271374 441922 271442 441978
rect 271498 441922 271568 441978
rect 271248 441888 271568 441922
rect 301968 442350 302288 442384
rect 301968 442294 302038 442350
rect 302094 442294 302162 442350
rect 302218 442294 302288 442350
rect 301968 442226 302288 442294
rect 301968 442170 302038 442226
rect 302094 442170 302162 442226
rect 302218 442170 302288 442226
rect 301968 442102 302288 442170
rect 301968 442046 302038 442102
rect 302094 442046 302162 442102
rect 302218 442046 302288 442102
rect 301968 441978 302288 442046
rect 301968 441922 302038 441978
rect 302094 441922 302162 441978
rect 302218 441922 302288 441978
rect 301968 441888 302288 441922
rect 332688 442350 333008 442384
rect 332688 442294 332758 442350
rect 332814 442294 332882 442350
rect 332938 442294 333008 442350
rect 332688 442226 333008 442294
rect 332688 442170 332758 442226
rect 332814 442170 332882 442226
rect 332938 442170 333008 442226
rect 332688 442102 333008 442170
rect 332688 442046 332758 442102
rect 332814 442046 332882 442102
rect 332938 442046 333008 442102
rect 332688 441978 333008 442046
rect 332688 441922 332758 441978
rect 332814 441922 332882 441978
rect 332938 441922 333008 441978
rect 332688 441888 333008 441922
rect 363408 442350 363728 442384
rect 363408 442294 363478 442350
rect 363534 442294 363602 442350
rect 363658 442294 363728 442350
rect 363408 442226 363728 442294
rect 363408 442170 363478 442226
rect 363534 442170 363602 442226
rect 363658 442170 363728 442226
rect 363408 442102 363728 442170
rect 363408 442046 363478 442102
rect 363534 442046 363602 442102
rect 363658 442046 363728 442102
rect 363408 441978 363728 442046
rect 363408 441922 363478 441978
rect 363534 441922 363602 441978
rect 363658 441922 363728 441978
rect 363408 441888 363728 441922
rect 394128 442350 394448 442384
rect 394128 442294 394198 442350
rect 394254 442294 394322 442350
rect 394378 442294 394448 442350
rect 394128 442226 394448 442294
rect 394128 442170 394198 442226
rect 394254 442170 394322 442226
rect 394378 442170 394448 442226
rect 394128 442102 394448 442170
rect 394128 442046 394198 442102
rect 394254 442046 394322 442102
rect 394378 442046 394448 442102
rect 394128 441978 394448 442046
rect 394128 441922 394198 441978
rect 394254 441922 394322 441978
rect 394378 441922 394448 441978
rect 394128 441888 394448 441922
rect 424848 442350 425168 442384
rect 424848 442294 424918 442350
rect 424974 442294 425042 442350
rect 425098 442294 425168 442350
rect 424848 442226 425168 442294
rect 424848 442170 424918 442226
rect 424974 442170 425042 442226
rect 425098 442170 425168 442226
rect 424848 442102 425168 442170
rect 424848 442046 424918 442102
rect 424974 442046 425042 442102
rect 425098 442046 425168 442102
rect 424848 441978 425168 442046
rect 424848 441922 424918 441978
rect 424974 441922 425042 441978
rect 425098 441922 425168 441978
rect 424848 441888 425168 441922
rect 455568 442350 455888 442384
rect 455568 442294 455638 442350
rect 455694 442294 455762 442350
rect 455818 442294 455888 442350
rect 455568 442226 455888 442294
rect 455568 442170 455638 442226
rect 455694 442170 455762 442226
rect 455818 442170 455888 442226
rect 455568 442102 455888 442170
rect 455568 442046 455638 442102
rect 455694 442046 455762 442102
rect 455818 442046 455888 442102
rect 455568 441978 455888 442046
rect 455568 441922 455638 441978
rect 455694 441922 455762 441978
rect 455818 441922 455888 441978
rect 455568 441888 455888 441922
rect 486288 442350 486608 442384
rect 486288 442294 486358 442350
rect 486414 442294 486482 442350
rect 486538 442294 486608 442350
rect 486288 442226 486608 442294
rect 486288 442170 486358 442226
rect 486414 442170 486482 442226
rect 486538 442170 486608 442226
rect 486288 442102 486608 442170
rect 486288 442046 486358 442102
rect 486414 442046 486482 442102
rect 486538 442046 486608 442102
rect 486288 441978 486608 442046
rect 486288 441922 486358 441978
rect 486414 441922 486482 441978
rect 486538 441922 486608 441978
rect 486288 441888 486608 441922
rect 517008 442350 517328 442384
rect 517008 442294 517078 442350
rect 517134 442294 517202 442350
rect 517258 442294 517328 442350
rect 517008 442226 517328 442294
rect 517008 442170 517078 442226
rect 517134 442170 517202 442226
rect 517258 442170 517328 442226
rect 517008 442102 517328 442170
rect 517008 442046 517078 442102
rect 517134 442046 517202 442102
rect 517258 442046 517328 442102
rect 517008 441978 517328 442046
rect 517008 441922 517078 441978
rect 517134 441922 517202 441978
rect 517258 441922 517328 441978
rect 517008 441888 517328 441922
rect 194448 436350 194768 436384
rect 194448 436294 194518 436350
rect 194574 436294 194642 436350
rect 194698 436294 194768 436350
rect 194448 436226 194768 436294
rect 194448 436170 194518 436226
rect 194574 436170 194642 436226
rect 194698 436170 194768 436226
rect 194448 436102 194768 436170
rect 194448 436046 194518 436102
rect 194574 436046 194642 436102
rect 194698 436046 194768 436102
rect 194448 435978 194768 436046
rect 194448 435922 194518 435978
rect 194574 435922 194642 435978
rect 194698 435922 194768 435978
rect 194448 435888 194768 435922
rect 225168 436350 225488 436384
rect 225168 436294 225238 436350
rect 225294 436294 225362 436350
rect 225418 436294 225488 436350
rect 225168 436226 225488 436294
rect 225168 436170 225238 436226
rect 225294 436170 225362 436226
rect 225418 436170 225488 436226
rect 225168 436102 225488 436170
rect 225168 436046 225238 436102
rect 225294 436046 225362 436102
rect 225418 436046 225488 436102
rect 225168 435978 225488 436046
rect 225168 435922 225238 435978
rect 225294 435922 225362 435978
rect 225418 435922 225488 435978
rect 225168 435888 225488 435922
rect 255888 436350 256208 436384
rect 255888 436294 255958 436350
rect 256014 436294 256082 436350
rect 256138 436294 256208 436350
rect 255888 436226 256208 436294
rect 255888 436170 255958 436226
rect 256014 436170 256082 436226
rect 256138 436170 256208 436226
rect 255888 436102 256208 436170
rect 255888 436046 255958 436102
rect 256014 436046 256082 436102
rect 256138 436046 256208 436102
rect 255888 435978 256208 436046
rect 255888 435922 255958 435978
rect 256014 435922 256082 435978
rect 256138 435922 256208 435978
rect 255888 435888 256208 435922
rect 286608 436350 286928 436384
rect 286608 436294 286678 436350
rect 286734 436294 286802 436350
rect 286858 436294 286928 436350
rect 286608 436226 286928 436294
rect 286608 436170 286678 436226
rect 286734 436170 286802 436226
rect 286858 436170 286928 436226
rect 286608 436102 286928 436170
rect 286608 436046 286678 436102
rect 286734 436046 286802 436102
rect 286858 436046 286928 436102
rect 286608 435978 286928 436046
rect 286608 435922 286678 435978
rect 286734 435922 286802 435978
rect 286858 435922 286928 435978
rect 286608 435888 286928 435922
rect 317328 436350 317648 436384
rect 317328 436294 317398 436350
rect 317454 436294 317522 436350
rect 317578 436294 317648 436350
rect 317328 436226 317648 436294
rect 317328 436170 317398 436226
rect 317454 436170 317522 436226
rect 317578 436170 317648 436226
rect 317328 436102 317648 436170
rect 317328 436046 317398 436102
rect 317454 436046 317522 436102
rect 317578 436046 317648 436102
rect 317328 435978 317648 436046
rect 317328 435922 317398 435978
rect 317454 435922 317522 435978
rect 317578 435922 317648 435978
rect 317328 435888 317648 435922
rect 348048 436350 348368 436384
rect 348048 436294 348118 436350
rect 348174 436294 348242 436350
rect 348298 436294 348368 436350
rect 348048 436226 348368 436294
rect 348048 436170 348118 436226
rect 348174 436170 348242 436226
rect 348298 436170 348368 436226
rect 348048 436102 348368 436170
rect 348048 436046 348118 436102
rect 348174 436046 348242 436102
rect 348298 436046 348368 436102
rect 348048 435978 348368 436046
rect 348048 435922 348118 435978
rect 348174 435922 348242 435978
rect 348298 435922 348368 435978
rect 348048 435888 348368 435922
rect 378768 436350 379088 436384
rect 378768 436294 378838 436350
rect 378894 436294 378962 436350
rect 379018 436294 379088 436350
rect 378768 436226 379088 436294
rect 378768 436170 378838 436226
rect 378894 436170 378962 436226
rect 379018 436170 379088 436226
rect 378768 436102 379088 436170
rect 378768 436046 378838 436102
rect 378894 436046 378962 436102
rect 379018 436046 379088 436102
rect 378768 435978 379088 436046
rect 378768 435922 378838 435978
rect 378894 435922 378962 435978
rect 379018 435922 379088 435978
rect 378768 435888 379088 435922
rect 409488 436350 409808 436384
rect 409488 436294 409558 436350
rect 409614 436294 409682 436350
rect 409738 436294 409808 436350
rect 409488 436226 409808 436294
rect 409488 436170 409558 436226
rect 409614 436170 409682 436226
rect 409738 436170 409808 436226
rect 409488 436102 409808 436170
rect 409488 436046 409558 436102
rect 409614 436046 409682 436102
rect 409738 436046 409808 436102
rect 409488 435978 409808 436046
rect 409488 435922 409558 435978
rect 409614 435922 409682 435978
rect 409738 435922 409808 435978
rect 409488 435888 409808 435922
rect 440208 436350 440528 436384
rect 440208 436294 440278 436350
rect 440334 436294 440402 436350
rect 440458 436294 440528 436350
rect 440208 436226 440528 436294
rect 440208 436170 440278 436226
rect 440334 436170 440402 436226
rect 440458 436170 440528 436226
rect 440208 436102 440528 436170
rect 440208 436046 440278 436102
rect 440334 436046 440402 436102
rect 440458 436046 440528 436102
rect 440208 435978 440528 436046
rect 440208 435922 440278 435978
rect 440334 435922 440402 435978
rect 440458 435922 440528 435978
rect 440208 435888 440528 435922
rect 470928 436350 471248 436384
rect 470928 436294 470998 436350
rect 471054 436294 471122 436350
rect 471178 436294 471248 436350
rect 470928 436226 471248 436294
rect 470928 436170 470998 436226
rect 471054 436170 471122 436226
rect 471178 436170 471248 436226
rect 470928 436102 471248 436170
rect 470928 436046 470998 436102
rect 471054 436046 471122 436102
rect 471178 436046 471248 436102
rect 470928 435978 471248 436046
rect 470928 435922 470998 435978
rect 471054 435922 471122 435978
rect 471178 435922 471248 435978
rect 470928 435888 471248 435922
rect 501648 436350 501968 436384
rect 501648 436294 501718 436350
rect 501774 436294 501842 436350
rect 501898 436294 501968 436350
rect 501648 436226 501968 436294
rect 501648 436170 501718 436226
rect 501774 436170 501842 436226
rect 501898 436170 501968 436226
rect 501648 436102 501968 436170
rect 501648 436046 501718 436102
rect 501774 436046 501842 436102
rect 501898 436046 501968 436102
rect 501648 435978 501968 436046
rect 501648 435922 501718 435978
rect 501774 435922 501842 435978
rect 501898 435922 501968 435978
rect 501648 435888 501968 435922
rect 532368 436350 532688 436384
rect 532368 436294 532438 436350
rect 532494 436294 532562 436350
rect 532618 436294 532688 436350
rect 532368 436226 532688 436294
rect 532368 436170 532438 436226
rect 532494 436170 532562 436226
rect 532618 436170 532688 436226
rect 532368 436102 532688 436170
rect 532368 436046 532438 436102
rect 532494 436046 532562 436102
rect 532618 436046 532688 436102
rect 532368 435978 532688 436046
rect 532368 435922 532438 435978
rect 532494 435922 532562 435978
rect 532618 435922 532688 435978
rect 532368 435888 532688 435922
rect 209808 424350 210128 424384
rect 209808 424294 209878 424350
rect 209934 424294 210002 424350
rect 210058 424294 210128 424350
rect 209808 424226 210128 424294
rect 209808 424170 209878 424226
rect 209934 424170 210002 424226
rect 210058 424170 210128 424226
rect 209808 424102 210128 424170
rect 209808 424046 209878 424102
rect 209934 424046 210002 424102
rect 210058 424046 210128 424102
rect 209808 423978 210128 424046
rect 209808 423922 209878 423978
rect 209934 423922 210002 423978
rect 210058 423922 210128 423978
rect 209808 423888 210128 423922
rect 240528 424350 240848 424384
rect 240528 424294 240598 424350
rect 240654 424294 240722 424350
rect 240778 424294 240848 424350
rect 240528 424226 240848 424294
rect 240528 424170 240598 424226
rect 240654 424170 240722 424226
rect 240778 424170 240848 424226
rect 240528 424102 240848 424170
rect 240528 424046 240598 424102
rect 240654 424046 240722 424102
rect 240778 424046 240848 424102
rect 240528 423978 240848 424046
rect 240528 423922 240598 423978
rect 240654 423922 240722 423978
rect 240778 423922 240848 423978
rect 240528 423888 240848 423922
rect 271248 424350 271568 424384
rect 271248 424294 271318 424350
rect 271374 424294 271442 424350
rect 271498 424294 271568 424350
rect 271248 424226 271568 424294
rect 271248 424170 271318 424226
rect 271374 424170 271442 424226
rect 271498 424170 271568 424226
rect 271248 424102 271568 424170
rect 271248 424046 271318 424102
rect 271374 424046 271442 424102
rect 271498 424046 271568 424102
rect 271248 423978 271568 424046
rect 271248 423922 271318 423978
rect 271374 423922 271442 423978
rect 271498 423922 271568 423978
rect 271248 423888 271568 423922
rect 301968 424350 302288 424384
rect 301968 424294 302038 424350
rect 302094 424294 302162 424350
rect 302218 424294 302288 424350
rect 301968 424226 302288 424294
rect 301968 424170 302038 424226
rect 302094 424170 302162 424226
rect 302218 424170 302288 424226
rect 301968 424102 302288 424170
rect 301968 424046 302038 424102
rect 302094 424046 302162 424102
rect 302218 424046 302288 424102
rect 301968 423978 302288 424046
rect 301968 423922 302038 423978
rect 302094 423922 302162 423978
rect 302218 423922 302288 423978
rect 301968 423888 302288 423922
rect 332688 424350 333008 424384
rect 332688 424294 332758 424350
rect 332814 424294 332882 424350
rect 332938 424294 333008 424350
rect 332688 424226 333008 424294
rect 332688 424170 332758 424226
rect 332814 424170 332882 424226
rect 332938 424170 333008 424226
rect 332688 424102 333008 424170
rect 332688 424046 332758 424102
rect 332814 424046 332882 424102
rect 332938 424046 333008 424102
rect 332688 423978 333008 424046
rect 332688 423922 332758 423978
rect 332814 423922 332882 423978
rect 332938 423922 333008 423978
rect 332688 423888 333008 423922
rect 363408 424350 363728 424384
rect 363408 424294 363478 424350
rect 363534 424294 363602 424350
rect 363658 424294 363728 424350
rect 363408 424226 363728 424294
rect 363408 424170 363478 424226
rect 363534 424170 363602 424226
rect 363658 424170 363728 424226
rect 363408 424102 363728 424170
rect 363408 424046 363478 424102
rect 363534 424046 363602 424102
rect 363658 424046 363728 424102
rect 363408 423978 363728 424046
rect 363408 423922 363478 423978
rect 363534 423922 363602 423978
rect 363658 423922 363728 423978
rect 363408 423888 363728 423922
rect 394128 424350 394448 424384
rect 394128 424294 394198 424350
rect 394254 424294 394322 424350
rect 394378 424294 394448 424350
rect 394128 424226 394448 424294
rect 394128 424170 394198 424226
rect 394254 424170 394322 424226
rect 394378 424170 394448 424226
rect 394128 424102 394448 424170
rect 394128 424046 394198 424102
rect 394254 424046 394322 424102
rect 394378 424046 394448 424102
rect 394128 423978 394448 424046
rect 394128 423922 394198 423978
rect 394254 423922 394322 423978
rect 394378 423922 394448 423978
rect 394128 423888 394448 423922
rect 424848 424350 425168 424384
rect 424848 424294 424918 424350
rect 424974 424294 425042 424350
rect 425098 424294 425168 424350
rect 424848 424226 425168 424294
rect 424848 424170 424918 424226
rect 424974 424170 425042 424226
rect 425098 424170 425168 424226
rect 424848 424102 425168 424170
rect 424848 424046 424918 424102
rect 424974 424046 425042 424102
rect 425098 424046 425168 424102
rect 424848 423978 425168 424046
rect 424848 423922 424918 423978
rect 424974 423922 425042 423978
rect 425098 423922 425168 423978
rect 424848 423888 425168 423922
rect 455568 424350 455888 424384
rect 455568 424294 455638 424350
rect 455694 424294 455762 424350
rect 455818 424294 455888 424350
rect 455568 424226 455888 424294
rect 455568 424170 455638 424226
rect 455694 424170 455762 424226
rect 455818 424170 455888 424226
rect 455568 424102 455888 424170
rect 455568 424046 455638 424102
rect 455694 424046 455762 424102
rect 455818 424046 455888 424102
rect 455568 423978 455888 424046
rect 455568 423922 455638 423978
rect 455694 423922 455762 423978
rect 455818 423922 455888 423978
rect 455568 423888 455888 423922
rect 486288 424350 486608 424384
rect 486288 424294 486358 424350
rect 486414 424294 486482 424350
rect 486538 424294 486608 424350
rect 486288 424226 486608 424294
rect 486288 424170 486358 424226
rect 486414 424170 486482 424226
rect 486538 424170 486608 424226
rect 486288 424102 486608 424170
rect 486288 424046 486358 424102
rect 486414 424046 486482 424102
rect 486538 424046 486608 424102
rect 486288 423978 486608 424046
rect 486288 423922 486358 423978
rect 486414 423922 486482 423978
rect 486538 423922 486608 423978
rect 486288 423888 486608 423922
rect 517008 424350 517328 424384
rect 517008 424294 517078 424350
rect 517134 424294 517202 424350
rect 517258 424294 517328 424350
rect 517008 424226 517328 424294
rect 517008 424170 517078 424226
rect 517134 424170 517202 424226
rect 517258 424170 517328 424226
rect 517008 424102 517328 424170
rect 517008 424046 517078 424102
rect 517134 424046 517202 424102
rect 517258 424046 517328 424102
rect 517008 423978 517328 424046
rect 517008 423922 517078 423978
rect 517134 423922 517202 423978
rect 517258 423922 517328 423978
rect 517008 423888 517328 423922
rect 194448 418350 194768 418384
rect 194448 418294 194518 418350
rect 194574 418294 194642 418350
rect 194698 418294 194768 418350
rect 194448 418226 194768 418294
rect 194448 418170 194518 418226
rect 194574 418170 194642 418226
rect 194698 418170 194768 418226
rect 194448 418102 194768 418170
rect 194448 418046 194518 418102
rect 194574 418046 194642 418102
rect 194698 418046 194768 418102
rect 194448 417978 194768 418046
rect 194448 417922 194518 417978
rect 194574 417922 194642 417978
rect 194698 417922 194768 417978
rect 194448 417888 194768 417922
rect 225168 418350 225488 418384
rect 225168 418294 225238 418350
rect 225294 418294 225362 418350
rect 225418 418294 225488 418350
rect 225168 418226 225488 418294
rect 225168 418170 225238 418226
rect 225294 418170 225362 418226
rect 225418 418170 225488 418226
rect 225168 418102 225488 418170
rect 225168 418046 225238 418102
rect 225294 418046 225362 418102
rect 225418 418046 225488 418102
rect 225168 417978 225488 418046
rect 225168 417922 225238 417978
rect 225294 417922 225362 417978
rect 225418 417922 225488 417978
rect 225168 417888 225488 417922
rect 255888 418350 256208 418384
rect 255888 418294 255958 418350
rect 256014 418294 256082 418350
rect 256138 418294 256208 418350
rect 255888 418226 256208 418294
rect 255888 418170 255958 418226
rect 256014 418170 256082 418226
rect 256138 418170 256208 418226
rect 255888 418102 256208 418170
rect 255888 418046 255958 418102
rect 256014 418046 256082 418102
rect 256138 418046 256208 418102
rect 255888 417978 256208 418046
rect 255888 417922 255958 417978
rect 256014 417922 256082 417978
rect 256138 417922 256208 417978
rect 255888 417888 256208 417922
rect 286608 418350 286928 418384
rect 286608 418294 286678 418350
rect 286734 418294 286802 418350
rect 286858 418294 286928 418350
rect 286608 418226 286928 418294
rect 286608 418170 286678 418226
rect 286734 418170 286802 418226
rect 286858 418170 286928 418226
rect 286608 418102 286928 418170
rect 286608 418046 286678 418102
rect 286734 418046 286802 418102
rect 286858 418046 286928 418102
rect 286608 417978 286928 418046
rect 286608 417922 286678 417978
rect 286734 417922 286802 417978
rect 286858 417922 286928 417978
rect 286608 417888 286928 417922
rect 317328 418350 317648 418384
rect 317328 418294 317398 418350
rect 317454 418294 317522 418350
rect 317578 418294 317648 418350
rect 317328 418226 317648 418294
rect 317328 418170 317398 418226
rect 317454 418170 317522 418226
rect 317578 418170 317648 418226
rect 317328 418102 317648 418170
rect 317328 418046 317398 418102
rect 317454 418046 317522 418102
rect 317578 418046 317648 418102
rect 317328 417978 317648 418046
rect 317328 417922 317398 417978
rect 317454 417922 317522 417978
rect 317578 417922 317648 417978
rect 317328 417888 317648 417922
rect 348048 418350 348368 418384
rect 348048 418294 348118 418350
rect 348174 418294 348242 418350
rect 348298 418294 348368 418350
rect 348048 418226 348368 418294
rect 348048 418170 348118 418226
rect 348174 418170 348242 418226
rect 348298 418170 348368 418226
rect 348048 418102 348368 418170
rect 348048 418046 348118 418102
rect 348174 418046 348242 418102
rect 348298 418046 348368 418102
rect 348048 417978 348368 418046
rect 348048 417922 348118 417978
rect 348174 417922 348242 417978
rect 348298 417922 348368 417978
rect 348048 417888 348368 417922
rect 378768 418350 379088 418384
rect 378768 418294 378838 418350
rect 378894 418294 378962 418350
rect 379018 418294 379088 418350
rect 378768 418226 379088 418294
rect 378768 418170 378838 418226
rect 378894 418170 378962 418226
rect 379018 418170 379088 418226
rect 378768 418102 379088 418170
rect 378768 418046 378838 418102
rect 378894 418046 378962 418102
rect 379018 418046 379088 418102
rect 378768 417978 379088 418046
rect 378768 417922 378838 417978
rect 378894 417922 378962 417978
rect 379018 417922 379088 417978
rect 378768 417888 379088 417922
rect 409488 418350 409808 418384
rect 409488 418294 409558 418350
rect 409614 418294 409682 418350
rect 409738 418294 409808 418350
rect 409488 418226 409808 418294
rect 409488 418170 409558 418226
rect 409614 418170 409682 418226
rect 409738 418170 409808 418226
rect 409488 418102 409808 418170
rect 409488 418046 409558 418102
rect 409614 418046 409682 418102
rect 409738 418046 409808 418102
rect 409488 417978 409808 418046
rect 409488 417922 409558 417978
rect 409614 417922 409682 417978
rect 409738 417922 409808 417978
rect 409488 417888 409808 417922
rect 440208 418350 440528 418384
rect 440208 418294 440278 418350
rect 440334 418294 440402 418350
rect 440458 418294 440528 418350
rect 440208 418226 440528 418294
rect 440208 418170 440278 418226
rect 440334 418170 440402 418226
rect 440458 418170 440528 418226
rect 440208 418102 440528 418170
rect 440208 418046 440278 418102
rect 440334 418046 440402 418102
rect 440458 418046 440528 418102
rect 440208 417978 440528 418046
rect 440208 417922 440278 417978
rect 440334 417922 440402 417978
rect 440458 417922 440528 417978
rect 440208 417888 440528 417922
rect 470928 418350 471248 418384
rect 470928 418294 470998 418350
rect 471054 418294 471122 418350
rect 471178 418294 471248 418350
rect 470928 418226 471248 418294
rect 470928 418170 470998 418226
rect 471054 418170 471122 418226
rect 471178 418170 471248 418226
rect 470928 418102 471248 418170
rect 470928 418046 470998 418102
rect 471054 418046 471122 418102
rect 471178 418046 471248 418102
rect 470928 417978 471248 418046
rect 470928 417922 470998 417978
rect 471054 417922 471122 417978
rect 471178 417922 471248 417978
rect 470928 417888 471248 417922
rect 501648 418350 501968 418384
rect 501648 418294 501718 418350
rect 501774 418294 501842 418350
rect 501898 418294 501968 418350
rect 501648 418226 501968 418294
rect 501648 418170 501718 418226
rect 501774 418170 501842 418226
rect 501898 418170 501968 418226
rect 501648 418102 501968 418170
rect 501648 418046 501718 418102
rect 501774 418046 501842 418102
rect 501898 418046 501968 418102
rect 501648 417978 501968 418046
rect 501648 417922 501718 417978
rect 501774 417922 501842 417978
rect 501898 417922 501968 417978
rect 501648 417888 501968 417922
rect 532368 418350 532688 418384
rect 532368 418294 532438 418350
rect 532494 418294 532562 418350
rect 532618 418294 532688 418350
rect 532368 418226 532688 418294
rect 532368 418170 532438 418226
rect 532494 418170 532562 418226
rect 532618 418170 532688 418226
rect 532368 418102 532688 418170
rect 532368 418046 532438 418102
rect 532494 418046 532562 418102
rect 532618 418046 532688 418102
rect 532368 417978 532688 418046
rect 532368 417922 532438 417978
rect 532494 417922 532562 417978
rect 532618 417922 532688 417978
rect 532368 417888 532688 417922
rect 308028 409332 308084 409342
rect 308028 409258 308084 409276
rect 308028 409192 308084 409202
rect 302652 409078 302708 409088
rect 302652 408884 302708 409022
rect 302652 408818 302708 408828
rect 376348 408996 376404 409006
rect 193116 282258 193172 282268
rect 193458 406350 194078 408578
rect 193458 406294 193554 406350
rect 193610 406294 193678 406350
rect 193734 406294 193802 406350
rect 193858 406294 193926 406350
rect 193982 406294 194078 406350
rect 193458 406226 194078 406294
rect 193458 406170 193554 406226
rect 193610 406170 193678 406226
rect 193734 406170 193802 406226
rect 193858 406170 193926 406226
rect 193982 406170 194078 406226
rect 193458 406102 194078 406170
rect 193458 406046 193554 406102
rect 193610 406046 193678 406102
rect 193734 406046 193802 406102
rect 193858 406046 193926 406102
rect 193982 406046 194078 406102
rect 193458 405978 194078 406046
rect 193458 405922 193554 405978
rect 193610 405922 193678 405978
rect 193734 405922 193802 405978
rect 193858 405922 193926 405978
rect 193982 405922 194078 405978
rect 193458 388350 194078 405922
rect 220458 400350 221078 408578
rect 220458 400294 220554 400350
rect 220610 400294 220678 400350
rect 220734 400294 220802 400350
rect 220858 400294 220926 400350
rect 220982 400294 221078 400350
rect 220458 400226 221078 400294
rect 220458 400170 220554 400226
rect 220610 400170 220678 400226
rect 220734 400170 220802 400226
rect 220858 400170 220926 400226
rect 220982 400170 221078 400226
rect 220458 400102 221078 400170
rect 220458 400046 220554 400102
rect 220610 400046 220678 400102
rect 220734 400046 220802 400102
rect 220858 400046 220926 400102
rect 220982 400046 221078 400102
rect 220458 399978 221078 400046
rect 220458 399922 220554 399978
rect 220610 399922 220678 399978
rect 220734 399922 220802 399978
rect 220858 399922 220926 399978
rect 220982 399922 221078 399978
rect 193458 388294 193554 388350
rect 193610 388294 193678 388350
rect 193734 388294 193802 388350
rect 193858 388294 193926 388350
rect 193982 388294 194078 388350
rect 193458 388226 194078 388294
rect 193458 388170 193554 388226
rect 193610 388170 193678 388226
rect 193734 388170 193802 388226
rect 193858 388170 193926 388226
rect 193982 388170 194078 388226
rect 193458 388102 194078 388170
rect 193458 388046 193554 388102
rect 193610 388046 193678 388102
rect 193734 388046 193802 388102
rect 193858 388046 193926 388102
rect 193982 388046 194078 388102
rect 193458 387978 194078 388046
rect 193458 387922 193554 387978
rect 193610 387922 193678 387978
rect 193734 387922 193802 387978
rect 193858 387922 193926 387978
rect 193982 387922 194078 387978
rect 193458 370350 194078 387922
rect 212492 388918 212548 388928
rect 209132 380548 209188 380558
rect 199724 377524 199780 377534
rect 199500 376404 199556 376414
rect 199276 375284 199332 375294
rect 199164 373044 199220 373054
rect 193458 370294 193554 370350
rect 193610 370294 193678 370350
rect 193734 370294 193802 370350
rect 193858 370294 193926 370350
rect 193982 370294 194078 370350
rect 193458 370226 194078 370294
rect 193458 370170 193554 370226
rect 193610 370170 193678 370226
rect 193734 370170 193802 370226
rect 193858 370170 193926 370226
rect 193982 370170 194078 370226
rect 193458 370102 194078 370170
rect 193458 370046 193554 370102
rect 193610 370046 193678 370102
rect 193734 370046 193802 370102
rect 193858 370046 193926 370102
rect 193982 370046 194078 370102
rect 193458 369978 194078 370046
rect 193458 369922 193554 369978
rect 193610 369922 193678 369978
rect 193734 369922 193802 369978
rect 193858 369922 193926 369978
rect 193982 369922 194078 369978
rect 193458 352350 194078 369922
rect 193458 352294 193554 352350
rect 193610 352294 193678 352350
rect 193734 352294 193802 352350
rect 193858 352294 193926 352350
rect 193982 352294 194078 352350
rect 193458 352226 194078 352294
rect 193458 352170 193554 352226
rect 193610 352170 193678 352226
rect 193734 352170 193802 352226
rect 193858 352170 193926 352226
rect 193982 352170 194078 352226
rect 193458 352102 194078 352170
rect 193458 352046 193554 352102
rect 193610 352046 193678 352102
rect 193734 352046 193802 352102
rect 193858 352046 193926 352102
rect 193982 352046 194078 352102
rect 193458 351978 194078 352046
rect 193458 351922 193554 351978
rect 193610 351922 193678 351978
rect 193734 351922 193802 351978
rect 193858 351922 193926 351978
rect 193982 351922 194078 351978
rect 193458 334350 194078 351922
rect 193458 334294 193554 334350
rect 193610 334294 193678 334350
rect 193734 334294 193802 334350
rect 193858 334294 193926 334350
rect 193982 334294 194078 334350
rect 193458 334226 194078 334294
rect 193458 334170 193554 334226
rect 193610 334170 193678 334226
rect 193734 334170 193802 334226
rect 193858 334170 193926 334226
rect 193982 334170 194078 334226
rect 193458 334102 194078 334170
rect 193458 334046 193554 334102
rect 193610 334046 193678 334102
rect 193734 334046 193802 334102
rect 193858 334046 193926 334102
rect 193982 334046 194078 334102
rect 193458 333978 194078 334046
rect 193458 333922 193554 333978
rect 193610 333922 193678 333978
rect 193734 333922 193802 333978
rect 193858 333922 193926 333978
rect 193982 333922 194078 333978
rect 193458 316350 194078 333922
rect 199052 371924 199108 371934
rect 199052 326116 199108 371868
rect 199164 349636 199220 372988
rect 199276 356356 199332 375228
rect 199276 356290 199332 356300
rect 199388 374164 199444 374174
rect 199388 352996 199444 374108
rect 199500 359716 199556 376348
rect 199724 363076 199780 377468
rect 199724 363010 199780 363020
rect 199500 359650 199556 359660
rect 199388 352930 199444 352940
rect 199164 349570 199220 349580
rect 199052 326050 199108 326060
rect 195244 322756 195300 322766
rect 195244 321972 195300 322700
rect 195244 321906 195300 321916
rect 193458 316294 193554 316350
rect 193610 316294 193678 316350
rect 193734 316294 193802 316350
rect 193858 316294 193926 316350
rect 193982 316294 194078 316350
rect 193458 316226 194078 316294
rect 193458 316170 193554 316226
rect 193610 316170 193678 316226
rect 193734 316170 193802 316226
rect 193858 316170 193926 316226
rect 193982 316170 194078 316226
rect 193458 316102 194078 316170
rect 193458 316046 193554 316102
rect 193610 316046 193678 316102
rect 193734 316046 193802 316102
rect 193858 316046 193926 316102
rect 193982 316046 194078 316102
rect 193458 315978 194078 316046
rect 193458 315922 193554 315978
rect 193610 315922 193678 315978
rect 193734 315922 193802 315978
rect 193858 315922 193926 315978
rect 193982 315922 194078 315978
rect 193458 298350 194078 315922
rect 193458 298294 193554 298350
rect 193610 298294 193678 298350
rect 193734 298294 193802 298350
rect 193858 298294 193926 298350
rect 193982 298294 194078 298350
rect 193458 298226 194078 298294
rect 193458 298170 193554 298226
rect 193610 298170 193678 298226
rect 193734 298170 193802 298226
rect 193858 298170 193926 298226
rect 193982 298170 194078 298226
rect 193458 298102 194078 298170
rect 193458 298046 193554 298102
rect 193610 298046 193678 298102
rect 193734 298046 193802 298102
rect 193858 298046 193926 298102
rect 193982 298046 194078 298102
rect 193458 297978 194078 298046
rect 193458 297922 193554 297978
rect 193610 297922 193678 297978
rect 193734 297922 193802 297978
rect 193858 297922 193926 297978
rect 193982 297922 194078 297978
rect 189738 274294 189834 274350
rect 189890 274294 189958 274350
rect 190014 274294 190082 274350
rect 190138 274294 190206 274350
rect 190262 274294 190358 274350
rect 189738 274226 190358 274294
rect 189738 274170 189834 274226
rect 189890 274170 189958 274226
rect 190014 274170 190082 274226
rect 190138 274170 190206 274226
rect 190262 274170 190358 274226
rect 189738 274102 190358 274170
rect 189738 274046 189834 274102
rect 189890 274046 189958 274102
rect 190014 274046 190082 274102
rect 190138 274046 190206 274102
rect 190262 274046 190358 274102
rect 189738 273978 190358 274046
rect 189084 273924 189140 273934
rect 189084 251972 189140 273868
rect 189738 273922 189834 273978
rect 189890 273922 189958 273978
rect 190014 273922 190082 273978
rect 190138 273922 190206 273978
rect 190262 273922 190358 273978
rect 189532 269892 189588 269902
rect 189532 268858 189588 269836
rect 189532 268792 189588 268802
rect 189196 261828 189252 261838
rect 189196 255108 189252 261772
rect 189196 255042 189252 255052
rect 189738 256350 190358 273922
rect 189738 256294 189834 256350
rect 189890 256294 189958 256350
rect 190014 256294 190082 256350
rect 190138 256294 190206 256350
rect 190262 256294 190358 256350
rect 189738 256226 190358 256294
rect 189738 256170 189834 256226
rect 189890 256170 189958 256226
rect 190014 256170 190082 256226
rect 190138 256170 190206 256226
rect 190262 256170 190358 256226
rect 189738 256102 190358 256170
rect 189738 256046 189834 256102
rect 189890 256046 189958 256102
rect 190014 256046 190082 256102
rect 190138 256046 190206 256102
rect 190262 256046 190358 256102
rect 189738 255978 190358 256046
rect 189738 255922 189834 255978
rect 189890 255922 189958 255978
rect 190014 255922 190082 255978
rect 190138 255922 190206 255978
rect 190262 255922 190358 255978
rect 189084 251906 189140 251916
rect 188972 246754 189028 246764
rect 162738 244294 162834 244350
rect 162890 244294 162958 244350
rect 163014 244294 163082 244350
rect 163138 244294 163206 244350
rect 163262 244294 163358 244350
rect 162738 244226 163358 244294
rect 162738 244170 162834 244226
rect 162890 244170 162958 244226
rect 163014 244170 163082 244226
rect 163138 244170 163206 244226
rect 163262 244170 163358 244226
rect 162738 244102 163358 244170
rect 162738 244046 162834 244102
rect 162890 244046 162958 244102
rect 163014 244046 163082 244102
rect 163138 244046 163206 244102
rect 163262 244046 163358 244102
rect 162738 243978 163358 244046
rect 162738 243922 162834 243978
rect 162890 243922 162958 243978
rect 163014 243922 163082 243978
rect 163138 243922 163206 243978
rect 163262 243922 163358 243978
rect 162738 226350 163358 243922
rect 162738 226294 162834 226350
rect 162890 226294 162958 226350
rect 163014 226294 163082 226350
rect 163138 226294 163206 226350
rect 163262 226294 163358 226350
rect 162738 226226 163358 226294
rect 162738 226170 162834 226226
rect 162890 226170 162958 226226
rect 163014 226170 163082 226226
rect 163138 226170 163206 226226
rect 163262 226170 163358 226226
rect 162738 226102 163358 226170
rect 162738 226046 162834 226102
rect 162890 226046 162958 226102
rect 163014 226046 163082 226102
rect 163138 226046 163206 226102
rect 163262 226046 163358 226102
rect 162738 225978 163358 226046
rect 162738 225922 162834 225978
rect 162890 225922 162958 225978
rect 163014 225922 163082 225978
rect 163138 225922 163206 225978
rect 163262 225922 163358 225978
rect 162738 210462 163358 225922
rect 189738 238350 190358 255922
rect 189738 238294 189834 238350
rect 189890 238294 189958 238350
rect 190014 238294 190082 238350
rect 190138 238294 190206 238350
rect 190262 238294 190358 238350
rect 189738 238226 190358 238294
rect 189738 238170 189834 238226
rect 189890 238170 189958 238226
rect 190014 238170 190082 238226
rect 190138 238170 190206 238226
rect 190262 238170 190358 238226
rect 189738 238102 190358 238170
rect 189738 238046 189834 238102
rect 189890 238046 189958 238102
rect 190014 238046 190082 238102
rect 190138 238046 190206 238102
rect 190262 238046 190358 238102
rect 189738 237978 190358 238046
rect 189738 237922 189834 237978
rect 189890 237922 189958 237978
rect 190014 237922 190082 237978
rect 190138 237922 190206 237978
rect 190262 237922 190358 237978
rect 189738 220350 190358 237922
rect 189738 220294 189834 220350
rect 189890 220294 189958 220350
rect 190014 220294 190082 220350
rect 190138 220294 190206 220350
rect 190262 220294 190358 220350
rect 189738 220226 190358 220294
rect 189738 220170 189834 220226
rect 189890 220170 189958 220226
rect 190014 220170 190082 220226
rect 190138 220170 190206 220226
rect 190262 220170 190358 220226
rect 189738 220102 190358 220170
rect 189738 220046 189834 220102
rect 189890 220046 189958 220102
rect 190014 220046 190082 220102
rect 190138 220046 190206 220102
rect 190262 220046 190358 220102
rect 189738 219978 190358 220046
rect 189738 219922 189834 219978
rect 189890 219922 189958 219978
rect 190014 219922 190082 219978
rect 190138 219922 190206 219978
rect 190262 219922 190358 219978
rect 189738 210462 190358 219922
rect 193458 280350 194078 297922
rect 209132 295764 209188 380492
rect 209132 295698 209188 295708
rect 193458 280294 193554 280350
rect 193610 280294 193678 280350
rect 193734 280294 193802 280350
rect 193858 280294 193926 280350
rect 193982 280294 194078 280350
rect 193458 280226 194078 280294
rect 193458 280170 193554 280226
rect 193610 280170 193678 280226
rect 193734 280170 193802 280226
rect 193858 280170 193926 280226
rect 193982 280170 194078 280226
rect 193458 280102 194078 280170
rect 193458 280046 193554 280102
rect 193610 280046 193678 280102
rect 193734 280046 193802 280102
rect 193858 280046 193926 280102
rect 193982 280046 194078 280102
rect 193458 279978 194078 280046
rect 193458 279922 193554 279978
rect 193610 279922 193678 279978
rect 193734 279922 193802 279978
rect 193858 279922 193926 279978
rect 193982 279922 194078 279978
rect 193458 262350 194078 279922
rect 193458 262294 193554 262350
rect 193610 262294 193678 262350
rect 193734 262294 193802 262350
rect 193858 262294 193926 262350
rect 193982 262294 194078 262350
rect 193458 262226 194078 262294
rect 193458 262170 193554 262226
rect 193610 262170 193678 262226
rect 193734 262170 193802 262226
rect 193858 262170 193926 262226
rect 193982 262170 194078 262226
rect 193458 262102 194078 262170
rect 193458 262046 193554 262102
rect 193610 262046 193678 262102
rect 193734 262046 193802 262102
rect 193858 262046 193926 262102
rect 193982 262046 194078 262102
rect 193458 261978 194078 262046
rect 193458 261922 193554 261978
rect 193610 261922 193678 261978
rect 193734 261922 193802 261978
rect 193858 261922 193926 261978
rect 193982 261922 194078 261978
rect 193458 244350 194078 261922
rect 193458 244294 193554 244350
rect 193610 244294 193678 244350
rect 193734 244294 193802 244350
rect 193858 244294 193926 244350
rect 193982 244294 194078 244350
rect 193458 244226 194078 244294
rect 193458 244170 193554 244226
rect 193610 244170 193678 244226
rect 193734 244170 193802 244226
rect 193858 244170 193926 244226
rect 193982 244170 194078 244226
rect 193458 244102 194078 244170
rect 193458 244046 193554 244102
rect 193610 244046 193678 244102
rect 193734 244046 193802 244102
rect 193858 244046 193926 244102
rect 193982 244046 194078 244102
rect 193458 243978 194078 244046
rect 193458 243922 193554 243978
rect 193610 243922 193678 243978
rect 193734 243922 193802 243978
rect 193858 243922 193926 243978
rect 193982 243922 194078 243978
rect 193458 226350 194078 243922
rect 212492 240548 212548 388862
rect 220458 382350 221078 399922
rect 220458 382294 220554 382350
rect 220610 382294 220678 382350
rect 220734 382294 220802 382350
rect 220858 382294 220926 382350
rect 220982 382294 221078 382350
rect 220458 382226 221078 382294
rect 220458 382170 220554 382226
rect 220610 382170 220678 382226
rect 220734 382170 220802 382226
rect 220858 382170 220926 382226
rect 220982 382170 221078 382226
rect 220458 382102 221078 382170
rect 220458 382046 220554 382102
rect 220610 382046 220678 382102
rect 220734 382046 220802 382102
rect 220858 382046 220926 382102
rect 220982 382046 221078 382102
rect 220458 381978 221078 382046
rect 220458 381922 220554 381978
rect 220610 381922 220678 381978
rect 220734 381922 220802 381978
rect 220858 381922 220926 381978
rect 220982 381922 221078 381978
rect 220458 364350 221078 381922
rect 220458 364294 220554 364350
rect 220610 364294 220678 364350
rect 220734 364294 220802 364350
rect 220858 364294 220926 364350
rect 220982 364294 221078 364350
rect 220458 364226 221078 364294
rect 220458 364170 220554 364226
rect 220610 364170 220678 364226
rect 220734 364170 220802 364226
rect 220858 364170 220926 364226
rect 220982 364170 221078 364226
rect 220458 364102 221078 364170
rect 220458 364046 220554 364102
rect 220610 364046 220678 364102
rect 220734 364046 220802 364102
rect 220858 364046 220926 364102
rect 220982 364046 221078 364102
rect 220458 363978 221078 364046
rect 220458 363922 220554 363978
rect 220610 363922 220678 363978
rect 220734 363922 220802 363978
rect 220858 363922 220926 363978
rect 220982 363922 221078 363978
rect 220458 346350 221078 363922
rect 220458 346294 220554 346350
rect 220610 346294 220678 346350
rect 220734 346294 220802 346350
rect 220858 346294 220926 346350
rect 220982 346294 221078 346350
rect 220458 346226 221078 346294
rect 220458 346170 220554 346226
rect 220610 346170 220678 346226
rect 220734 346170 220802 346226
rect 220858 346170 220926 346226
rect 220982 346170 221078 346226
rect 220458 346102 221078 346170
rect 220458 346046 220554 346102
rect 220610 346046 220678 346102
rect 220734 346046 220802 346102
rect 220858 346046 220926 346102
rect 220982 346046 221078 346102
rect 220458 345978 221078 346046
rect 220458 345922 220554 345978
rect 220610 345922 220678 345978
rect 220734 345922 220802 345978
rect 220858 345922 220926 345978
rect 220982 345922 221078 345978
rect 212492 240482 212548 240492
rect 219996 332724 220052 332734
rect 193458 226294 193554 226350
rect 193610 226294 193678 226350
rect 193734 226294 193802 226350
rect 193858 226294 193926 226350
rect 193982 226294 194078 226350
rect 193458 226226 194078 226294
rect 193458 226170 193554 226226
rect 193610 226170 193678 226226
rect 193734 226170 193802 226226
rect 193858 226170 193926 226226
rect 193982 226170 194078 226226
rect 193458 226102 194078 226170
rect 193458 226046 193554 226102
rect 193610 226046 193678 226102
rect 193734 226046 193802 226102
rect 193858 226046 193926 226102
rect 193982 226046 194078 226102
rect 193458 225978 194078 226046
rect 193458 225922 193554 225978
rect 193610 225922 193678 225978
rect 193734 225922 193802 225978
rect 193858 225922 193926 225978
rect 193982 225922 194078 225978
rect 193458 210462 194078 225922
rect 219996 214228 220052 332668
rect 219996 214162 220052 214172
rect 220458 328350 221078 345922
rect 224178 406350 224798 408578
rect 238140 407764 238196 407774
rect 238140 407458 238196 407708
rect 245196 407652 245252 407676
rect 245196 407572 245252 407582
rect 250348 407652 250404 407662
rect 238140 407392 238196 407402
rect 250348 406868 250404 407596
rect 224178 406294 224274 406350
rect 224330 406294 224398 406350
rect 224454 406294 224522 406350
rect 224578 406294 224646 406350
rect 224702 406294 224798 406350
rect 224178 406226 224798 406294
rect 224178 406170 224274 406226
rect 224330 406170 224398 406226
rect 224454 406170 224522 406226
rect 224578 406170 224646 406226
rect 224702 406170 224798 406226
rect 224178 406102 224798 406170
rect 224178 406046 224274 406102
rect 224330 406046 224398 406102
rect 224454 406046 224522 406102
rect 224578 406046 224646 406102
rect 224702 406046 224798 406102
rect 224178 405978 224798 406046
rect 224178 405922 224274 405978
rect 224330 405922 224398 405978
rect 224454 405922 224522 405978
rect 224578 405922 224646 405978
rect 224702 405922 224798 405978
rect 224178 388350 224798 405922
rect 230972 406532 231028 406542
rect 224178 388294 224274 388350
rect 224330 388294 224398 388350
rect 224454 388294 224522 388350
rect 224578 388294 224646 388350
rect 224702 388294 224798 388350
rect 224178 388226 224798 388294
rect 224178 388170 224274 388226
rect 224330 388170 224398 388226
rect 224454 388170 224522 388226
rect 224578 388170 224646 388226
rect 224702 388170 224798 388226
rect 224178 388102 224798 388170
rect 224178 388046 224274 388102
rect 224330 388046 224398 388102
rect 224454 388046 224522 388102
rect 224578 388046 224646 388102
rect 224702 388046 224798 388102
rect 224178 387978 224798 388046
rect 224178 387922 224274 387978
rect 224330 387922 224398 387978
rect 224454 387922 224522 387978
rect 224578 387922 224646 387978
rect 224702 387922 224798 387978
rect 224178 370350 224798 387922
rect 224178 370294 224274 370350
rect 224330 370294 224398 370350
rect 224454 370294 224522 370350
rect 224578 370294 224646 370350
rect 224702 370294 224798 370350
rect 224178 370226 224798 370294
rect 224178 370170 224274 370226
rect 224330 370170 224398 370226
rect 224454 370170 224522 370226
rect 224578 370170 224646 370226
rect 224702 370170 224798 370226
rect 224178 370102 224798 370170
rect 224178 370046 224274 370102
rect 224330 370046 224398 370102
rect 224454 370046 224522 370102
rect 224578 370046 224646 370102
rect 224702 370046 224798 370102
rect 224178 369978 224798 370046
rect 224178 369922 224274 369978
rect 224330 369922 224398 369978
rect 224454 369922 224522 369978
rect 224578 369922 224646 369978
rect 224702 369922 224798 369978
rect 224178 352350 224798 369922
rect 224178 352294 224274 352350
rect 224330 352294 224398 352350
rect 224454 352294 224522 352350
rect 224578 352294 224646 352350
rect 224702 352294 224798 352350
rect 224178 352226 224798 352294
rect 224178 352170 224274 352226
rect 224330 352170 224398 352226
rect 224454 352170 224522 352226
rect 224578 352170 224646 352226
rect 224702 352170 224798 352226
rect 224178 352102 224798 352170
rect 224178 352046 224274 352102
rect 224330 352046 224398 352102
rect 224454 352046 224522 352102
rect 224578 352046 224646 352102
rect 224702 352046 224798 352102
rect 224178 351978 224798 352046
rect 224178 351922 224274 351978
rect 224330 351922 224398 351978
rect 224454 351922 224522 351978
rect 224578 351922 224646 351978
rect 224702 351922 224798 351978
rect 224178 334350 224798 351922
rect 224178 334294 224274 334350
rect 224330 334294 224398 334350
rect 224454 334294 224522 334350
rect 224578 334294 224646 334350
rect 224702 334294 224798 334350
rect 224178 334226 224798 334294
rect 224178 334170 224274 334226
rect 224330 334170 224398 334226
rect 224454 334170 224522 334226
rect 224578 334170 224646 334226
rect 224702 334170 224798 334226
rect 224178 334102 224798 334170
rect 224178 334046 224274 334102
rect 224330 334046 224398 334102
rect 224454 334046 224522 334102
rect 224578 334046 224646 334102
rect 224702 334046 224798 334102
rect 224178 333978 224798 334046
rect 224178 333922 224274 333978
rect 224330 333922 224398 333978
rect 224454 333922 224522 333978
rect 224578 333922 224646 333978
rect 224702 333922 224798 333978
rect 220458 328294 220554 328350
rect 220610 328294 220678 328350
rect 220734 328294 220802 328350
rect 220858 328294 220926 328350
rect 220982 328294 221078 328350
rect 220458 328226 221078 328294
rect 220458 328170 220554 328226
rect 220610 328170 220678 328226
rect 220734 328170 220802 328226
rect 220858 328170 220926 328226
rect 220982 328170 221078 328226
rect 220458 328102 221078 328170
rect 220458 328046 220554 328102
rect 220610 328046 220678 328102
rect 220734 328046 220802 328102
rect 220858 328046 220926 328102
rect 220982 328046 221078 328102
rect 220458 327978 221078 328046
rect 220458 327922 220554 327978
rect 220610 327922 220678 327978
rect 220734 327922 220802 327978
rect 220858 327922 220926 327978
rect 220982 327922 221078 327978
rect 220458 310350 221078 327922
rect 220458 310294 220554 310350
rect 220610 310294 220678 310350
rect 220734 310294 220802 310350
rect 220858 310294 220926 310350
rect 220982 310294 221078 310350
rect 220458 310226 221078 310294
rect 220458 310170 220554 310226
rect 220610 310170 220678 310226
rect 220734 310170 220802 310226
rect 220858 310170 220926 310226
rect 220982 310170 221078 310226
rect 220458 310102 221078 310170
rect 220458 310046 220554 310102
rect 220610 310046 220678 310102
rect 220734 310046 220802 310102
rect 220858 310046 220926 310102
rect 220982 310046 221078 310102
rect 220458 309978 221078 310046
rect 220458 309922 220554 309978
rect 220610 309922 220678 309978
rect 220734 309922 220802 309978
rect 220858 309922 220926 309978
rect 220982 309922 221078 309978
rect 220458 292350 221078 309922
rect 220458 292294 220554 292350
rect 220610 292294 220678 292350
rect 220734 292294 220802 292350
rect 220858 292294 220926 292350
rect 220982 292294 221078 292350
rect 220458 292226 221078 292294
rect 220458 292170 220554 292226
rect 220610 292170 220678 292226
rect 220734 292170 220802 292226
rect 220858 292170 220926 292226
rect 220982 292170 221078 292226
rect 220458 292102 221078 292170
rect 220458 292046 220554 292102
rect 220610 292046 220678 292102
rect 220734 292046 220802 292102
rect 220858 292046 220926 292102
rect 220982 292046 221078 292102
rect 220458 291978 221078 292046
rect 220458 291922 220554 291978
rect 220610 291922 220678 291978
rect 220734 291922 220802 291978
rect 220858 291922 220926 291978
rect 220982 291922 221078 291978
rect 220458 274350 221078 291922
rect 220458 274294 220554 274350
rect 220610 274294 220678 274350
rect 220734 274294 220802 274350
rect 220858 274294 220926 274350
rect 220982 274294 221078 274350
rect 220458 274226 221078 274294
rect 220458 274170 220554 274226
rect 220610 274170 220678 274226
rect 220734 274170 220802 274226
rect 220858 274170 220926 274226
rect 220982 274170 221078 274226
rect 220458 274102 221078 274170
rect 220458 274046 220554 274102
rect 220610 274046 220678 274102
rect 220734 274046 220802 274102
rect 220858 274046 220926 274102
rect 220982 274046 221078 274102
rect 220458 273978 221078 274046
rect 220458 273922 220554 273978
rect 220610 273922 220678 273978
rect 220734 273922 220802 273978
rect 220858 273922 220926 273978
rect 220982 273922 221078 273978
rect 220458 256350 221078 273922
rect 220458 256294 220554 256350
rect 220610 256294 220678 256350
rect 220734 256294 220802 256350
rect 220858 256294 220926 256350
rect 220982 256294 221078 256350
rect 220458 256226 221078 256294
rect 220458 256170 220554 256226
rect 220610 256170 220678 256226
rect 220734 256170 220802 256226
rect 220858 256170 220926 256226
rect 220982 256170 221078 256226
rect 220458 256102 221078 256170
rect 220458 256046 220554 256102
rect 220610 256046 220678 256102
rect 220734 256046 220802 256102
rect 220858 256046 220926 256102
rect 220982 256046 221078 256102
rect 220458 255978 221078 256046
rect 220458 255922 220554 255978
rect 220610 255922 220678 255978
rect 220734 255922 220802 255978
rect 220858 255922 220926 255978
rect 220982 255922 221078 255978
rect 220458 238350 221078 255922
rect 220458 238294 220554 238350
rect 220610 238294 220678 238350
rect 220734 238294 220802 238350
rect 220858 238294 220926 238350
rect 220982 238294 221078 238350
rect 220458 238226 221078 238294
rect 220458 238170 220554 238226
rect 220610 238170 220678 238226
rect 220734 238170 220802 238226
rect 220858 238170 220926 238226
rect 220982 238170 221078 238226
rect 220458 238102 221078 238170
rect 220458 238046 220554 238102
rect 220610 238046 220678 238102
rect 220734 238046 220802 238102
rect 220858 238046 220926 238102
rect 220982 238046 221078 238102
rect 220458 237978 221078 238046
rect 220458 237922 220554 237978
rect 220610 237922 220678 237978
rect 220734 237922 220802 237978
rect 220858 237922 220926 237978
rect 220982 237922 221078 237978
rect 220458 220350 221078 237922
rect 223356 333844 223412 333854
rect 223356 236740 223412 333788
rect 223356 236674 223412 236684
rect 224178 316350 224798 333922
rect 230076 397348 230132 397358
rect 226716 328244 226772 328254
rect 224178 316294 224274 316350
rect 224330 316294 224398 316350
rect 224454 316294 224522 316350
rect 224578 316294 224646 316350
rect 224702 316294 224798 316350
rect 224178 316226 224798 316294
rect 224178 316170 224274 316226
rect 224330 316170 224398 316226
rect 224454 316170 224522 316226
rect 224578 316170 224646 316226
rect 224702 316170 224798 316226
rect 224178 316102 224798 316170
rect 224178 316046 224274 316102
rect 224330 316046 224398 316102
rect 224454 316046 224522 316102
rect 224578 316046 224646 316102
rect 224702 316046 224798 316102
rect 224178 315978 224798 316046
rect 224178 315922 224274 315978
rect 224330 315922 224398 315978
rect 224454 315922 224522 315978
rect 224578 315922 224646 315978
rect 224702 315922 224798 315978
rect 224178 298350 224798 315922
rect 224178 298294 224274 298350
rect 224330 298294 224398 298350
rect 224454 298294 224522 298350
rect 224578 298294 224646 298350
rect 224702 298294 224798 298350
rect 224178 298226 224798 298294
rect 224178 298170 224274 298226
rect 224330 298170 224398 298226
rect 224454 298170 224522 298226
rect 224578 298170 224646 298226
rect 224702 298170 224798 298226
rect 224178 298102 224798 298170
rect 224178 298046 224274 298102
rect 224330 298046 224398 298102
rect 224454 298046 224522 298102
rect 224578 298046 224646 298102
rect 224702 298046 224798 298102
rect 224178 297978 224798 298046
rect 224178 297922 224274 297978
rect 224330 297922 224398 297978
rect 224454 297922 224522 297978
rect 224578 297922 224646 297978
rect 224702 297922 224798 297978
rect 224178 280350 224798 297922
rect 224178 280294 224274 280350
rect 224330 280294 224398 280350
rect 224454 280294 224522 280350
rect 224578 280294 224646 280350
rect 224702 280294 224798 280350
rect 224178 280226 224798 280294
rect 224178 280170 224274 280226
rect 224330 280170 224398 280226
rect 224454 280170 224522 280226
rect 224578 280170 224646 280226
rect 224702 280170 224798 280226
rect 224178 280102 224798 280170
rect 224178 280046 224274 280102
rect 224330 280046 224398 280102
rect 224454 280046 224522 280102
rect 224578 280046 224646 280102
rect 224702 280046 224798 280102
rect 224178 279978 224798 280046
rect 224178 279922 224274 279978
rect 224330 279922 224398 279978
rect 224454 279922 224522 279978
rect 224578 279922 224646 279978
rect 224702 279922 224798 279978
rect 224178 262350 224798 279922
rect 224178 262294 224274 262350
rect 224330 262294 224398 262350
rect 224454 262294 224522 262350
rect 224578 262294 224646 262350
rect 224702 262294 224798 262350
rect 224178 262226 224798 262294
rect 224178 262170 224274 262226
rect 224330 262170 224398 262226
rect 224454 262170 224522 262226
rect 224578 262170 224646 262226
rect 224702 262170 224798 262226
rect 224178 262102 224798 262170
rect 224178 262046 224274 262102
rect 224330 262046 224398 262102
rect 224454 262046 224522 262102
rect 224578 262046 224646 262102
rect 224702 262046 224798 262102
rect 224178 261978 224798 262046
rect 224178 261922 224274 261978
rect 224330 261922 224398 261978
rect 224454 261922 224522 261978
rect 224578 261922 224646 261978
rect 224702 261922 224798 261978
rect 224178 244350 224798 261922
rect 224178 244294 224274 244350
rect 224330 244294 224398 244350
rect 224454 244294 224522 244350
rect 224578 244294 224646 244350
rect 224702 244294 224798 244350
rect 224178 244226 224798 244294
rect 224178 244170 224274 244226
rect 224330 244170 224398 244226
rect 224454 244170 224522 244226
rect 224578 244170 224646 244226
rect 224702 244170 224798 244226
rect 224178 244102 224798 244170
rect 224178 244046 224274 244102
rect 224330 244046 224398 244102
rect 224454 244046 224522 244102
rect 224578 244046 224646 244102
rect 224702 244046 224798 244102
rect 224178 243978 224798 244046
rect 224178 243922 224274 243978
rect 224330 243922 224398 243978
rect 224454 243922 224522 243978
rect 224578 243922 224646 243978
rect 224702 243922 224798 243978
rect 220458 220294 220554 220350
rect 220610 220294 220678 220350
rect 220734 220294 220802 220350
rect 220858 220294 220926 220350
rect 220982 220294 221078 220350
rect 220458 220226 221078 220294
rect 220458 220170 220554 220226
rect 220610 220170 220678 220226
rect 220734 220170 220802 220226
rect 220858 220170 220926 220226
rect 220982 220170 221078 220226
rect 220458 220102 221078 220170
rect 220458 220046 220554 220102
rect 220610 220046 220678 220102
rect 220734 220046 220802 220102
rect 220858 220046 220926 220102
rect 220982 220046 221078 220102
rect 220458 219978 221078 220046
rect 220458 219922 220554 219978
rect 220610 219922 220678 219978
rect 220734 219922 220802 219978
rect 220858 219922 220926 219978
rect 220982 219922 221078 219978
rect 220458 210462 221078 219922
rect 224178 226350 224798 243922
rect 224178 226294 224274 226350
rect 224330 226294 224398 226350
rect 224454 226294 224522 226350
rect 224578 226294 224646 226350
rect 224702 226294 224798 226350
rect 224178 226226 224798 226294
rect 224178 226170 224274 226226
rect 224330 226170 224398 226226
rect 224454 226170 224522 226226
rect 224578 226170 224646 226226
rect 224702 226170 224798 226226
rect 224178 226102 224798 226170
rect 224178 226046 224274 226102
rect 224330 226046 224398 226102
rect 224454 226046 224522 226102
rect 224578 226046 224646 226102
rect 224702 226046 224798 226102
rect 224178 225978 224798 226046
rect 224178 225922 224274 225978
rect 224330 225922 224398 225978
rect 224454 225922 224522 225978
rect 224578 225922 224646 225978
rect 224702 225922 224798 225978
rect 224178 210462 224798 225922
rect 226604 323764 226660 323774
rect 226604 209412 226660 323708
rect 226716 211092 226772 328188
rect 229964 327124 230020 327134
rect 228396 326004 228452 326014
rect 228284 304948 228340 304958
rect 228284 298004 228340 304892
rect 228284 297938 228340 297948
rect 226716 211026 226772 211036
rect 228396 209524 228452 325948
rect 229852 321524 229908 321534
rect 229852 211204 229908 321468
rect 229852 211138 229908 211148
rect 229964 209636 230020 327068
rect 230076 277844 230132 397292
rect 230076 277778 230132 277788
rect 230972 249418 231028 406476
rect 231756 404038 231812 404048
rect 231532 402500 231588 402510
rect 231420 324884 231476 324894
rect 231308 322644 231364 322654
rect 231196 320404 231252 320414
rect 230972 249352 231028 249362
rect 231084 278068 231140 278078
rect 231084 246708 231140 278012
rect 231084 246642 231140 246652
rect 231196 211316 231252 320348
rect 231196 211250 231252 211260
rect 231308 209860 231364 322588
rect 231308 209794 231364 209804
rect 231420 209748 231476 324828
rect 231532 278964 231588 402444
rect 231532 278898 231588 278908
rect 231644 402388 231700 402398
rect 231644 275604 231700 402332
rect 231756 276724 231812 403982
rect 236012 400932 236068 400942
rect 234892 399028 234948 399038
rect 234780 387268 234836 387278
rect 234444 329364 234500 329374
rect 231756 276658 231812 276668
rect 232428 319284 232484 319294
rect 231644 275538 231700 275548
rect 231756 272244 231812 272254
rect 231532 271348 231588 271358
rect 231532 250292 231588 271292
rect 231756 255332 231812 272188
rect 231756 255266 231812 255276
rect 231532 250226 231588 250236
rect 231868 246932 231924 246942
rect 231868 246178 231924 246876
rect 231868 246112 231924 246122
rect 232428 212996 232484 319228
rect 233212 318164 233268 318174
rect 233100 315924 233156 315934
rect 232652 314804 232708 314814
rect 232540 313684 232596 313694
rect 232540 256228 232596 313628
rect 232540 256162 232596 256172
rect 232652 254660 232708 314748
rect 232876 312564 232932 312574
rect 232652 254594 232708 254604
rect 232764 311444 232820 311454
rect 232764 234388 232820 311388
rect 232764 234322 232820 234332
rect 232876 217812 232932 312508
rect 232876 217746 232932 217756
rect 232988 310324 233044 310334
rect 232988 213220 233044 310268
rect 233100 216580 233156 315868
rect 233100 216514 233156 216524
rect 233212 216356 233268 318108
rect 233212 216290 233268 216300
rect 233324 317044 233380 317054
rect 233324 214340 233380 316988
rect 233324 214274 233380 214284
rect 232988 213154 233044 213164
rect 232428 212930 232484 212940
rect 234444 209972 234500 329308
rect 234780 274484 234836 387212
rect 234892 280084 234948 398972
rect 235900 382618 235956 382628
rect 235900 339220 235956 382562
rect 235900 339154 235956 339164
rect 234892 280018 234948 280028
rect 235004 330484 235060 330494
rect 234780 274418 234836 274428
rect 234668 268884 234724 268894
rect 234556 266644 234612 266654
rect 234556 239428 234612 266588
rect 234668 241108 234724 268828
rect 234892 267764 234948 267774
rect 234668 241042 234724 241052
rect 234780 265524 234836 265534
rect 234556 239362 234612 239372
rect 234780 236516 234836 265468
rect 234780 236450 234836 236460
rect 234892 236404 234948 267708
rect 234892 236338 234948 236348
rect 235004 211428 235060 330428
rect 235788 273364 235844 273374
rect 235116 271124 235172 271134
rect 235116 255220 235172 271068
rect 235340 270004 235396 270014
rect 235340 255388 235396 269948
rect 235676 267988 235732 267998
rect 235676 264898 235732 267932
rect 235452 264842 235732 264898
rect 235452 255780 235508 264842
rect 235564 264628 235620 264638
rect 235564 256438 235620 264572
rect 235788 256564 235844 273308
rect 235788 256498 235844 256508
rect 235900 266308 235956 266318
rect 235564 256382 235844 256438
rect 235452 255714 235508 255724
rect 235340 255332 235620 255388
rect 235116 255154 235172 255164
rect 235564 239540 235620 255332
rect 235788 254772 235844 256382
rect 235900 256340 235956 266252
rect 235900 256274 235956 256284
rect 235788 254706 235844 254716
rect 236012 251748 236068 400876
rect 236236 392532 236292 392542
rect 236012 251682 236068 251692
rect 236124 385364 236180 385374
rect 235564 239474 235620 239484
rect 236124 236628 236180 385308
rect 236124 236562 236180 236572
rect 235004 211362 235060 211372
rect 236236 211078 236292 392476
rect 237916 392420 237972 392430
rect 237804 385924 237860 385934
rect 237692 385678 237748 385688
rect 237580 268858 237636 268868
rect 237580 257460 237636 268802
rect 237580 257394 237636 257404
rect 236236 211012 236292 211022
rect 237692 210980 237748 385622
rect 237804 211540 237860 385868
rect 237804 211474 237860 211484
rect 237692 210914 237748 210924
rect 237916 210898 237972 392364
rect 238252 389818 238308 389828
rect 238252 388164 238308 389762
rect 238252 388098 238308 388108
rect 250348 384580 250404 406812
rect 250348 384514 250404 384524
rect 254898 406350 255518 408578
rect 254898 406294 254994 406350
rect 255050 406294 255118 406350
rect 255174 406294 255242 406350
rect 255298 406294 255366 406350
rect 255422 406294 255518 406350
rect 254898 406226 255518 406294
rect 254898 406170 254994 406226
rect 255050 406170 255118 406226
rect 255174 406170 255242 406226
rect 255298 406170 255366 406226
rect 255422 406170 255518 406226
rect 254898 406102 255518 406170
rect 254898 406046 254994 406102
rect 255050 406046 255118 406102
rect 255174 406046 255242 406102
rect 255298 406046 255366 406102
rect 255422 406046 255518 406102
rect 254898 405978 255518 406046
rect 254898 405922 254994 405978
rect 255050 405922 255118 405978
rect 255174 405922 255242 405978
rect 255298 405922 255366 405978
rect 255422 405922 255518 405978
rect 254898 388350 255518 405922
rect 261212 407988 261268 407998
rect 261212 404852 261268 407932
rect 261212 404786 261268 404796
rect 285618 406350 286238 408578
rect 285618 406294 285714 406350
rect 285770 406294 285838 406350
rect 285894 406294 285962 406350
rect 286018 406294 286086 406350
rect 286142 406294 286238 406350
rect 285618 406226 286238 406294
rect 285618 406170 285714 406226
rect 285770 406170 285838 406226
rect 285894 406170 285962 406226
rect 286018 406170 286086 406226
rect 286142 406170 286238 406226
rect 285618 406102 286238 406170
rect 285618 406046 285714 406102
rect 285770 406046 285838 406102
rect 285894 406046 285962 406102
rect 286018 406046 286086 406102
rect 286142 406046 286238 406102
rect 285618 405978 286238 406046
rect 285618 405922 285714 405978
rect 285770 405922 285838 405978
rect 285894 405922 285962 405978
rect 286018 405922 286086 405978
rect 286142 405922 286238 405978
rect 254898 388294 254994 388350
rect 255050 388294 255118 388350
rect 255174 388294 255242 388350
rect 255298 388294 255366 388350
rect 255422 388294 255518 388350
rect 254898 388226 255518 388294
rect 254898 388170 254994 388226
rect 255050 388170 255118 388226
rect 255174 388170 255242 388226
rect 255298 388170 255366 388226
rect 255422 388170 255518 388226
rect 254898 388102 255518 388170
rect 254898 388046 254994 388102
rect 255050 388046 255118 388102
rect 255174 388046 255242 388102
rect 255298 388046 255366 388102
rect 255422 388046 255518 388102
rect 282156 388738 282212 388748
rect 282156 388164 282212 388682
rect 282156 388098 282212 388108
rect 285618 388350 286238 405922
rect 285618 388294 285714 388350
rect 285770 388294 285838 388350
rect 285894 388294 285962 388350
rect 286018 388294 286086 388350
rect 286142 388294 286238 388350
rect 285618 388226 286238 388294
rect 285618 388170 285714 388226
rect 285770 388170 285838 388226
rect 285894 388170 285962 388226
rect 286018 388170 286086 388226
rect 286142 388170 286238 388226
rect 285618 388102 286238 388170
rect 254898 387978 255518 388046
rect 254898 387922 254994 387978
rect 255050 387922 255118 387978
rect 255174 387922 255242 387978
rect 255298 387922 255366 387978
rect 255422 387922 255518 387978
rect 254898 383870 255518 387922
rect 285618 388046 285714 388102
rect 285770 388046 285838 388102
rect 285894 388046 285962 388102
rect 286018 388046 286086 388102
rect 286142 388046 286238 388102
rect 285618 387978 286238 388046
rect 285618 387922 285714 387978
rect 285770 387922 285838 387978
rect 285894 387922 285962 387978
rect 286018 387922 286086 387978
rect 286142 387922 286238 387978
rect 267820 385498 267876 385514
rect 267820 385410 267876 385420
rect 273196 385498 273252 385514
rect 273196 385410 273252 385420
rect 266028 385364 266084 385374
rect 266028 384244 266084 385308
rect 269612 385364 269668 385374
rect 269612 385252 269668 385262
rect 271404 385364 271460 385374
rect 271404 385252 271460 385262
rect 275884 385364 275940 385374
rect 275884 384468 275940 385308
rect 281260 385364 281316 385374
rect 281260 384580 281316 385308
rect 281260 384514 281316 384524
rect 283052 385364 283108 385374
rect 275884 384402 275940 384412
rect 283052 384468 283108 385308
rect 283052 384402 283108 384412
rect 266028 384178 266084 384188
rect 285618 383870 286238 387922
rect 286300 406980 286356 406990
rect 286300 385678 286356 406924
rect 303996 406980 304052 406990
rect 297388 388918 297444 388928
rect 297388 388164 297444 388862
rect 297388 388098 297444 388108
rect 286300 385612 286356 385622
rect 303996 385678 304052 406924
rect 303996 385612 304052 385622
rect 316338 406350 316958 408578
rect 316338 406294 316434 406350
rect 316490 406294 316558 406350
rect 316614 406294 316682 406350
rect 316738 406294 316806 406350
rect 316862 406294 316958 406350
rect 316338 406226 316958 406294
rect 316338 406170 316434 406226
rect 316490 406170 316558 406226
rect 316614 406170 316682 406226
rect 316738 406170 316806 406226
rect 316862 406170 316958 406226
rect 316338 406102 316958 406170
rect 316338 406046 316434 406102
rect 316490 406046 316558 406102
rect 316614 406046 316682 406102
rect 316738 406046 316806 406102
rect 316862 406046 316958 406102
rect 316338 405978 316958 406046
rect 316338 405922 316434 405978
rect 316490 405922 316558 405978
rect 316614 405922 316682 405978
rect 316738 405922 316806 405978
rect 316862 405922 316958 405978
rect 316338 388350 316958 405922
rect 316338 388294 316434 388350
rect 316490 388294 316558 388350
rect 316614 388294 316682 388350
rect 316738 388294 316806 388350
rect 316862 388294 316958 388350
rect 316338 388226 316958 388294
rect 316338 388170 316434 388226
rect 316490 388170 316558 388226
rect 316614 388170 316682 388226
rect 316738 388170 316806 388226
rect 316862 388170 316958 388226
rect 316338 388102 316958 388170
rect 316338 388046 316434 388102
rect 316490 388046 316558 388102
rect 316614 388046 316682 388102
rect 316738 388046 316806 388102
rect 316862 388046 316958 388102
rect 316338 387978 316958 388046
rect 316338 387922 316434 387978
rect 316490 387922 316558 387978
rect 316614 387922 316682 387978
rect 316738 387922 316806 387978
rect 316862 387922 316958 387978
rect 287532 385364 287588 385374
rect 287532 384418 287588 385308
rect 287532 384352 287588 384362
rect 288428 385364 288484 385374
rect 288428 384238 288484 385308
rect 288428 384172 288484 384182
rect 289324 385364 289380 385374
rect 289324 383878 289380 385308
rect 290220 385364 290276 385374
rect 290220 384058 290276 385308
rect 291116 385364 291172 385374
rect 291116 384244 291172 385308
rect 291116 384178 291172 384188
rect 292908 385364 292964 385374
rect 292908 384132 292964 385308
rect 292908 384066 292964 384076
rect 293804 385364 293860 385374
rect 290220 383992 290276 384002
rect 293804 384020 293860 385308
rect 293804 383954 293860 383964
rect 294700 385364 294756 385374
rect 294700 383908 294756 385308
rect 309036 385364 309092 385374
rect 309036 384356 309092 385308
rect 309036 384290 309092 384300
rect 316338 383870 316958 387922
rect 347058 406350 347678 408578
rect 347058 406294 347154 406350
rect 347210 406294 347278 406350
rect 347334 406294 347402 406350
rect 347458 406294 347526 406350
rect 347582 406294 347678 406350
rect 347058 406226 347678 406294
rect 347058 406170 347154 406226
rect 347210 406170 347278 406226
rect 347334 406170 347402 406226
rect 347458 406170 347526 406226
rect 347582 406170 347678 406226
rect 347058 406102 347678 406170
rect 347058 406046 347154 406102
rect 347210 406046 347278 406102
rect 347334 406046 347402 406102
rect 347458 406046 347526 406102
rect 347582 406046 347678 406102
rect 347058 405978 347678 406046
rect 347058 405922 347154 405978
rect 347210 405922 347278 405978
rect 347334 405922 347402 405978
rect 347458 405922 347526 405978
rect 347582 405922 347678 405978
rect 347058 388350 347678 405922
rect 375452 407652 375508 407662
rect 347058 388294 347154 388350
rect 347210 388294 347278 388350
rect 347334 388294 347402 388350
rect 347458 388294 347526 388350
rect 347582 388294 347678 388350
rect 347058 388226 347678 388294
rect 347058 388170 347154 388226
rect 347210 388170 347278 388226
rect 347334 388170 347402 388226
rect 347458 388170 347526 388226
rect 347582 388170 347678 388226
rect 347058 388102 347678 388170
rect 347058 388046 347154 388102
rect 347210 388046 347278 388102
rect 347334 388046 347402 388102
rect 347458 388046 347526 388102
rect 347582 388046 347678 388102
rect 347058 387978 347678 388046
rect 347058 387922 347154 387978
rect 347210 387922 347278 387978
rect 347334 387922 347402 387978
rect 347458 387922 347526 387978
rect 347582 387922 347678 387978
rect 347058 383870 347678 387922
rect 372988 393204 373044 393214
rect 372316 386148 372372 386158
rect 294700 383842 294756 383852
rect 289324 383812 289380 383822
rect 240448 382269 240768 382284
rect 240448 382213 240518 382269
rect 240574 382213 240642 382269
rect 240698 382213 240768 382269
rect 240448 382145 240768 382213
rect 240448 382089 240518 382145
rect 240574 382089 240642 382145
rect 240698 382089 240768 382145
rect 240448 382021 240768 382089
rect 240448 381965 240518 382021
rect 240574 381965 240642 382021
rect 240698 381965 240768 382021
rect 240448 381897 240768 381965
rect 240448 381841 240518 381897
rect 240574 381841 240642 381897
rect 240698 381841 240768 381897
rect 240448 381826 240768 381841
rect 271168 382269 271488 382284
rect 271168 382213 271238 382269
rect 271294 382213 271362 382269
rect 271418 382213 271488 382269
rect 271168 382145 271488 382213
rect 271168 382089 271238 382145
rect 271294 382089 271362 382145
rect 271418 382089 271488 382145
rect 271168 382021 271488 382089
rect 271168 381965 271238 382021
rect 271294 381965 271362 382021
rect 271418 381965 271488 382021
rect 271168 381897 271488 381965
rect 271168 381841 271238 381897
rect 271294 381841 271362 381897
rect 271418 381841 271488 381897
rect 271168 381826 271488 381841
rect 301888 382269 302208 382284
rect 301888 382213 301958 382269
rect 302014 382213 302082 382269
rect 302138 382213 302208 382269
rect 301888 382145 302208 382213
rect 301888 382089 301958 382145
rect 302014 382089 302082 382145
rect 302138 382089 302208 382145
rect 301888 382021 302208 382089
rect 301888 381965 301958 382021
rect 302014 381965 302082 382021
rect 302138 381965 302208 382021
rect 301888 381897 302208 381965
rect 301888 381841 301958 381897
rect 302014 381841 302082 381897
rect 302138 381841 302208 381897
rect 301888 381826 302208 381841
rect 332608 382269 332928 382284
rect 332608 382213 332678 382269
rect 332734 382213 332802 382269
rect 332858 382213 332928 382269
rect 332608 382145 332928 382213
rect 332608 382089 332678 382145
rect 332734 382089 332802 382145
rect 332858 382089 332928 382145
rect 332608 382021 332928 382089
rect 332608 381965 332678 382021
rect 332734 381965 332802 382021
rect 332858 381965 332928 382021
rect 332608 381897 332928 381965
rect 332608 381841 332678 381897
rect 332734 381841 332802 381897
rect 332858 381841 332928 381897
rect 332608 381826 332928 381841
rect 363328 382269 363648 382284
rect 363328 382213 363398 382269
rect 363454 382213 363522 382269
rect 363578 382213 363648 382269
rect 363328 382145 363648 382213
rect 363328 382089 363398 382145
rect 363454 382089 363522 382145
rect 363578 382089 363648 382145
rect 363328 382021 363648 382089
rect 363328 381965 363398 382021
rect 363454 381965 363522 382021
rect 363578 381965 363648 382021
rect 363328 381897 363648 381965
rect 363328 381841 363398 381897
rect 363454 381841 363522 381897
rect 363578 381841 363648 381897
rect 363328 381826 363648 381841
rect 255808 370350 256128 370384
rect 255808 370294 255878 370350
rect 255934 370294 256002 370350
rect 256058 370294 256128 370350
rect 255808 370226 256128 370294
rect 255808 370170 255878 370226
rect 255934 370170 256002 370226
rect 256058 370170 256128 370226
rect 255808 370102 256128 370170
rect 255808 370046 255878 370102
rect 255934 370046 256002 370102
rect 256058 370046 256128 370102
rect 255808 369978 256128 370046
rect 255808 369922 255878 369978
rect 255934 369922 256002 369978
rect 256058 369922 256128 369978
rect 255808 369888 256128 369922
rect 286528 370350 286848 370384
rect 286528 370294 286598 370350
rect 286654 370294 286722 370350
rect 286778 370294 286848 370350
rect 286528 370226 286848 370294
rect 286528 370170 286598 370226
rect 286654 370170 286722 370226
rect 286778 370170 286848 370226
rect 286528 370102 286848 370170
rect 286528 370046 286598 370102
rect 286654 370046 286722 370102
rect 286778 370046 286848 370102
rect 286528 369978 286848 370046
rect 286528 369922 286598 369978
rect 286654 369922 286722 369978
rect 286778 369922 286848 369978
rect 286528 369888 286848 369922
rect 317248 370350 317568 370384
rect 317248 370294 317318 370350
rect 317374 370294 317442 370350
rect 317498 370294 317568 370350
rect 317248 370226 317568 370294
rect 317248 370170 317318 370226
rect 317374 370170 317442 370226
rect 317498 370170 317568 370226
rect 317248 370102 317568 370170
rect 317248 370046 317318 370102
rect 317374 370046 317442 370102
rect 317498 370046 317568 370102
rect 317248 369978 317568 370046
rect 317248 369922 317318 369978
rect 317374 369922 317442 369978
rect 317498 369922 317568 369978
rect 317248 369888 317568 369922
rect 347968 370350 348288 370384
rect 347968 370294 348038 370350
rect 348094 370294 348162 370350
rect 348218 370294 348288 370350
rect 347968 370226 348288 370294
rect 347968 370170 348038 370226
rect 348094 370170 348162 370226
rect 348218 370170 348288 370226
rect 347968 370102 348288 370170
rect 347968 370046 348038 370102
rect 348094 370046 348162 370102
rect 348218 370046 348288 370102
rect 347968 369978 348288 370046
rect 347968 369922 348038 369978
rect 348094 369922 348162 369978
rect 348218 369922 348288 369978
rect 347968 369888 348288 369922
rect 240448 364350 240768 364384
rect 240448 364294 240518 364350
rect 240574 364294 240642 364350
rect 240698 364294 240768 364350
rect 240448 364226 240768 364294
rect 240448 364170 240518 364226
rect 240574 364170 240642 364226
rect 240698 364170 240768 364226
rect 240448 364102 240768 364170
rect 240448 364046 240518 364102
rect 240574 364046 240642 364102
rect 240698 364046 240768 364102
rect 240448 363978 240768 364046
rect 240448 363922 240518 363978
rect 240574 363922 240642 363978
rect 240698 363922 240768 363978
rect 240448 363888 240768 363922
rect 271168 364350 271488 364384
rect 271168 364294 271238 364350
rect 271294 364294 271362 364350
rect 271418 364294 271488 364350
rect 271168 364226 271488 364294
rect 271168 364170 271238 364226
rect 271294 364170 271362 364226
rect 271418 364170 271488 364226
rect 271168 364102 271488 364170
rect 271168 364046 271238 364102
rect 271294 364046 271362 364102
rect 271418 364046 271488 364102
rect 271168 363978 271488 364046
rect 271168 363922 271238 363978
rect 271294 363922 271362 363978
rect 271418 363922 271488 363978
rect 271168 363888 271488 363922
rect 301888 364350 302208 364384
rect 301888 364294 301958 364350
rect 302014 364294 302082 364350
rect 302138 364294 302208 364350
rect 301888 364226 302208 364294
rect 301888 364170 301958 364226
rect 302014 364170 302082 364226
rect 302138 364170 302208 364226
rect 301888 364102 302208 364170
rect 301888 364046 301958 364102
rect 302014 364046 302082 364102
rect 302138 364046 302208 364102
rect 301888 363978 302208 364046
rect 301888 363922 301958 363978
rect 302014 363922 302082 363978
rect 302138 363922 302208 363978
rect 301888 363888 302208 363922
rect 332608 364350 332928 364384
rect 332608 364294 332678 364350
rect 332734 364294 332802 364350
rect 332858 364294 332928 364350
rect 332608 364226 332928 364294
rect 332608 364170 332678 364226
rect 332734 364170 332802 364226
rect 332858 364170 332928 364226
rect 332608 364102 332928 364170
rect 332608 364046 332678 364102
rect 332734 364046 332802 364102
rect 332858 364046 332928 364102
rect 332608 363978 332928 364046
rect 332608 363922 332678 363978
rect 332734 363922 332802 363978
rect 332858 363922 332928 363978
rect 332608 363888 332928 363922
rect 363328 364350 363648 364384
rect 363328 364294 363398 364350
rect 363454 364294 363522 364350
rect 363578 364294 363648 364350
rect 363328 364226 363648 364294
rect 363328 364170 363398 364226
rect 363454 364170 363522 364226
rect 363578 364170 363648 364226
rect 363328 364102 363648 364170
rect 363328 364046 363398 364102
rect 363454 364046 363522 364102
rect 363578 364046 363648 364102
rect 363328 363978 363648 364046
rect 363328 363922 363398 363978
rect 363454 363922 363522 363978
rect 363578 363922 363648 363978
rect 363328 363888 363648 363922
rect 255808 352350 256128 352384
rect 255808 352294 255878 352350
rect 255934 352294 256002 352350
rect 256058 352294 256128 352350
rect 255808 352226 256128 352294
rect 255808 352170 255878 352226
rect 255934 352170 256002 352226
rect 256058 352170 256128 352226
rect 255808 352102 256128 352170
rect 255808 352046 255878 352102
rect 255934 352046 256002 352102
rect 256058 352046 256128 352102
rect 255808 351978 256128 352046
rect 255808 351922 255878 351978
rect 255934 351922 256002 351978
rect 256058 351922 256128 351978
rect 255808 351888 256128 351922
rect 286528 352350 286848 352384
rect 286528 352294 286598 352350
rect 286654 352294 286722 352350
rect 286778 352294 286848 352350
rect 286528 352226 286848 352294
rect 286528 352170 286598 352226
rect 286654 352170 286722 352226
rect 286778 352170 286848 352226
rect 286528 352102 286848 352170
rect 286528 352046 286598 352102
rect 286654 352046 286722 352102
rect 286778 352046 286848 352102
rect 286528 351978 286848 352046
rect 286528 351922 286598 351978
rect 286654 351922 286722 351978
rect 286778 351922 286848 351978
rect 286528 351888 286848 351922
rect 317248 352350 317568 352384
rect 317248 352294 317318 352350
rect 317374 352294 317442 352350
rect 317498 352294 317568 352350
rect 317248 352226 317568 352294
rect 317248 352170 317318 352226
rect 317374 352170 317442 352226
rect 317498 352170 317568 352226
rect 317248 352102 317568 352170
rect 317248 352046 317318 352102
rect 317374 352046 317442 352102
rect 317498 352046 317568 352102
rect 317248 351978 317568 352046
rect 317248 351922 317318 351978
rect 317374 351922 317442 351978
rect 317498 351922 317568 351978
rect 317248 351888 317568 351922
rect 347968 352350 348288 352384
rect 347968 352294 348038 352350
rect 348094 352294 348162 352350
rect 348218 352294 348288 352350
rect 347968 352226 348288 352294
rect 347968 352170 348038 352226
rect 348094 352170 348162 352226
rect 348218 352170 348288 352226
rect 347968 352102 348288 352170
rect 347968 352046 348038 352102
rect 348094 352046 348162 352102
rect 348218 352046 348288 352102
rect 347968 351978 348288 352046
rect 347968 351922 348038 351978
rect 348094 351922 348162 351978
rect 348218 351922 348288 351978
rect 347968 351888 348288 351922
rect 240448 346350 240768 346384
rect 240448 346294 240518 346350
rect 240574 346294 240642 346350
rect 240698 346294 240768 346350
rect 240448 346226 240768 346294
rect 240448 346170 240518 346226
rect 240574 346170 240642 346226
rect 240698 346170 240768 346226
rect 240448 346102 240768 346170
rect 240448 346046 240518 346102
rect 240574 346046 240642 346102
rect 240698 346046 240768 346102
rect 240448 345978 240768 346046
rect 240448 345922 240518 345978
rect 240574 345922 240642 345978
rect 240698 345922 240768 345978
rect 240448 345888 240768 345922
rect 271168 346350 271488 346384
rect 271168 346294 271238 346350
rect 271294 346294 271362 346350
rect 271418 346294 271488 346350
rect 271168 346226 271488 346294
rect 271168 346170 271238 346226
rect 271294 346170 271362 346226
rect 271418 346170 271488 346226
rect 271168 346102 271488 346170
rect 271168 346046 271238 346102
rect 271294 346046 271362 346102
rect 271418 346046 271488 346102
rect 271168 345978 271488 346046
rect 271168 345922 271238 345978
rect 271294 345922 271362 345978
rect 271418 345922 271488 345978
rect 271168 345888 271488 345922
rect 301888 346350 302208 346384
rect 301888 346294 301958 346350
rect 302014 346294 302082 346350
rect 302138 346294 302208 346350
rect 301888 346226 302208 346294
rect 301888 346170 301958 346226
rect 302014 346170 302082 346226
rect 302138 346170 302208 346226
rect 301888 346102 302208 346170
rect 301888 346046 301958 346102
rect 302014 346046 302082 346102
rect 302138 346046 302208 346102
rect 301888 345978 302208 346046
rect 301888 345922 301958 345978
rect 302014 345922 302082 345978
rect 302138 345922 302208 345978
rect 301888 345888 302208 345922
rect 332608 346350 332928 346384
rect 332608 346294 332678 346350
rect 332734 346294 332802 346350
rect 332858 346294 332928 346350
rect 332608 346226 332928 346294
rect 332608 346170 332678 346226
rect 332734 346170 332802 346226
rect 332858 346170 332928 346226
rect 332608 346102 332928 346170
rect 332608 346046 332678 346102
rect 332734 346046 332802 346102
rect 332858 346046 332928 346102
rect 332608 345978 332928 346046
rect 332608 345922 332678 345978
rect 332734 345922 332802 345978
rect 332858 345922 332928 345978
rect 332608 345888 332928 345922
rect 363328 346350 363648 346384
rect 363328 346294 363398 346350
rect 363454 346294 363522 346350
rect 363578 346294 363648 346350
rect 363328 346226 363648 346294
rect 363328 346170 363398 346226
rect 363454 346170 363522 346226
rect 363578 346170 363648 346226
rect 363328 346102 363648 346170
rect 363328 346046 363398 346102
rect 363454 346046 363522 346102
rect 363578 346046 363648 346102
rect 363328 345978 363648 346046
rect 363328 345922 363398 345978
rect 363454 345922 363522 345978
rect 363578 345922 363648 345978
rect 363328 345888 363648 345922
rect 255808 334350 256128 334384
rect 255808 334294 255878 334350
rect 255934 334294 256002 334350
rect 256058 334294 256128 334350
rect 255808 334226 256128 334294
rect 255808 334170 255878 334226
rect 255934 334170 256002 334226
rect 256058 334170 256128 334226
rect 255808 334102 256128 334170
rect 255808 334046 255878 334102
rect 255934 334046 256002 334102
rect 256058 334046 256128 334102
rect 255808 333978 256128 334046
rect 255808 333922 255878 333978
rect 255934 333922 256002 333978
rect 256058 333922 256128 333978
rect 255808 333888 256128 333922
rect 286528 334350 286848 334384
rect 286528 334294 286598 334350
rect 286654 334294 286722 334350
rect 286778 334294 286848 334350
rect 286528 334226 286848 334294
rect 286528 334170 286598 334226
rect 286654 334170 286722 334226
rect 286778 334170 286848 334226
rect 286528 334102 286848 334170
rect 286528 334046 286598 334102
rect 286654 334046 286722 334102
rect 286778 334046 286848 334102
rect 286528 333978 286848 334046
rect 286528 333922 286598 333978
rect 286654 333922 286722 333978
rect 286778 333922 286848 333978
rect 286528 333888 286848 333922
rect 317248 334350 317568 334384
rect 317248 334294 317318 334350
rect 317374 334294 317442 334350
rect 317498 334294 317568 334350
rect 317248 334226 317568 334294
rect 317248 334170 317318 334226
rect 317374 334170 317442 334226
rect 317498 334170 317568 334226
rect 317248 334102 317568 334170
rect 317248 334046 317318 334102
rect 317374 334046 317442 334102
rect 317498 334046 317568 334102
rect 317248 333978 317568 334046
rect 317248 333922 317318 333978
rect 317374 333922 317442 333978
rect 317498 333922 317568 333978
rect 317248 333888 317568 333922
rect 347968 334350 348288 334384
rect 347968 334294 348038 334350
rect 348094 334294 348162 334350
rect 348218 334294 348288 334350
rect 347968 334226 348288 334294
rect 347968 334170 348038 334226
rect 348094 334170 348162 334226
rect 348218 334170 348288 334226
rect 347968 334102 348288 334170
rect 347968 334046 348038 334102
rect 348094 334046 348162 334102
rect 348218 334046 348288 334102
rect 347968 333978 348288 334046
rect 347968 333922 348038 333978
rect 348094 333922 348162 333978
rect 348218 333922 348288 333978
rect 347968 333888 348288 333922
rect 240448 328350 240768 328384
rect 240448 328294 240518 328350
rect 240574 328294 240642 328350
rect 240698 328294 240768 328350
rect 240448 328226 240768 328294
rect 240448 328170 240518 328226
rect 240574 328170 240642 328226
rect 240698 328170 240768 328226
rect 240448 328102 240768 328170
rect 240448 328046 240518 328102
rect 240574 328046 240642 328102
rect 240698 328046 240768 328102
rect 240448 327978 240768 328046
rect 240448 327922 240518 327978
rect 240574 327922 240642 327978
rect 240698 327922 240768 327978
rect 240448 327888 240768 327922
rect 271168 328350 271488 328384
rect 271168 328294 271238 328350
rect 271294 328294 271362 328350
rect 271418 328294 271488 328350
rect 271168 328226 271488 328294
rect 271168 328170 271238 328226
rect 271294 328170 271362 328226
rect 271418 328170 271488 328226
rect 271168 328102 271488 328170
rect 271168 328046 271238 328102
rect 271294 328046 271362 328102
rect 271418 328046 271488 328102
rect 271168 327978 271488 328046
rect 271168 327922 271238 327978
rect 271294 327922 271362 327978
rect 271418 327922 271488 327978
rect 271168 327888 271488 327922
rect 301888 328350 302208 328384
rect 301888 328294 301958 328350
rect 302014 328294 302082 328350
rect 302138 328294 302208 328350
rect 301888 328226 302208 328294
rect 301888 328170 301958 328226
rect 302014 328170 302082 328226
rect 302138 328170 302208 328226
rect 301888 328102 302208 328170
rect 301888 328046 301958 328102
rect 302014 328046 302082 328102
rect 302138 328046 302208 328102
rect 301888 327978 302208 328046
rect 301888 327922 301958 327978
rect 302014 327922 302082 327978
rect 302138 327922 302208 327978
rect 301888 327888 302208 327922
rect 332608 328350 332928 328384
rect 332608 328294 332678 328350
rect 332734 328294 332802 328350
rect 332858 328294 332928 328350
rect 332608 328226 332928 328294
rect 332608 328170 332678 328226
rect 332734 328170 332802 328226
rect 332858 328170 332928 328226
rect 332608 328102 332928 328170
rect 332608 328046 332678 328102
rect 332734 328046 332802 328102
rect 332858 328046 332928 328102
rect 332608 327978 332928 328046
rect 332608 327922 332678 327978
rect 332734 327922 332802 327978
rect 332858 327922 332928 327978
rect 332608 327888 332928 327922
rect 363328 328350 363648 328384
rect 363328 328294 363398 328350
rect 363454 328294 363522 328350
rect 363578 328294 363648 328350
rect 363328 328226 363648 328294
rect 363328 328170 363398 328226
rect 363454 328170 363522 328226
rect 363578 328170 363648 328226
rect 363328 328102 363648 328170
rect 363328 328046 363398 328102
rect 363454 328046 363522 328102
rect 363578 328046 363648 328102
rect 363328 327978 363648 328046
rect 363328 327922 363398 327978
rect 363454 327922 363522 327978
rect 363578 327922 363648 327978
rect 363328 327888 363648 327922
rect 255808 316350 256128 316384
rect 255808 316294 255878 316350
rect 255934 316294 256002 316350
rect 256058 316294 256128 316350
rect 255808 316226 256128 316294
rect 255808 316170 255878 316226
rect 255934 316170 256002 316226
rect 256058 316170 256128 316226
rect 255808 316102 256128 316170
rect 255808 316046 255878 316102
rect 255934 316046 256002 316102
rect 256058 316046 256128 316102
rect 255808 315978 256128 316046
rect 255808 315922 255878 315978
rect 255934 315922 256002 315978
rect 256058 315922 256128 315978
rect 255808 315888 256128 315922
rect 286528 316350 286848 316384
rect 286528 316294 286598 316350
rect 286654 316294 286722 316350
rect 286778 316294 286848 316350
rect 286528 316226 286848 316294
rect 286528 316170 286598 316226
rect 286654 316170 286722 316226
rect 286778 316170 286848 316226
rect 286528 316102 286848 316170
rect 286528 316046 286598 316102
rect 286654 316046 286722 316102
rect 286778 316046 286848 316102
rect 286528 315978 286848 316046
rect 286528 315922 286598 315978
rect 286654 315922 286722 315978
rect 286778 315922 286848 315978
rect 286528 315888 286848 315922
rect 317248 316350 317568 316384
rect 317248 316294 317318 316350
rect 317374 316294 317442 316350
rect 317498 316294 317568 316350
rect 317248 316226 317568 316294
rect 317248 316170 317318 316226
rect 317374 316170 317442 316226
rect 317498 316170 317568 316226
rect 317248 316102 317568 316170
rect 317248 316046 317318 316102
rect 317374 316046 317442 316102
rect 317498 316046 317568 316102
rect 317248 315978 317568 316046
rect 317248 315922 317318 315978
rect 317374 315922 317442 315978
rect 317498 315922 317568 315978
rect 317248 315888 317568 315922
rect 347968 316350 348288 316384
rect 347968 316294 348038 316350
rect 348094 316294 348162 316350
rect 348218 316294 348288 316350
rect 347968 316226 348288 316294
rect 347968 316170 348038 316226
rect 348094 316170 348162 316226
rect 348218 316170 348288 316226
rect 347968 316102 348288 316170
rect 347968 316046 348038 316102
rect 348094 316046 348162 316102
rect 348218 316046 348288 316102
rect 347968 315978 348288 316046
rect 347968 315922 348038 315978
rect 348094 315922 348162 315978
rect 348218 315922 348288 315978
rect 347968 315888 348288 315922
rect 240448 310350 240768 310384
rect 240448 310294 240518 310350
rect 240574 310294 240642 310350
rect 240698 310294 240768 310350
rect 240448 310226 240768 310294
rect 240448 310170 240518 310226
rect 240574 310170 240642 310226
rect 240698 310170 240768 310226
rect 240448 310102 240768 310170
rect 240448 310046 240518 310102
rect 240574 310046 240642 310102
rect 240698 310046 240768 310102
rect 240448 309978 240768 310046
rect 240448 309922 240518 309978
rect 240574 309922 240642 309978
rect 240698 309922 240768 309978
rect 240448 309888 240768 309922
rect 271168 310350 271488 310384
rect 271168 310294 271238 310350
rect 271294 310294 271362 310350
rect 271418 310294 271488 310350
rect 271168 310226 271488 310294
rect 271168 310170 271238 310226
rect 271294 310170 271362 310226
rect 271418 310170 271488 310226
rect 271168 310102 271488 310170
rect 271168 310046 271238 310102
rect 271294 310046 271362 310102
rect 271418 310046 271488 310102
rect 271168 309978 271488 310046
rect 271168 309922 271238 309978
rect 271294 309922 271362 309978
rect 271418 309922 271488 309978
rect 271168 309888 271488 309922
rect 301888 310350 302208 310384
rect 301888 310294 301958 310350
rect 302014 310294 302082 310350
rect 302138 310294 302208 310350
rect 301888 310226 302208 310294
rect 301888 310170 301958 310226
rect 302014 310170 302082 310226
rect 302138 310170 302208 310226
rect 301888 310102 302208 310170
rect 301888 310046 301958 310102
rect 302014 310046 302082 310102
rect 302138 310046 302208 310102
rect 301888 309978 302208 310046
rect 301888 309922 301958 309978
rect 302014 309922 302082 309978
rect 302138 309922 302208 309978
rect 301888 309888 302208 309922
rect 332608 310350 332928 310384
rect 332608 310294 332678 310350
rect 332734 310294 332802 310350
rect 332858 310294 332928 310350
rect 332608 310226 332928 310294
rect 332608 310170 332678 310226
rect 332734 310170 332802 310226
rect 332858 310170 332928 310226
rect 332608 310102 332928 310170
rect 332608 310046 332678 310102
rect 332734 310046 332802 310102
rect 332858 310046 332928 310102
rect 332608 309978 332928 310046
rect 332608 309922 332678 309978
rect 332734 309922 332802 309978
rect 332858 309922 332928 309978
rect 332608 309888 332928 309922
rect 363328 310350 363648 310384
rect 363328 310294 363398 310350
rect 363454 310294 363522 310350
rect 363578 310294 363648 310350
rect 363328 310226 363648 310294
rect 363328 310170 363398 310226
rect 363454 310170 363522 310226
rect 363578 310170 363648 310226
rect 363328 310102 363648 310170
rect 363328 310046 363398 310102
rect 363454 310046 363522 310102
rect 363578 310046 363648 310102
rect 363328 309978 363648 310046
rect 363328 309922 363398 309978
rect 363454 309922 363522 309978
rect 363578 309922 363648 309978
rect 363328 309888 363648 309922
rect 255808 298350 256128 298384
rect 255808 298294 255878 298350
rect 255934 298294 256002 298350
rect 256058 298294 256128 298350
rect 255808 298226 256128 298294
rect 255808 298170 255878 298226
rect 255934 298170 256002 298226
rect 256058 298170 256128 298226
rect 255808 298102 256128 298170
rect 255808 298046 255878 298102
rect 255934 298046 256002 298102
rect 256058 298046 256128 298102
rect 255808 297978 256128 298046
rect 255808 297922 255878 297978
rect 255934 297922 256002 297978
rect 256058 297922 256128 297978
rect 255808 297888 256128 297922
rect 286528 298350 286848 298384
rect 286528 298294 286598 298350
rect 286654 298294 286722 298350
rect 286778 298294 286848 298350
rect 286528 298226 286848 298294
rect 286528 298170 286598 298226
rect 286654 298170 286722 298226
rect 286778 298170 286848 298226
rect 286528 298102 286848 298170
rect 286528 298046 286598 298102
rect 286654 298046 286722 298102
rect 286778 298046 286848 298102
rect 286528 297978 286848 298046
rect 286528 297922 286598 297978
rect 286654 297922 286722 297978
rect 286778 297922 286848 297978
rect 286528 297888 286848 297922
rect 317248 298350 317568 298384
rect 317248 298294 317318 298350
rect 317374 298294 317442 298350
rect 317498 298294 317568 298350
rect 317248 298226 317568 298294
rect 317248 298170 317318 298226
rect 317374 298170 317442 298226
rect 317498 298170 317568 298226
rect 317248 298102 317568 298170
rect 317248 298046 317318 298102
rect 317374 298046 317442 298102
rect 317498 298046 317568 298102
rect 317248 297978 317568 298046
rect 317248 297922 317318 297978
rect 317374 297922 317442 297978
rect 317498 297922 317568 297978
rect 317248 297888 317568 297922
rect 347968 298350 348288 298384
rect 347968 298294 348038 298350
rect 348094 298294 348162 298350
rect 348218 298294 348288 298350
rect 347968 298226 348288 298294
rect 347968 298170 348038 298226
rect 348094 298170 348162 298226
rect 348218 298170 348288 298226
rect 347968 298102 348288 298170
rect 347968 298046 348038 298102
rect 348094 298046 348162 298102
rect 348218 298046 348288 298102
rect 347968 297978 348288 298046
rect 347968 297922 348038 297978
rect 348094 297922 348162 297978
rect 348218 297922 348288 297978
rect 347968 297888 348288 297922
rect 240448 292350 240768 292384
rect 240448 292294 240518 292350
rect 240574 292294 240642 292350
rect 240698 292294 240768 292350
rect 240448 292226 240768 292294
rect 240448 292170 240518 292226
rect 240574 292170 240642 292226
rect 240698 292170 240768 292226
rect 240448 292102 240768 292170
rect 240448 292046 240518 292102
rect 240574 292046 240642 292102
rect 240698 292046 240768 292102
rect 240448 291978 240768 292046
rect 240448 291922 240518 291978
rect 240574 291922 240642 291978
rect 240698 291922 240768 291978
rect 240448 291888 240768 291922
rect 271168 292350 271488 292384
rect 271168 292294 271238 292350
rect 271294 292294 271362 292350
rect 271418 292294 271488 292350
rect 271168 292226 271488 292294
rect 271168 292170 271238 292226
rect 271294 292170 271362 292226
rect 271418 292170 271488 292226
rect 271168 292102 271488 292170
rect 271168 292046 271238 292102
rect 271294 292046 271362 292102
rect 271418 292046 271488 292102
rect 271168 291978 271488 292046
rect 271168 291922 271238 291978
rect 271294 291922 271362 291978
rect 271418 291922 271488 291978
rect 271168 291888 271488 291922
rect 301888 292350 302208 292384
rect 301888 292294 301958 292350
rect 302014 292294 302082 292350
rect 302138 292294 302208 292350
rect 301888 292226 302208 292294
rect 301888 292170 301958 292226
rect 302014 292170 302082 292226
rect 302138 292170 302208 292226
rect 301888 292102 302208 292170
rect 301888 292046 301958 292102
rect 302014 292046 302082 292102
rect 302138 292046 302208 292102
rect 301888 291978 302208 292046
rect 301888 291922 301958 291978
rect 302014 291922 302082 291978
rect 302138 291922 302208 291978
rect 301888 291888 302208 291922
rect 332608 292350 332928 292384
rect 332608 292294 332678 292350
rect 332734 292294 332802 292350
rect 332858 292294 332928 292350
rect 332608 292226 332928 292294
rect 332608 292170 332678 292226
rect 332734 292170 332802 292226
rect 332858 292170 332928 292226
rect 332608 292102 332928 292170
rect 332608 292046 332678 292102
rect 332734 292046 332802 292102
rect 332858 292046 332928 292102
rect 332608 291978 332928 292046
rect 332608 291922 332678 291978
rect 332734 291922 332802 291978
rect 332858 291922 332928 291978
rect 332608 291888 332928 291922
rect 363328 292350 363648 292384
rect 363328 292294 363398 292350
rect 363454 292294 363522 292350
rect 363578 292294 363648 292350
rect 363328 292226 363648 292294
rect 363328 292170 363398 292226
rect 363454 292170 363522 292226
rect 363578 292170 363648 292226
rect 363328 292102 363648 292170
rect 363328 292046 363398 292102
rect 363454 292046 363522 292102
rect 363578 292046 363648 292102
rect 363328 291978 363648 292046
rect 363328 291922 363398 291978
rect 363454 291922 363522 291978
rect 363578 291922 363648 291978
rect 363328 291888 363648 291922
rect 255808 280350 256128 280384
rect 255808 280294 255878 280350
rect 255934 280294 256002 280350
rect 256058 280294 256128 280350
rect 255808 280226 256128 280294
rect 255808 280170 255878 280226
rect 255934 280170 256002 280226
rect 256058 280170 256128 280226
rect 255808 280102 256128 280170
rect 255808 280046 255878 280102
rect 255934 280046 256002 280102
rect 256058 280046 256128 280102
rect 255808 279978 256128 280046
rect 255808 279922 255878 279978
rect 255934 279922 256002 279978
rect 256058 279922 256128 279978
rect 255808 279888 256128 279922
rect 286528 280350 286848 280384
rect 286528 280294 286598 280350
rect 286654 280294 286722 280350
rect 286778 280294 286848 280350
rect 286528 280226 286848 280294
rect 286528 280170 286598 280226
rect 286654 280170 286722 280226
rect 286778 280170 286848 280226
rect 286528 280102 286848 280170
rect 286528 280046 286598 280102
rect 286654 280046 286722 280102
rect 286778 280046 286848 280102
rect 286528 279978 286848 280046
rect 286528 279922 286598 279978
rect 286654 279922 286722 279978
rect 286778 279922 286848 279978
rect 286528 279888 286848 279922
rect 317248 280350 317568 280384
rect 317248 280294 317318 280350
rect 317374 280294 317442 280350
rect 317498 280294 317568 280350
rect 317248 280226 317568 280294
rect 317248 280170 317318 280226
rect 317374 280170 317442 280226
rect 317498 280170 317568 280226
rect 317248 280102 317568 280170
rect 317248 280046 317318 280102
rect 317374 280046 317442 280102
rect 317498 280046 317568 280102
rect 317248 279978 317568 280046
rect 317248 279922 317318 279978
rect 317374 279922 317442 279978
rect 317498 279922 317568 279978
rect 317248 279888 317568 279922
rect 347968 280350 348288 280384
rect 347968 280294 348038 280350
rect 348094 280294 348162 280350
rect 348218 280294 348288 280350
rect 347968 280226 348288 280294
rect 347968 280170 348038 280226
rect 348094 280170 348162 280226
rect 348218 280170 348288 280226
rect 347968 280102 348288 280170
rect 347968 280046 348038 280102
rect 348094 280046 348162 280102
rect 348218 280046 348288 280102
rect 347968 279978 348288 280046
rect 347968 279922 348038 279978
rect 348094 279922 348162 279978
rect 348218 279922 348288 279978
rect 347968 279888 348288 279922
rect 240448 274350 240768 274384
rect 240448 274294 240518 274350
rect 240574 274294 240642 274350
rect 240698 274294 240768 274350
rect 240448 274226 240768 274294
rect 240448 274170 240518 274226
rect 240574 274170 240642 274226
rect 240698 274170 240768 274226
rect 240448 274102 240768 274170
rect 240448 274046 240518 274102
rect 240574 274046 240642 274102
rect 240698 274046 240768 274102
rect 240448 273978 240768 274046
rect 240448 273922 240518 273978
rect 240574 273922 240642 273978
rect 240698 273922 240768 273978
rect 240448 273888 240768 273922
rect 271168 274350 271488 274384
rect 271168 274294 271238 274350
rect 271294 274294 271362 274350
rect 271418 274294 271488 274350
rect 271168 274226 271488 274294
rect 271168 274170 271238 274226
rect 271294 274170 271362 274226
rect 271418 274170 271488 274226
rect 271168 274102 271488 274170
rect 271168 274046 271238 274102
rect 271294 274046 271362 274102
rect 271418 274046 271488 274102
rect 271168 273978 271488 274046
rect 271168 273922 271238 273978
rect 271294 273922 271362 273978
rect 271418 273922 271488 273978
rect 271168 273888 271488 273922
rect 301888 274350 302208 274384
rect 301888 274294 301958 274350
rect 302014 274294 302082 274350
rect 302138 274294 302208 274350
rect 301888 274226 302208 274294
rect 301888 274170 301958 274226
rect 302014 274170 302082 274226
rect 302138 274170 302208 274226
rect 301888 274102 302208 274170
rect 301888 274046 301958 274102
rect 302014 274046 302082 274102
rect 302138 274046 302208 274102
rect 301888 273978 302208 274046
rect 301888 273922 301958 273978
rect 302014 273922 302082 273978
rect 302138 273922 302208 273978
rect 301888 273888 302208 273922
rect 332608 274350 332928 274384
rect 332608 274294 332678 274350
rect 332734 274294 332802 274350
rect 332858 274294 332928 274350
rect 332608 274226 332928 274294
rect 332608 274170 332678 274226
rect 332734 274170 332802 274226
rect 332858 274170 332928 274226
rect 332608 274102 332928 274170
rect 332608 274046 332678 274102
rect 332734 274046 332802 274102
rect 332858 274046 332928 274102
rect 332608 273978 332928 274046
rect 332608 273922 332678 273978
rect 332734 273922 332802 273978
rect 332858 273922 332928 273978
rect 332608 273888 332928 273922
rect 363328 274350 363648 274384
rect 363328 274294 363398 274350
rect 363454 274294 363522 274350
rect 363578 274294 363648 274350
rect 363328 274226 363648 274294
rect 363328 274170 363398 274226
rect 363454 274170 363522 274226
rect 363578 274170 363648 274226
rect 363328 274102 363648 274170
rect 363328 274046 363398 274102
rect 363454 274046 363522 274102
rect 363578 274046 363648 274102
rect 363328 273978 363648 274046
rect 363328 273922 363398 273978
rect 363454 273922 363522 273978
rect 363578 273922 363648 273978
rect 363328 273888 363648 273922
rect 255808 262350 256128 262384
rect 255808 262294 255878 262350
rect 255934 262294 256002 262350
rect 256058 262294 256128 262350
rect 255808 262226 256128 262294
rect 255808 262170 255878 262226
rect 255934 262170 256002 262226
rect 256058 262170 256128 262226
rect 255808 262102 256128 262170
rect 255808 262046 255878 262102
rect 255934 262046 256002 262102
rect 256058 262046 256128 262102
rect 255808 261978 256128 262046
rect 255808 261922 255878 261978
rect 255934 261922 256002 261978
rect 256058 261922 256128 261978
rect 255808 261888 256128 261922
rect 286528 262350 286848 262384
rect 286528 262294 286598 262350
rect 286654 262294 286722 262350
rect 286778 262294 286848 262350
rect 286528 262226 286848 262294
rect 286528 262170 286598 262226
rect 286654 262170 286722 262226
rect 286778 262170 286848 262226
rect 286528 262102 286848 262170
rect 286528 262046 286598 262102
rect 286654 262046 286722 262102
rect 286778 262046 286848 262102
rect 286528 261978 286848 262046
rect 286528 261922 286598 261978
rect 286654 261922 286722 261978
rect 286778 261922 286848 261978
rect 286528 261888 286848 261922
rect 317248 262350 317568 262384
rect 317248 262294 317318 262350
rect 317374 262294 317442 262350
rect 317498 262294 317568 262350
rect 317248 262226 317568 262294
rect 317248 262170 317318 262226
rect 317374 262170 317442 262226
rect 317498 262170 317568 262226
rect 317248 262102 317568 262170
rect 317248 262046 317318 262102
rect 317374 262046 317442 262102
rect 317498 262046 317568 262102
rect 317248 261978 317568 262046
rect 317248 261922 317318 261978
rect 317374 261922 317442 261978
rect 317498 261922 317568 261978
rect 317248 261888 317568 261922
rect 347968 262350 348288 262384
rect 347968 262294 348038 262350
rect 348094 262294 348162 262350
rect 348218 262294 348288 262350
rect 347968 262226 348288 262294
rect 347968 262170 348038 262226
rect 348094 262170 348162 262226
rect 348218 262170 348288 262226
rect 347968 262102 348288 262170
rect 347968 262046 348038 262102
rect 348094 262046 348162 262102
rect 348218 262046 348288 262102
rect 347968 261978 348288 262046
rect 347968 261922 348038 261978
rect 348094 261922 348162 261978
rect 348218 261922 348288 261978
rect 347968 261888 348288 261922
rect 358652 257878 358708 257888
rect 237916 210832 237972 210842
rect 251178 256350 251798 257490
rect 251178 256294 251274 256350
rect 251330 256294 251398 256350
rect 251454 256294 251522 256350
rect 251578 256294 251646 256350
rect 251702 256294 251798 256350
rect 251178 256226 251798 256294
rect 251178 256170 251274 256226
rect 251330 256170 251398 256226
rect 251454 256170 251522 256226
rect 251578 256170 251646 256226
rect 251702 256170 251798 256226
rect 251178 256102 251798 256170
rect 251178 256046 251274 256102
rect 251330 256046 251398 256102
rect 251454 256046 251522 256102
rect 251578 256046 251646 256102
rect 251702 256046 251798 256102
rect 251178 255978 251798 256046
rect 251178 255922 251274 255978
rect 251330 255922 251398 255978
rect 251454 255922 251522 255978
rect 251578 255922 251646 255978
rect 251702 255922 251798 255978
rect 251178 238350 251798 255922
rect 251916 253652 251972 253662
rect 251916 252838 251972 253596
rect 251916 252772 251972 252782
rect 252588 253652 252644 253662
rect 252588 252478 252644 253596
rect 252588 252412 252644 252422
rect 251178 238294 251274 238350
rect 251330 238294 251398 238350
rect 251454 238294 251522 238350
rect 251578 238294 251646 238350
rect 251702 238294 251798 238350
rect 251178 238226 251798 238294
rect 251178 238170 251274 238226
rect 251330 238170 251398 238226
rect 251454 238170 251522 238226
rect 251578 238170 251646 238226
rect 251702 238170 251798 238226
rect 251178 238102 251798 238170
rect 251178 238046 251274 238102
rect 251330 238046 251398 238102
rect 251454 238046 251522 238102
rect 251578 238046 251646 238102
rect 251702 238046 251798 238102
rect 251178 237978 251798 238046
rect 251178 237922 251274 237978
rect 251330 237922 251398 237978
rect 251454 237922 251522 237978
rect 251578 237922 251646 237978
rect 251702 237922 251798 237978
rect 251178 220350 251798 237922
rect 251178 220294 251274 220350
rect 251330 220294 251398 220350
rect 251454 220294 251522 220350
rect 251578 220294 251646 220350
rect 251702 220294 251798 220350
rect 251178 220226 251798 220294
rect 251178 220170 251274 220226
rect 251330 220170 251398 220226
rect 251454 220170 251522 220226
rect 251578 220170 251646 220226
rect 251702 220170 251798 220226
rect 251178 220102 251798 220170
rect 251178 220046 251274 220102
rect 251330 220046 251398 220102
rect 251454 220046 251522 220102
rect 251578 220046 251646 220102
rect 251702 220046 251798 220102
rect 251178 219978 251798 220046
rect 251178 219922 251274 219978
rect 251330 219922 251398 219978
rect 251454 219922 251522 219978
rect 251578 219922 251646 219978
rect 251702 219922 251798 219978
rect 251178 210462 251798 219922
rect 254898 244350 255518 257490
rect 269276 257348 269332 257358
rect 258860 253652 258916 253662
rect 258860 252658 258916 253596
rect 258860 252592 258916 252602
rect 259756 253652 259812 253662
rect 259756 252298 259812 253596
rect 259756 252232 259812 252242
rect 260652 253652 260708 253662
rect 260652 252118 260708 253596
rect 260652 252052 260708 252062
rect 254898 244294 254994 244350
rect 255050 244294 255118 244350
rect 255174 244294 255242 244350
rect 255298 244294 255366 244350
rect 255422 244294 255518 244350
rect 254898 244226 255518 244294
rect 254898 244170 254994 244226
rect 255050 244170 255118 244226
rect 255174 244170 255242 244226
rect 255298 244170 255366 244226
rect 255422 244170 255518 244226
rect 254898 244102 255518 244170
rect 254898 244046 254994 244102
rect 255050 244046 255118 244102
rect 255174 244046 255242 244102
rect 255298 244046 255366 244102
rect 255422 244046 255518 244102
rect 254898 243978 255518 244046
rect 254898 243922 254994 243978
rect 255050 243922 255118 243978
rect 255174 243922 255242 243978
rect 255298 243922 255366 243978
rect 255422 243922 255518 243978
rect 254898 226350 255518 243922
rect 254898 226294 254994 226350
rect 255050 226294 255118 226350
rect 255174 226294 255242 226350
rect 255298 226294 255366 226350
rect 255422 226294 255518 226350
rect 254898 226226 255518 226294
rect 254898 226170 254994 226226
rect 255050 226170 255118 226226
rect 255174 226170 255242 226226
rect 255298 226170 255366 226226
rect 255422 226170 255518 226226
rect 254898 226102 255518 226170
rect 254898 226046 254994 226102
rect 255050 226046 255118 226102
rect 255174 226046 255242 226102
rect 255298 226046 255366 226102
rect 255422 226046 255518 226102
rect 254898 225978 255518 226046
rect 254898 225922 254994 225978
rect 255050 225922 255118 225978
rect 255174 225922 255242 225978
rect 255298 225922 255366 225978
rect 255422 225922 255518 225978
rect 254898 210462 255518 225922
rect 267148 249396 267204 249406
rect 234444 209906 234500 209916
rect 231420 209682 231476 209692
rect 229964 209570 230020 209580
rect 228396 209458 228452 209468
rect 226604 209346 226660 209356
rect 75168 202350 75488 202384
rect 75168 202294 75238 202350
rect 75294 202294 75362 202350
rect 75418 202294 75488 202350
rect 75168 202226 75488 202294
rect 75168 202170 75238 202226
rect 75294 202170 75362 202226
rect 75418 202170 75488 202226
rect 75168 202102 75488 202170
rect 75168 202046 75238 202102
rect 75294 202046 75362 202102
rect 75418 202046 75488 202102
rect 75168 201978 75488 202046
rect 75168 201922 75238 201978
rect 75294 201922 75362 201978
rect 75418 201922 75488 201978
rect 75168 201888 75488 201922
rect 105888 202350 106208 202384
rect 105888 202294 105958 202350
rect 106014 202294 106082 202350
rect 106138 202294 106208 202350
rect 105888 202226 106208 202294
rect 105888 202170 105958 202226
rect 106014 202170 106082 202226
rect 106138 202170 106208 202226
rect 105888 202102 106208 202170
rect 105888 202046 105958 202102
rect 106014 202046 106082 202102
rect 106138 202046 106208 202102
rect 105888 201978 106208 202046
rect 105888 201922 105958 201978
rect 106014 201922 106082 201978
rect 106138 201922 106208 201978
rect 105888 201888 106208 201922
rect 136608 202350 136928 202384
rect 136608 202294 136678 202350
rect 136734 202294 136802 202350
rect 136858 202294 136928 202350
rect 136608 202226 136928 202294
rect 136608 202170 136678 202226
rect 136734 202170 136802 202226
rect 136858 202170 136928 202226
rect 136608 202102 136928 202170
rect 136608 202046 136678 202102
rect 136734 202046 136802 202102
rect 136858 202046 136928 202102
rect 136608 201978 136928 202046
rect 136608 201922 136678 201978
rect 136734 201922 136802 201978
rect 136858 201922 136928 201978
rect 136608 201888 136928 201922
rect 167328 202350 167648 202384
rect 167328 202294 167398 202350
rect 167454 202294 167522 202350
rect 167578 202294 167648 202350
rect 167328 202226 167648 202294
rect 167328 202170 167398 202226
rect 167454 202170 167522 202226
rect 167578 202170 167648 202226
rect 167328 202102 167648 202170
rect 167328 202046 167398 202102
rect 167454 202046 167522 202102
rect 167578 202046 167648 202102
rect 167328 201978 167648 202046
rect 167328 201922 167398 201978
rect 167454 201922 167522 201978
rect 167578 201922 167648 201978
rect 167328 201888 167648 201922
rect 198048 202350 198368 202384
rect 198048 202294 198118 202350
rect 198174 202294 198242 202350
rect 198298 202294 198368 202350
rect 198048 202226 198368 202294
rect 198048 202170 198118 202226
rect 198174 202170 198242 202226
rect 198298 202170 198368 202226
rect 198048 202102 198368 202170
rect 198048 202046 198118 202102
rect 198174 202046 198242 202102
rect 198298 202046 198368 202102
rect 198048 201978 198368 202046
rect 198048 201922 198118 201978
rect 198174 201922 198242 201978
rect 198298 201922 198368 201978
rect 198048 201888 198368 201922
rect 228768 202350 229088 202384
rect 228768 202294 228838 202350
rect 228894 202294 228962 202350
rect 229018 202294 229088 202350
rect 228768 202226 229088 202294
rect 228768 202170 228838 202226
rect 228894 202170 228962 202226
rect 229018 202170 229088 202226
rect 228768 202102 229088 202170
rect 228768 202046 228838 202102
rect 228894 202046 228962 202102
rect 229018 202046 229088 202102
rect 228768 201978 229088 202046
rect 228768 201922 228838 201978
rect 228894 201922 228962 201978
rect 229018 201922 229088 201978
rect 228768 201888 229088 201922
rect 259488 202350 259808 202384
rect 259488 202294 259558 202350
rect 259614 202294 259682 202350
rect 259738 202294 259808 202350
rect 259488 202226 259808 202294
rect 259488 202170 259558 202226
rect 259614 202170 259682 202226
rect 259738 202170 259808 202226
rect 259488 202102 259808 202170
rect 259488 202046 259558 202102
rect 259614 202046 259682 202102
rect 259738 202046 259808 202102
rect 259488 201978 259808 202046
rect 259488 201922 259558 201978
rect 259614 201922 259682 201978
rect 259738 201922 259808 201978
rect 259488 201888 259808 201922
rect 59808 190350 60128 190384
rect 59808 190294 59878 190350
rect 59934 190294 60002 190350
rect 60058 190294 60128 190350
rect 59808 190226 60128 190294
rect 59808 190170 59878 190226
rect 59934 190170 60002 190226
rect 60058 190170 60128 190226
rect 59808 190102 60128 190170
rect 59808 190046 59878 190102
rect 59934 190046 60002 190102
rect 60058 190046 60128 190102
rect 59808 189978 60128 190046
rect 59808 189922 59878 189978
rect 59934 189922 60002 189978
rect 60058 189922 60128 189978
rect 59808 189888 60128 189922
rect 90528 190350 90848 190384
rect 90528 190294 90598 190350
rect 90654 190294 90722 190350
rect 90778 190294 90848 190350
rect 90528 190226 90848 190294
rect 90528 190170 90598 190226
rect 90654 190170 90722 190226
rect 90778 190170 90848 190226
rect 90528 190102 90848 190170
rect 90528 190046 90598 190102
rect 90654 190046 90722 190102
rect 90778 190046 90848 190102
rect 90528 189978 90848 190046
rect 90528 189922 90598 189978
rect 90654 189922 90722 189978
rect 90778 189922 90848 189978
rect 90528 189888 90848 189922
rect 121248 190350 121568 190384
rect 121248 190294 121318 190350
rect 121374 190294 121442 190350
rect 121498 190294 121568 190350
rect 121248 190226 121568 190294
rect 121248 190170 121318 190226
rect 121374 190170 121442 190226
rect 121498 190170 121568 190226
rect 121248 190102 121568 190170
rect 121248 190046 121318 190102
rect 121374 190046 121442 190102
rect 121498 190046 121568 190102
rect 121248 189978 121568 190046
rect 121248 189922 121318 189978
rect 121374 189922 121442 189978
rect 121498 189922 121568 189978
rect 121248 189888 121568 189922
rect 151968 190350 152288 190384
rect 151968 190294 152038 190350
rect 152094 190294 152162 190350
rect 152218 190294 152288 190350
rect 151968 190226 152288 190294
rect 151968 190170 152038 190226
rect 152094 190170 152162 190226
rect 152218 190170 152288 190226
rect 151968 190102 152288 190170
rect 151968 190046 152038 190102
rect 152094 190046 152162 190102
rect 152218 190046 152288 190102
rect 151968 189978 152288 190046
rect 151968 189922 152038 189978
rect 152094 189922 152162 189978
rect 152218 189922 152288 189978
rect 151968 189888 152288 189922
rect 182688 190350 183008 190384
rect 182688 190294 182758 190350
rect 182814 190294 182882 190350
rect 182938 190294 183008 190350
rect 182688 190226 183008 190294
rect 182688 190170 182758 190226
rect 182814 190170 182882 190226
rect 182938 190170 183008 190226
rect 182688 190102 183008 190170
rect 182688 190046 182758 190102
rect 182814 190046 182882 190102
rect 182938 190046 183008 190102
rect 182688 189978 183008 190046
rect 182688 189922 182758 189978
rect 182814 189922 182882 189978
rect 182938 189922 183008 189978
rect 182688 189888 183008 189922
rect 213408 190350 213728 190384
rect 213408 190294 213478 190350
rect 213534 190294 213602 190350
rect 213658 190294 213728 190350
rect 213408 190226 213728 190294
rect 213408 190170 213478 190226
rect 213534 190170 213602 190226
rect 213658 190170 213728 190226
rect 213408 190102 213728 190170
rect 213408 190046 213478 190102
rect 213534 190046 213602 190102
rect 213658 190046 213728 190102
rect 213408 189978 213728 190046
rect 213408 189922 213478 189978
rect 213534 189922 213602 189978
rect 213658 189922 213728 189978
rect 213408 189888 213728 189922
rect 244128 190350 244448 190384
rect 244128 190294 244198 190350
rect 244254 190294 244322 190350
rect 244378 190294 244448 190350
rect 244128 190226 244448 190294
rect 244128 190170 244198 190226
rect 244254 190170 244322 190226
rect 244378 190170 244448 190226
rect 244128 190102 244448 190170
rect 244128 190046 244198 190102
rect 244254 190046 244322 190102
rect 244378 190046 244448 190102
rect 244128 189978 244448 190046
rect 244128 189922 244198 189978
rect 244254 189922 244322 189978
rect 244378 189922 244448 189978
rect 244128 189888 244448 189922
rect 75168 184350 75488 184384
rect 75168 184294 75238 184350
rect 75294 184294 75362 184350
rect 75418 184294 75488 184350
rect 75168 184226 75488 184294
rect 75168 184170 75238 184226
rect 75294 184170 75362 184226
rect 75418 184170 75488 184226
rect 75168 184102 75488 184170
rect 75168 184046 75238 184102
rect 75294 184046 75362 184102
rect 75418 184046 75488 184102
rect 75168 183978 75488 184046
rect 75168 183922 75238 183978
rect 75294 183922 75362 183978
rect 75418 183922 75488 183978
rect 75168 183888 75488 183922
rect 105888 184350 106208 184384
rect 105888 184294 105958 184350
rect 106014 184294 106082 184350
rect 106138 184294 106208 184350
rect 105888 184226 106208 184294
rect 105888 184170 105958 184226
rect 106014 184170 106082 184226
rect 106138 184170 106208 184226
rect 105888 184102 106208 184170
rect 105888 184046 105958 184102
rect 106014 184046 106082 184102
rect 106138 184046 106208 184102
rect 105888 183978 106208 184046
rect 105888 183922 105958 183978
rect 106014 183922 106082 183978
rect 106138 183922 106208 183978
rect 105888 183888 106208 183922
rect 136608 184350 136928 184384
rect 136608 184294 136678 184350
rect 136734 184294 136802 184350
rect 136858 184294 136928 184350
rect 136608 184226 136928 184294
rect 136608 184170 136678 184226
rect 136734 184170 136802 184226
rect 136858 184170 136928 184226
rect 136608 184102 136928 184170
rect 136608 184046 136678 184102
rect 136734 184046 136802 184102
rect 136858 184046 136928 184102
rect 136608 183978 136928 184046
rect 136608 183922 136678 183978
rect 136734 183922 136802 183978
rect 136858 183922 136928 183978
rect 136608 183888 136928 183922
rect 167328 184350 167648 184384
rect 167328 184294 167398 184350
rect 167454 184294 167522 184350
rect 167578 184294 167648 184350
rect 167328 184226 167648 184294
rect 167328 184170 167398 184226
rect 167454 184170 167522 184226
rect 167578 184170 167648 184226
rect 167328 184102 167648 184170
rect 167328 184046 167398 184102
rect 167454 184046 167522 184102
rect 167578 184046 167648 184102
rect 167328 183978 167648 184046
rect 167328 183922 167398 183978
rect 167454 183922 167522 183978
rect 167578 183922 167648 183978
rect 167328 183888 167648 183922
rect 198048 184350 198368 184384
rect 198048 184294 198118 184350
rect 198174 184294 198242 184350
rect 198298 184294 198368 184350
rect 198048 184226 198368 184294
rect 198048 184170 198118 184226
rect 198174 184170 198242 184226
rect 198298 184170 198368 184226
rect 198048 184102 198368 184170
rect 198048 184046 198118 184102
rect 198174 184046 198242 184102
rect 198298 184046 198368 184102
rect 198048 183978 198368 184046
rect 198048 183922 198118 183978
rect 198174 183922 198242 183978
rect 198298 183922 198368 183978
rect 198048 183888 198368 183922
rect 228768 184350 229088 184384
rect 228768 184294 228838 184350
rect 228894 184294 228962 184350
rect 229018 184294 229088 184350
rect 228768 184226 229088 184294
rect 228768 184170 228838 184226
rect 228894 184170 228962 184226
rect 229018 184170 229088 184226
rect 228768 184102 229088 184170
rect 228768 184046 228838 184102
rect 228894 184046 228962 184102
rect 229018 184046 229088 184102
rect 228768 183978 229088 184046
rect 228768 183922 228838 183978
rect 228894 183922 228962 183978
rect 229018 183922 229088 183978
rect 228768 183888 229088 183922
rect 259488 184350 259808 184384
rect 259488 184294 259558 184350
rect 259614 184294 259682 184350
rect 259738 184294 259808 184350
rect 259488 184226 259808 184294
rect 259488 184170 259558 184226
rect 259614 184170 259682 184226
rect 259738 184170 259808 184226
rect 259488 184102 259808 184170
rect 259488 184046 259558 184102
rect 259614 184046 259682 184102
rect 259738 184046 259808 184102
rect 259488 183978 259808 184046
rect 259488 183922 259558 183978
rect 259614 183922 259682 183978
rect 259738 183922 259808 183978
rect 259488 183888 259808 183922
rect 59808 172350 60128 172384
rect 59808 172294 59878 172350
rect 59934 172294 60002 172350
rect 60058 172294 60128 172350
rect 59808 172226 60128 172294
rect 59808 172170 59878 172226
rect 59934 172170 60002 172226
rect 60058 172170 60128 172226
rect 59808 172102 60128 172170
rect 59808 172046 59878 172102
rect 59934 172046 60002 172102
rect 60058 172046 60128 172102
rect 59808 171978 60128 172046
rect 59808 171922 59878 171978
rect 59934 171922 60002 171978
rect 60058 171922 60128 171978
rect 59808 171888 60128 171922
rect 90528 172350 90848 172384
rect 90528 172294 90598 172350
rect 90654 172294 90722 172350
rect 90778 172294 90848 172350
rect 90528 172226 90848 172294
rect 90528 172170 90598 172226
rect 90654 172170 90722 172226
rect 90778 172170 90848 172226
rect 90528 172102 90848 172170
rect 90528 172046 90598 172102
rect 90654 172046 90722 172102
rect 90778 172046 90848 172102
rect 90528 171978 90848 172046
rect 90528 171922 90598 171978
rect 90654 171922 90722 171978
rect 90778 171922 90848 171978
rect 90528 171888 90848 171922
rect 121248 172350 121568 172384
rect 121248 172294 121318 172350
rect 121374 172294 121442 172350
rect 121498 172294 121568 172350
rect 121248 172226 121568 172294
rect 121248 172170 121318 172226
rect 121374 172170 121442 172226
rect 121498 172170 121568 172226
rect 121248 172102 121568 172170
rect 121248 172046 121318 172102
rect 121374 172046 121442 172102
rect 121498 172046 121568 172102
rect 121248 171978 121568 172046
rect 121248 171922 121318 171978
rect 121374 171922 121442 171978
rect 121498 171922 121568 171978
rect 121248 171888 121568 171922
rect 151968 172350 152288 172384
rect 151968 172294 152038 172350
rect 152094 172294 152162 172350
rect 152218 172294 152288 172350
rect 151968 172226 152288 172294
rect 151968 172170 152038 172226
rect 152094 172170 152162 172226
rect 152218 172170 152288 172226
rect 151968 172102 152288 172170
rect 151968 172046 152038 172102
rect 152094 172046 152162 172102
rect 152218 172046 152288 172102
rect 151968 171978 152288 172046
rect 151968 171922 152038 171978
rect 152094 171922 152162 171978
rect 152218 171922 152288 171978
rect 151968 171888 152288 171922
rect 182688 172350 183008 172384
rect 182688 172294 182758 172350
rect 182814 172294 182882 172350
rect 182938 172294 183008 172350
rect 182688 172226 183008 172294
rect 182688 172170 182758 172226
rect 182814 172170 182882 172226
rect 182938 172170 183008 172226
rect 182688 172102 183008 172170
rect 182688 172046 182758 172102
rect 182814 172046 182882 172102
rect 182938 172046 183008 172102
rect 182688 171978 183008 172046
rect 182688 171922 182758 171978
rect 182814 171922 182882 171978
rect 182938 171922 183008 171978
rect 182688 171888 183008 171922
rect 213408 172350 213728 172384
rect 213408 172294 213478 172350
rect 213534 172294 213602 172350
rect 213658 172294 213728 172350
rect 213408 172226 213728 172294
rect 213408 172170 213478 172226
rect 213534 172170 213602 172226
rect 213658 172170 213728 172226
rect 213408 172102 213728 172170
rect 213408 172046 213478 172102
rect 213534 172046 213602 172102
rect 213658 172046 213728 172102
rect 213408 171978 213728 172046
rect 213408 171922 213478 171978
rect 213534 171922 213602 171978
rect 213658 171922 213728 171978
rect 213408 171888 213728 171922
rect 244128 172350 244448 172384
rect 244128 172294 244198 172350
rect 244254 172294 244322 172350
rect 244378 172294 244448 172350
rect 244128 172226 244448 172294
rect 244128 172170 244198 172226
rect 244254 172170 244322 172226
rect 244378 172170 244448 172226
rect 244128 172102 244448 172170
rect 244128 172046 244198 172102
rect 244254 172046 244322 172102
rect 244378 172046 244448 172102
rect 244128 171978 244448 172046
rect 244128 171922 244198 171978
rect 244254 171922 244322 171978
rect 244378 171922 244448 171978
rect 244128 171888 244448 171922
rect 75168 166350 75488 166384
rect 75168 166294 75238 166350
rect 75294 166294 75362 166350
rect 75418 166294 75488 166350
rect 75168 166226 75488 166294
rect 75168 166170 75238 166226
rect 75294 166170 75362 166226
rect 75418 166170 75488 166226
rect 75168 166102 75488 166170
rect 75168 166046 75238 166102
rect 75294 166046 75362 166102
rect 75418 166046 75488 166102
rect 75168 165978 75488 166046
rect 75168 165922 75238 165978
rect 75294 165922 75362 165978
rect 75418 165922 75488 165978
rect 75168 165888 75488 165922
rect 105888 166350 106208 166384
rect 105888 166294 105958 166350
rect 106014 166294 106082 166350
rect 106138 166294 106208 166350
rect 105888 166226 106208 166294
rect 105888 166170 105958 166226
rect 106014 166170 106082 166226
rect 106138 166170 106208 166226
rect 105888 166102 106208 166170
rect 105888 166046 105958 166102
rect 106014 166046 106082 166102
rect 106138 166046 106208 166102
rect 105888 165978 106208 166046
rect 105888 165922 105958 165978
rect 106014 165922 106082 165978
rect 106138 165922 106208 165978
rect 105888 165888 106208 165922
rect 136608 166350 136928 166384
rect 136608 166294 136678 166350
rect 136734 166294 136802 166350
rect 136858 166294 136928 166350
rect 136608 166226 136928 166294
rect 136608 166170 136678 166226
rect 136734 166170 136802 166226
rect 136858 166170 136928 166226
rect 136608 166102 136928 166170
rect 136608 166046 136678 166102
rect 136734 166046 136802 166102
rect 136858 166046 136928 166102
rect 136608 165978 136928 166046
rect 136608 165922 136678 165978
rect 136734 165922 136802 165978
rect 136858 165922 136928 165978
rect 136608 165888 136928 165922
rect 167328 166350 167648 166384
rect 167328 166294 167398 166350
rect 167454 166294 167522 166350
rect 167578 166294 167648 166350
rect 167328 166226 167648 166294
rect 167328 166170 167398 166226
rect 167454 166170 167522 166226
rect 167578 166170 167648 166226
rect 167328 166102 167648 166170
rect 167328 166046 167398 166102
rect 167454 166046 167522 166102
rect 167578 166046 167648 166102
rect 167328 165978 167648 166046
rect 167328 165922 167398 165978
rect 167454 165922 167522 165978
rect 167578 165922 167648 165978
rect 167328 165888 167648 165922
rect 198048 166350 198368 166384
rect 198048 166294 198118 166350
rect 198174 166294 198242 166350
rect 198298 166294 198368 166350
rect 198048 166226 198368 166294
rect 198048 166170 198118 166226
rect 198174 166170 198242 166226
rect 198298 166170 198368 166226
rect 198048 166102 198368 166170
rect 198048 166046 198118 166102
rect 198174 166046 198242 166102
rect 198298 166046 198368 166102
rect 198048 165978 198368 166046
rect 198048 165922 198118 165978
rect 198174 165922 198242 165978
rect 198298 165922 198368 165978
rect 198048 165888 198368 165922
rect 228768 166350 229088 166384
rect 228768 166294 228838 166350
rect 228894 166294 228962 166350
rect 229018 166294 229088 166350
rect 228768 166226 229088 166294
rect 228768 166170 228838 166226
rect 228894 166170 228962 166226
rect 229018 166170 229088 166226
rect 228768 166102 229088 166170
rect 228768 166046 228838 166102
rect 228894 166046 228962 166102
rect 229018 166046 229088 166102
rect 228768 165978 229088 166046
rect 228768 165922 228838 165978
rect 228894 165922 228962 165978
rect 229018 165922 229088 165978
rect 228768 165888 229088 165922
rect 259488 166350 259808 166384
rect 259488 166294 259558 166350
rect 259614 166294 259682 166350
rect 259738 166294 259808 166350
rect 259488 166226 259808 166294
rect 259488 166170 259558 166226
rect 259614 166170 259682 166226
rect 259738 166170 259808 166226
rect 259488 166102 259808 166170
rect 259488 166046 259558 166102
rect 259614 166046 259682 166102
rect 259738 166046 259808 166102
rect 259488 165978 259808 166046
rect 259488 165922 259558 165978
rect 259614 165922 259682 165978
rect 259738 165922 259808 165978
rect 259488 165888 259808 165922
rect 59808 154350 60128 154384
rect 59808 154294 59878 154350
rect 59934 154294 60002 154350
rect 60058 154294 60128 154350
rect 59808 154226 60128 154294
rect 59808 154170 59878 154226
rect 59934 154170 60002 154226
rect 60058 154170 60128 154226
rect 59808 154102 60128 154170
rect 59808 154046 59878 154102
rect 59934 154046 60002 154102
rect 60058 154046 60128 154102
rect 59808 153978 60128 154046
rect 59808 153922 59878 153978
rect 59934 153922 60002 153978
rect 60058 153922 60128 153978
rect 59808 153888 60128 153922
rect 90528 154350 90848 154384
rect 90528 154294 90598 154350
rect 90654 154294 90722 154350
rect 90778 154294 90848 154350
rect 90528 154226 90848 154294
rect 90528 154170 90598 154226
rect 90654 154170 90722 154226
rect 90778 154170 90848 154226
rect 90528 154102 90848 154170
rect 90528 154046 90598 154102
rect 90654 154046 90722 154102
rect 90778 154046 90848 154102
rect 90528 153978 90848 154046
rect 90528 153922 90598 153978
rect 90654 153922 90722 153978
rect 90778 153922 90848 153978
rect 90528 153888 90848 153922
rect 121248 154350 121568 154384
rect 121248 154294 121318 154350
rect 121374 154294 121442 154350
rect 121498 154294 121568 154350
rect 121248 154226 121568 154294
rect 121248 154170 121318 154226
rect 121374 154170 121442 154226
rect 121498 154170 121568 154226
rect 121248 154102 121568 154170
rect 121248 154046 121318 154102
rect 121374 154046 121442 154102
rect 121498 154046 121568 154102
rect 121248 153978 121568 154046
rect 121248 153922 121318 153978
rect 121374 153922 121442 153978
rect 121498 153922 121568 153978
rect 121248 153888 121568 153922
rect 151968 154350 152288 154384
rect 151968 154294 152038 154350
rect 152094 154294 152162 154350
rect 152218 154294 152288 154350
rect 151968 154226 152288 154294
rect 151968 154170 152038 154226
rect 152094 154170 152162 154226
rect 152218 154170 152288 154226
rect 151968 154102 152288 154170
rect 151968 154046 152038 154102
rect 152094 154046 152162 154102
rect 152218 154046 152288 154102
rect 151968 153978 152288 154046
rect 151968 153922 152038 153978
rect 152094 153922 152162 153978
rect 152218 153922 152288 153978
rect 151968 153888 152288 153922
rect 182688 154350 183008 154384
rect 182688 154294 182758 154350
rect 182814 154294 182882 154350
rect 182938 154294 183008 154350
rect 182688 154226 183008 154294
rect 182688 154170 182758 154226
rect 182814 154170 182882 154226
rect 182938 154170 183008 154226
rect 182688 154102 183008 154170
rect 182688 154046 182758 154102
rect 182814 154046 182882 154102
rect 182938 154046 183008 154102
rect 182688 153978 183008 154046
rect 182688 153922 182758 153978
rect 182814 153922 182882 153978
rect 182938 153922 183008 153978
rect 182688 153888 183008 153922
rect 213408 154350 213728 154384
rect 213408 154294 213478 154350
rect 213534 154294 213602 154350
rect 213658 154294 213728 154350
rect 213408 154226 213728 154294
rect 213408 154170 213478 154226
rect 213534 154170 213602 154226
rect 213658 154170 213728 154226
rect 213408 154102 213728 154170
rect 213408 154046 213478 154102
rect 213534 154046 213602 154102
rect 213658 154046 213728 154102
rect 213408 153978 213728 154046
rect 213408 153922 213478 153978
rect 213534 153922 213602 153978
rect 213658 153922 213728 153978
rect 213408 153888 213728 153922
rect 244128 154350 244448 154384
rect 244128 154294 244198 154350
rect 244254 154294 244322 154350
rect 244378 154294 244448 154350
rect 244128 154226 244448 154294
rect 244128 154170 244198 154226
rect 244254 154170 244322 154226
rect 244378 154170 244448 154226
rect 244128 154102 244448 154170
rect 244128 154046 244198 154102
rect 244254 154046 244322 154102
rect 244378 154046 244448 154102
rect 244128 153978 244448 154046
rect 244128 153922 244198 153978
rect 244254 153922 244322 153978
rect 244378 153922 244448 153978
rect 244128 153888 244448 153922
rect 75168 148350 75488 148384
rect 75168 148294 75238 148350
rect 75294 148294 75362 148350
rect 75418 148294 75488 148350
rect 75168 148226 75488 148294
rect 75168 148170 75238 148226
rect 75294 148170 75362 148226
rect 75418 148170 75488 148226
rect 75168 148102 75488 148170
rect 75168 148046 75238 148102
rect 75294 148046 75362 148102
rect 75418 148046 75488 148102
rect 75168 147978 75488 148046
rect 75168 147922 75238 147978
rect 75294 147922 75362 147978
rect 75418 147922 75488 147978
rect 75168 147888 75488 147922
rect 105888 148350 106208 148384
rect 105888 148294 105958 148350
rect 106014 148294 106082 148350
rect 106138 148294 106208 148350
rect 105888 148226 106208 148294
rect 105888 148170 105958 148226
rect 106014 148170 106082 148226
rect 106138 148170 106208 148226
rect 105888 148102 106208 148170
rect 105888 148046 105958 148102
rect 106014 148046 106082 148102
rect 106138 148046 106208 148102
rect 105888 147978 106208 148046
rect 105888 147922 105958 147978
rect 106014 147922 106082 147978
rect 106138 147922 106208 147978
rect 105888 147888 106208 147922
rect 136608 148350 136928 148384
rect 136608 148294 136678 148350
rect 136734 148294 136802 148350
rect 136858 148294 136928 148350
rect 136608 148226 136928 148294
rect 136608 148170 136678 148226
rect 136734 148170 136802 148226
rect 136858 148170 136928 148226
rect 136608 148102 136928 148170
rect 136608 148046 136678 148102
rect 136734 148046 136802 148102
rect 136858 148046 136928 148102
rect 136608 147978 136928 148046
rect 136608 147922 136678 147978
rect 136734 147922 136802 147978
rect 136858 147922 136928 147978
rect 136608 147888 136928 147922
rect 167328 148350 167648 148384
rect 167328 148294 167398 148350
rect 167454 148294 167522 148350
rect 167578 148294 167648 148350
rect 167328 148226 167648 148294
rect 167328 148170 167398 148226
rect 167454 148170 167522 148226
rect 167578 148170 167648 148226
rect 167328 148102 167648 148170
rect 167328 148046 167398 148102
rect 167454 148046 167522 148102
rect 167578 148046 167648 148102
rect 167328 147978 167648 148046
rect 167328 147922 167398 147978
rect 167454 147922 167522 147978
rect 167578 147922 167648 147978
rect 167328 147888 167648 147922
rect 198048 148350 198368 148384
rect 198048 148294 198118 148350
rect 198174 148294 198242 148350
rect 198298 148294 198368 148350
rect 198048 148226 198368 148294
rect 198048 148170 198118 148226
rect 198174 148170 198242 148226
rect 198298 148170 198368 148226
rect 198048 148102 198368 148170
rect 198048 148046 198118 148102
rect 198174 148046 198242 148102
rect 198298 148046 198368 148102
rect 198048 147978 198368 148046
rect 198048 147922 198118 147978
rect 198174 147922 198242 147978
rect 198298 147922 198368 147978
rect 198048 147888 198368 147922
rect 228768 148350 229088 148384
rect 228768 148294 228838 148350
rect 228894 148294 228962 148350
rect 229018 148294 229088 148350
rect 228768 148226 229088 148294
rect 228768 148170 228838 148226
rect 228894 148170 228962 148226
rect 229018 148170 229088 148226
rect 228768 148102 229088 148170
rect 228768 148046 228838 148102
rect 228894 148046 228962 148102
rect 229018 148046 229088 148102
rect 228768 147978 229088 148046
rect 228768 147922 228838 147978
rect 228894 147922 228962 147978
rect 229018 147922 229088 147978
rect 228768 147888 229088 147922
rect 259488 148350 259808 148384
rect 259488 148294 259558 148350
rect 259614 148294 259682 148350
rect 259738 148294 259808 148350
rect 259488 148226 259808 148294
rect 259488 148170 259558 148226
rect 259614 148170 259682 148226
rect 259738 148170 259808 148226
rect 259488 148102 259808 148170
rect 259488 148046 259558 148102
rect 259614 148046 259682 148102
rect 259738 148046 259808 148102
rect 259488 147978 259808 148046
rect 259488 147922 259558 147978
rect 259614 147922 259682 147978
rect 259738 147922 259808 147978
rect 259488 147888 259808 147922
rect 59808 136350 60128 136384
rect 59808 136294 59878 136350
rect 59934 136294 60002 136350
rect 60058 136294 60128 136350
rect 59808 136226 60128 136294
rect 59808 136170 59878 136226
rect 59934 136170 60002 136226
rect 60058 136170 60128 136226
rect 59808 136102 60128 136170
rect 59808 136046 59878 136102
rect 59934 136046 60002 136102
rect 60058 136046 60128 136102
rect 59808 135978 60128 136046
rect 59808 135922 59878 135978
rect 59934 135922 60002 135978
rect 60058 135922 60128 135978
rect 59808 135888 60128 135922
rect 90528 136350 90848 136384
rect 90528 136294 90598 136350
rect 90654 136294 90722 136350
rect 90778 136294 90848 136350
rect 90528 136226 90848 136294
rect 90528 136170 90598 136226
rect 90654 136170 90722 136226
rect 90778 136170 90848 136226
rect 90528 136102 90848 136170
rect 90528 136046 90598 136102
rect 90654 136046 90722 136102
rect 90778 136046 90848 136102
rect 90528 135978 90848 136046
rect 90528 135922 90598 135978
rect 90654 135922 90722 135978
rect 90778 135922 90848 135978
rect 90528 135888 90848 135922
rect 121248 136350 121568 136384
rect 121248 136294 121318 136350
rect 121374 136294 121442 136350
rect 121498 136294 121568 136350
rect 121248 136226 121568 136294
rect 121248 136170 121318 136226
rect 121374 136170 121442 136226
rect 121498 136170 121568 136226
rect 121248 136102 121568 136170
rect 121248 136046 121318 136102
rect 121374 136046 121442 136102
rect 121498 136046 121568 136102
rect 121248 135978 121568 136046
rect 121248 135922 121318 135978
rect 121374 135922 121442 135978
rect 121498 135922 121568 135978
rect 121248 135888 121568 135922
rect 151968 136350 152288 136384
rect 151968 136294 152038 136350
rect 152094 136294 152162 136350
rect 152218 136294 152288 136350
rect 151968 136226 152288 136294
rect 151968 136170 152038 136226
rect 152094 136170 152162 136226
rect 152218 136170 152288 136226
rect 151968 136102 152288 136170
rect 151968 136046 152038 136102
rect 152094 136046 152162 136102
rect 152218 136046 152288 136102
rect 151968 135978 152288 136046
rect 151968 135922 152038 135978
rect 152094 135922 152162 135978
rect 152218 135922 152288 135978
rect 151968 135888 152288 135922
rect 182688 136350 183008 136384
rect 182688 136294 182758 136350
rect 182814 136294 182882 136350
rect 182938 136294 183008 136350
rect 182688 136226 183008 136294
rect 182688 136170 182758 136226
rect 182814 136170 182882 136226
rect 182938 136170 183008 136226
rect 182688 136102 183008 136170
rect 182688 136046 182758 136102
rect 182814 136046 182882 136102
rect 182938 136046 183008 136102
rect 182688 135978 183008 136046
rect 182688 135922 182758 135978
rect 182814 135922 182882 135978
rect 182938 135922 183008 135978
rect 182688 135888 183008 135922
rect 213408 136350 213728 136384
rect 213408 136294 213478 136350
rect 213534 136294 213602 136350
rect 213658 136294 213728 136350
rect 213408 136226 213728 136294
rect 213408 136170 213478 136226
rect 213534 136170 213602 136226
rect 213658 136170 213728 136226
rect 213408 136102 213728 136170
rect 213408 136046 213478 136102
rect 213534 136046 213602 136102
rect 213658 136046 213728 136102
rect 213408 135978 213728 136046
rect 213408 135922 213478 135978
rect 213534 135922 213602 135978
rect 213658 135922 213728 135978
rect 213408 135888 213728 135922
rect 244128 136350 244448 136384
rect 244128 136294 244198 136350
rect 244254 136294 244322 136350
rect 244378 136294 244448 136350
rect 244128 136226 244448 136294
rect 244128 136170 244198 136226
rect 244254 136170 244322 136226
rect 244378 136170 244448 136226
rect 244128 136102 244448 136170
rect 244128 136046 244198 136102
rect 244254 136046 244322 136102
rect 244378 136046 244448 136102
rect 244128 135978 244448 136046
rect 244128 135922 244198 135978
rect 244254 135922 244322 135978
rect 244378 135922 244448 135978
rect 244128 135888 244448 135922
rect 75168 130350 75488 130384
rect 75168 130294 75238 130350
rect 75294 130294 75362 130350
rect 75418 130294 75488 130350
rect 75168 130226 75488 130294
rect 75168 130170 75238 130226
rect 75294 130170 75362 130226
rect 75418 130170 75488 130226
rect 75168 130102 75488 130170
rect 75168 130046 75238 130102
rect 75294 130046 75362 130102
rect 75418 130046 75488 130102
rect 75168 129978 75488 130046
rect 75168 129922 75238 129978
rect 75294 129922 75362 129978
rect 75418 129922 75488 129978
rect 75168 129888 75488 129922
rect 105888 130350 106208 130384
rect 105888 130294 105958 130350
rect 106014 130294 106082 130350
rect 106138 130294 106208 130350
rect 105888 130226 106208 130294
rect 105888 130170 105958 130226
rect 106014 130170 106082 130226
rect 106138 130170 106208 130226
rect 105888 130102 106208 130170
rect 105888 130046 105958 130102
rect 106014 130046 106082 130102
rect 106138 130046 106208 130102
rect 105888 129978 106208 130046
rect 105888 129922 105958 129978
rect 106014 129922 106082 129978
rect 106138 129922 106208 129978
rect 105888 129888 106208 129922
rect 136608 130350 136928 130384
rect 136608 130294 136678 130350
rect 136734 130294 136802 130350
rect 136858 130294 136928 130350
rect 136608 130226 136928 130294
rect 136608 130170 136678 130226
rect 136734 130170 136802 130226
rect 136858 130170 136928 130226
rect 136608 130102 136928 130170
rect 136608 130046 136678 130102
rect 136734 130046 136802 130102
rect 136858 130046 136928 130102
rect 136608 129978 136928 130046
rect 136608 129922 136678 129978
rect 136734 129922 136802 129978
rect 136858 129922 136928 129978
rect 136608 129888 136928 129922
rect 167328 130350 167648 130384
rect 167328 130294 167398 130350
rect 167454 130294 167522 130350
rect 167578 130294 167648 130350
rect 167328 130226 167648 130294
rect 167328 130170 167398 130226
rect 167454 130170 167522 130226
rect 167578 130170 167648 130226
rect 167328 130102 167648 130170
rect 167328 130046 167398 130102
rect 167454 130046 167522 130102
rect 167578 130046 167648 130102
rect 167328 129978 167648 130046
rect 167328 129922 167398 129978
rect 167454 129922 167522 129978
rect 167578 129922 167648 129978
rect 167328 129888 167648 129922
rect 198048 130350 198368 130384
rect 198048 130294 198118 130350
rect 198174 130294 198242 130350
rect 198298 130294 198368 130350
rect 198048 130226 198368 130294
rect 198048 130170 198118 130226
rect 198174 130170 198242 130226
rect 198298 130170 198368 130226
rect 198048 130102 198368 130170
rect 198048 130046 198118 130102
rect 198174 130046 198242 130102
rect 198298 130046 198368 130102
rect 198048 129978 198368 130046
rect 198048 129922 198118 129978
rect 198174 129922 198242 129978
rect 198298 129922 198368 129978
rect 198048 129888 198368 129922
rect 228768 130350 229088 130384
rect 228768 130294 228838 130350
rect 228894 130294 228962 130350
rect 229018 130294 229088 130350
rect 228768 130226 229088 130294
rect 228768 130170 228838 130226
rect 228894 130170 228962 130226
rect 229018 130170 229088 130226
rect 228768 130102 229088 130170
rect 228768 130046 228838 130102
rect 228894 130046 228962 130102
rect 229018 130046 229088 130102
rect 228768 129978 229088 130046
rect 228768 129922 228838 129978
rect 228894 129922 228962 129978
rect 229018 129922 229088 129978
rect 228768 129888 229088 129922
rect 259488 130350 259808 130384
rect 259488 130294 259558 130350
rect 259614 130294 259682 130350
rect 259738 130294 259808 130350
rect 259488 130226 259808 130294
rect 259488 130170 259558 130226
rect 259614 130170 259682 130226
rect 259738 130170 259808 130226
rect 259488 130102 259808 130170
rect 259488 130046 259558 130102
rect 259614 130046 259682 130102
rect 259738 130046 259808 130102
rect 259488 129978 259808 130046
rect 259488 129922 259558 129978
rect 259614 129922 259682 129978
rect 259738 129922 259808 129978
rect 259488 129888 259808 129922
rect 59808 118350 60128 118384
rect 59808 118294 59878 118350
rect 59934 118294 60002 118350
rect 60058 118294 60128 118350
rect 59808 118226 60128 118294
rect 59808 118170 59878 118226
rect 59934 118170 60002 118226
rect 60058 118170 60128 118226
rect 59808 118102 60128 118170
rect 59808 118046 59878 118102
rect 59934 118046 60002 118102
rect 60058 118046 60128 118102
rect 59808 117978 60128 118046
rect 59808 117922 59878 117978
rect 59934 117922 60002 117978
rect 60058 117922 60128 117978
rect 59808 117888 60128 117922
rect 90528 118350 90848 118384
rect 90528 118294 90598 118350
rect 90654 118294 90722 118350
rect 90778 118294 90848 118350
rect 90528 118226 90848 118294
rect 90528 118170 90598 118226
rect 90654 118170 90722 118226
rect 90778 118170 90848 118226
rect 90528 118102 90848 118170
rect 90528 118046 90598 118102
rect 90654 118046 90722 118102
rect 90778 118046 90848 118102
rect 90528 117978 90848 118046
rect 90528 117922 90598 117978
rect 90654 117922 90722 117978
rect 90778 117922 90848 117978
rect 90528 117888 90848 117922
rect 121248 118350 121568 118384
rect 121248 118294 121318 118350
rect 121374 118294 121442 118350
rect 121498 118294 121568 118350
rect 121248 118226 121568 118294
rect 121248 118170 121318 118226
rect 121374 118170 121442 118226
rect 121498 118170 121568 118226
rect 121248 118102 121568 118170
rect 121248 118046 121318 118102
rect 121374 118046 121442 118102
rect 121498 118046 121568 118102
rect 121248 117978 121568 118046
rect 121248 117922 121318 117978
rect 121374 117922 121442 117978
rect 121498 117922 121568 117978
rect 121248 117888 121568 117922
rect 151968 118350 152288 118384
rect 151968 118294 152038 118350
rect 152094 118294 152162 118350
rect 152218 118294 152288 118350
rect 151968 118226 152288 118294
rect 151968 118170 152038 118226
rect 152094 118170 152162 118226
rect 152218 118170 152288 118226
rect 151968 118102 152288 118170
rect 151968 118046 152038 118102
rect 152094 118046 152162 118102
rect 152218 118046 152288 118102
rect 151968 117978 152288 118046
rect 151968 117922 152038 117978
rect 152094 117922 152162 117978
rect 152218 117922 152288 117978
rect 151968 117888 152288 117922
rect 182688 118350 183008 118384
rect 182688 118294 182758 118350
rect 182814 118294 182882 118350
rect 182938 118294 183008 118350
rect 182688 118226 183008 118294
rect 182688 118170 182758 118226
rect 182814 118170 182882 118226
rect 182938 118170 183008 118226
rect 182688 118102 183008 118170
rect 182688 118046 182758 118102
rect 182814 118046 182882 118102
rect 182938 118046 183008 118102
rect 182688 117978 183008 118046
rect 182688 117922 182758 117978
rect 182814 117922 182882 117978
rect 182938 117922 183008 117978
rect 182688 117888 183008 117922
rect 213408 118350 213728 118384
rect 213408 118294 213478 118350
rect 213534 118294 213602 118350
rect 213658 118294 213728 118350
rect 213408 118226 213728 118294
rect 213408 118170 213478 118226
rect 213534 118170 213602 118226
rect 213658 118170 213728 118226
rect 213408 118102 213728 118170
rect 213408 118046 213478 118102
rect 213534 118046 213602 118102
rect 213658 118046 213728 118102
rect 213408 117978 213728 118046
rect 213408 117922 213478 117978
rect 213534 117922 213602 117978
rect 213658 117922 213728 117978
rect 213408 117888 213728 117922
rect 244128 118350 244448 118384
rect 244128 118294 244198 118350
rect 244254 118294 244322 118350
rect 244378 118294 244448 118350
rect 244128 118226 244448 118294
rect 244128 118170 244198 118226
rect 244254 118170 244322 118226
rect 244378 118170 244448 118226
rect 244128 118102 244448 118170
rect 244128 118046 244198 118102
rect 244254 118046 244322 118102
rect 244378 118046 244448 118102
rect 244128 117978 244448 118046
rect 244128 117922 244198 117978
rect 244254 117922 244322 117978
rect 244378 117922 244448 117978
rect 244128 117888 244448 117922
rect 75168 112350 75488 112384
rect 75168 112294 75238 112350
rect 75294 112294 75362 112350
rect 75418 112294 75488 112350
rect 75168 112226 75488 112294
rect 75168 112170 75238 112226
rect 75294 112170 75362 112226
rect 75418 112170 75488 112226
rect 75168 112102 75488 112170
rect 75168 112046 75238 112102
rect 75294 112046 75362 112102
rect 75418 112046 75488 112102
rect 75168 111978 75488 112046
rect 75168 111922 75238 111978
rect 75294 111922 75362 111978
rect 75418 111922 75488 111978
rect 75168 111888 75488 111922
rect 105888 112350 106208 112384
rect 105888 112294 105958 112350
rect 106014 112294 106082 112350
rect 106138 112294 106208 112350
rect 105888 112226 106208 112294
rect 105888 112170 105958 112226
rect 106014 112170 106082 112226
rect 106138 112170 106208 112226
rect 105888 112102 106208 112170
rect 105888 112046 105958 112102
rect 106014 112046 106082 112102
rect 106138 112046 106208 112102
rect 105888 111978 106208 112046
rect 105888 111922 105958 111978
rect 106014 111922 106082 111978
rect 106138 111922 106208 111978
rect 105888 111888 106208 111922
rect 136608 112350 136928 112384
rect 136608 112294 136678 112350
rect 136734 112294 136802 112350
rect 136858 112294 136928 112350
rect 136608 112226 136928 112294
rect 136608 112170 136678 112226
rect 136734 112170 136802 112226
rect 136858 112170 136928 112226
rect 136608 112102 136928 112170
rect 136608 112046 136678 112102
rect 136734 112046 136802 112102
rect 136858 112046 136928 112102
rect 136608 111978 136928 112046
rect 136608 111922 136678 111978
rect 136734 111922 136802 111978
rect 136858 111922 136928 111978
rect 136608 111888 136928 111922
rect 167328 112350 167648 112384
rect 167328 112294 167398 112350
rect 167454 112294 167522 112350
rect 167578 112294 167648 112350
rect 167328 112226 167648 112294
rect 167328 112170 167398 112226
rect 167454 112170 167522 112226
rect 167578 112170 167648 112226
rect 167328 112102 167648 112170
rect 167328 112046 167398 112102
rect 167454 112046 167522 112102
rect 167578 112046 167648 112102
rect 167328 111978 167648 112046
rect 167328 111922 167398 111978
rect 167454 111922 167522 111978
rect 167578 111922 167648 111978
rect 167328 111888 167648 111922
rect 198048 112350 198368 112384
rect 198048 112294 198118 112350
rect 198174 112294 198242 112350
rect 198298 112294 198368 112350
rect 198048 112226 198368 112294
rect 198048 112170 198118 112226
rect 198174 112170 198242 112226
rect 198298 112170 198368 112226
rect 198048 112102 198368 112170
rect 198048 112046 198118 112102
rect 198174 112046 198242 112102
rect 198298 112046 198368 112102
rect 198048 111978 198368 112046
rect 198048 111922 198118 111978
rect 198174 111922 198242 111978
rect 198298 111922 198368 111978
rect 198048 111888 198368 111922
rect 228768 112350 229088 112384
rect 228768 112294 228838 112350
rect 228894 112294 228962 112350
rect 229018 112294 229088 112350
rect 228768 112226 229088 112294
rect 228768 112170 228838 112226
rect 228894 112170 228962 112226
rect 229018 112170 229088 112226
rect 228768 112102 229088 112170
rect 228768 112046 228838 112102
rect 228894 112046 228962 112102
rect 229018 112046 229088 112102
rect 228768 111978 229088 112046
rect 228768 111922 228838 111978
rect 228894 111922 228962 111978
rect 229018 111922 229088 111978
rect 228768 111888 229088 111922
rect 259488 112350 259808 112384
rect 259488 112294 259558 112350
rect 259614 112294 259682 112350
rect 259738 112294 259808 112350
rect 259488 112226 259808 112294
rect 259488 112170 259558 112226
rect 259614 112170 259682 112226
rect 259738 112170 259808 112226
rect 259488 112102 259808 112170
rect 259488 112046 259558 112102
rect 259614 112046 259682 112102
rect 259738 112046 259808 112102
rect 259488 111978 259808 112046
rect 259488 111922 259558 111978
rect 259614 111922 259682 111978
rect 259738 111922 259808 111978
rect 259488 111888 259808 111922
rect 59808 100350 60128 100384
rect 59808 100294 59878 100350
rect 59934 100294 60002 100350
rect 60058 100294 60128 100350
rect 59808 100226 60128 100294
rect 59808 100170 59878 100226
rect 59934 100170 60002 100226
rect 60058 100170 60128 100226
rect 59808 100102 60128 100170
rect 59808 100046 59878 100102
rect 59934 100046 60002 100102
rect 60058 100046 60128 100102
rect 59808 99978 60128 100046
rect 59808 99922 59878 99978
rect 59934 99922 60002 99978
rect 60058 99922 60128 99978
rect 59808 99888 60128 99922
rect 90528 100350 90848 100384
rect 90528 100294 90598 100350
rect 90654 100294 90722 100350
rect 90778 100294 90848 100350
rect 90528 100226 90848 100294
rect 90528 100170 90598 100226
rect 90654 100170 90722 100226
rect 90778 100170 90848 100226
rect 90528 100102 90848 100170
rect 90528 100046 90598 100102
rect 90654 100046 90722 100102
rect 90778 100046 90848 100102
rect 90528 99978 90848 100046
rect 90528 99922 90598 99978
rect 90654 99922 90722 99978
rect 90778 99922 90848 99978
rect 90528 99888 90848 99922
rect 121248 100350 121568 100384
rect 121248 100294 121318 100350
rect 121374 100294 121442 100350
rect 121498 100294 121568 100350
rect 121248 100226 121568 100294
rect 121248 100170 121318 100226
rect 121374 100170 121442 100226
rect 121498 100170 121568 100226
rect 121248 100102 121568 100170
rect 121248 100046 121318 100102
rect 121374 100046 121442 100102
rect 121498 100046 121568 100102
rect 121248 99978 121568 100046
rect 121248 99922 121318 99978
rect 121374 99922 121442 99978
rect 121498 99922 121568 99978
rect 121248 99888 121568 99922
rect 151968 100350 152288 100384
rect 151968 100294 152038 100350
rect 152094 100294 152162 100350
rect 152218 100294 152288 100350
rect 151968 100226 152288 100294
rect 151968 100170 152038 100226
rect 152094 100170 152162 100226
rect 152218 100170 152288 100226
rect 151968 100102 152288 100170
rect 151968 100046 152038 100102
rect 152094 100046 152162 100102
rect 152218 100046 152288 100102
rect 151968 99978 152288 100046
rect 151968 99922 152038 99978
rect 152094 99922 152162 99978
rect 152218 99922 152288 99978
rect 151968 99888 152288 99922
rect 182688 100350 183008 100384
rect 182688 100294 182758 100350
rect 182814 100294 182882 100350
rect 182938 100294 183008 100350
rect 182688 100226 183008 100294
rect 182688 100170 182758 100226
rect 182814 100170 182882 100226
rect 182938 100170 183008 100226
rect 182688 100102 183008 100170
rect 182688 100046 182758 100102
rect 182814 100046 182882 100102
rect 182938 100046 183008 100102
rect 182688 99978 183008 100046
rect 182688 99922 182758 99978
rect 182814 99922 182882 99978
rect 182938 99922 183008 99978
rect 182688 99888 183008 99922
rect 213408 100350 213728 100384
rect 213408 100294 213478 100350
rect 213534 100294 213602 100350
rect 213658 100294 213728 100350
rect 213408 100226 213728 100294
rect 213408 100170 213478 100226
rect 213534 100170 213602 100226
rect 213658 100170 213728 100226
rect 213408 100102 213728 100170
rect 213408 100046 213478 100102
rect 213534 100046 213602 100102
rect 213658 100046 213728 100102
rect 213408 99978 213728 100046
rect 213408 99922 213478 99978
rect 213534 99922 213602 99978
rect 213658 99922 213728 99978
rect 213408 99888 213728 99922
rect 244128 100350 244448 100384
rect 244128 100294 244198 100350
rect 244254 100294 244322 100350
rect 244378 100294 244448 100350
rect 244128 100226 244448 100294
rect 244128 100170 244198 100226
rect 244254 100170 244322 100226
rect 244378 100170 244448 100226
rect 244128 100102 244448 100170
rect 244128 100046 244198 100102
rect 244254 100046 244322 100102
rect 244378 100046 244448 100102
rect 244128 99978 244448 100046
rect 244128 99922 244198 99978
rect 244254 99922 244322 99978
rect 244378 99922 244448 99978
rect 244128 99888 244448 99922
rect 75168 94350 75488 94384
rect 75168 94294 75238 94350
rect 75294 94294 75362 94350
rect 75418 94294 75488 94350
rect 75168 94226 75488 94294
rect 75168 94170 75238 94226
rect 75294 94170 75362 94226
rect 75418 94170 75488 94226
rect 75168 94102 75488 94170
rect 75168 94046 75238 94102
rect 75294 94046 75362 94102
rect 75418 94046 75488 94102
rect 75168 93978 75488 94046
rect 75168 93922 75238 93978
rect 75294 93922 75362 93978
rect 75418 93922 75488 93978
rect 75168 93888 75488 93922
rect 105888 94350 106208 94384
rect 105888 94294 105958 94350
rect 106014 94294 106082 94350
rect 106138 94294 106208 94350
rect 105888 94226 106208 94294
rect 105888 94170 105958 94226
rect 106014 94170 106082 94226
rect 106138 94170 106208 94226
rect 105888 94102 106208 94170
rect 105888 94046 105958 94102
rect 106014 94046 106082 94102
rect 106138 94046 106208 94102
rect 105888 93978 106208 94046
rect 105888 93922 105958 93978
rect 106014 93922 106082 93978
rect 106138 93922 106208 93978
rect 105888 93888 106208 93922
rect 136608 94350 136928 94384
rect 136608 94294 136678 94350
rect 136734 94294 136802 94350
rect 136858 94294 136928 94350
rect 136608 94226 136928 94294
rect 136608 94170 136678 94226
rect 136734 94170 136802 94226
rect 136858 94170 136928 94226
rect 136608 94102 136928 94170
rect 136608 94046 136678 94102
rect 136734 94046 136802 94102
rect 136858 94046 136928 94102
rect 136608 93978 136928 94046
rect 136608 93922 136678 93978
rect 136734 93922 136802 93978
rect 136858 93922 136928 93978
rect 136608 93888 136928 93922
rect 167328 94350 167648 94384
rect 167328 94294 167398 94350
rect 167454 94294 167522 94350
rect 167578 94294 167648 94350
rect 167328 94226 167648 94294
rect 167328 94170 167398 94226
rect 167454 94170 167522 94226
rect 167578 94170 167648 94226
rect 167328 94102 167648 94170
rect 167328 94046 167398 94102
rect 167454 94046 167522 94102
rect 167578 94046 167648 94102
rect 167328 93978 167648 94046
rect 167328 93922 167398 93978
rect 167454 93922 167522 93978
rect 167578 93922 167648 93978
rect 167328 93888 167648 93922
rect 198048 94350 198368 94384
rect 198048 94294 198118 94350
rect 198174 94294 198242 94350
rect 198298 94294 198368 94350
rect 198048 94226 198368 94294
rect 198048 94170 198118 94226
rect 198174 94170 198242 94226
rect 198298 94170 198368 94226
rect 198048 94102 198368 94170
rect 198048 94046 198118 94102
rect 198174 94046 198242 94102
rect 198298 94046 198368 94102
rect 198048 93978 198368 94046
rect 198048 93922 198118 93978
rect 198174 93922 198242 93978
rect 198298 93922 198368 93978
rect 198048 93888 198368 93922
rect 228768 94350 229088 94384
rect 228768 94294 228838 94350
rect 228894 94294 228962 94350
rect 229018 94294 229088 94350
rect 228768 94226 229088 94294
rect 228768 94170 228838 94226
rect 228894 94170 228962 94226
rect 229018 94170 229088 94226
rect 228768 94102 229088 94170
rect 228768 94046 228838 94102
rect 228894 94046 228962 94102
rect 229018 94046 229088 94102
rect 228768 93978 229088 94046
rect 228768 93922 228838 93978
rect 228894 93922 228962 93978
rect 229018 93922 229088 93978
rect 228768 93888 229088 93922
rect 259488 94350 259808 94384
rect 259488 94294 259558 94350
rect 259614 94294 259682 94350
rect 259738 94294 259808 94350
rect 259488 94226 259808 94294
rect 259488 94170 259558 94226
rect 259614 94170 259682 94226
rect 259738 94170 259808 94226
rect 259488 94102 259808 94170
rect 259488 94046 259558 94102
rect 259614 94046 259682 94102
rect 259738 94046 259808 94102
rect 259488 93978 259808 94046
rect 259488 93922 259558 93978
rect 259614 93922 259682 93978
rect 259738 93922 259808 93978
rect 259488 93888 259808 93922
rect 59808 82350 60128 82384
rect 59808 82294 59878 82350
rect 59934 82294 60002 82350
rect 60058 82294 60128 82350
rect 59808 82226 60128 82294
rect 59808 82170 59878 82226
rect 59934 82170 60002 82226
rect 60058 82170 60128 82226
rect 59808 82102 60128 82170
rect 59808 82046 59878 82102
rect 59934 82046 60002 82102
rect 60058 82046 60128 82102
rect 59808 81978 60128 82046
rect 59808 81922 59878 81978
rect 59934 81922 60002 81978
rect 60058 81922 60128 81978
rect 59808 81888 60128 81922
rect 90528 82350 90848 82384
rect 90528 82294 90598 82350
rect 90654 82294 90722 82350
rect 90778 82294 90848 82350
rect 90528 82226 90848 82294
rect 90528 82170 90598 82226
rect 90654 82170 90722 82226
rect 90778 82170 90848 82226
rect 90528 82102 90848 82170
rect 90528 82046 90598 82102
rect 90654 82046 90722 82102
rect 90778 82046 90848 82102
rect 90528 81978 90848 82046
rect 90528 81922 90598 81978
rect 90654 81922 90722 81978
rect 90778 81922 90848 81978
rect 90528 81888 90848 81922
rect 121248 82350 121568 82384
rect 121248 82294 121318 82350
rect 121374 82294 121442 82350
rect 121498 82294 121568 82350
rect 121248 82226 121568 82294
rect 121248 82170 121318 82226
rect 121374 82170 121442 82226
rect 121498 82170 121568 82226
rect 121248 82102 121568 82170
rect 121248 82046 121318 82102
rect 121374 82046 121442 82102
rect 121498 82046 121568 82102
rect 121248 81978 121568 82046
rect 121248 81922 121318 81978
rect 121374 81922 121442 81978
rect 121498 81922 121568 81978
rect 121248 81888 121568 81922
rect 151968 82350 152288 82384
rect 151968 82294 152038 82350
rect 152094 82294 152162 82350
rect 152218 82294 152288 82350
rect 151968 82226 152288 82294
rect 151968 82170 152038 82226
rect 152094 82170 152162 82226
rect 152218 82170 152288 82226
rect 151968 82102 152288 82170
rect 151968 82046 152038 82102
rect 152094 82046 152162 82102
rect 152218 82046 152288 82102
rect 151968 81978 152288 82046
rect 151968 81922 152038 81978
rect 152094 81922 152162 81978
rect 152218 81922 152288 81978
rect 151968 81888 152288 81922
rect 182688 82350 183008 82384
rect 182688 82294 182758 82350
rect 182814 82294 182882 82350
rect 182938 82294 183008 82350
rect 182688 82226 183008 82294
rect 182688 82170 182758 82226
rect 182814 82170 182882 82226
rect 182938 82170 183008 82226
rect 182688 82102 183008 82170
rect 182688 82046 182758 82102
rect 182814 82046 182882 82102
rect 182938 82046 183008 82102
rect 182688 81978 183008 82046
rect 182688 81922 182758 81978
rect 182814 81922 182882 81978
rect 182938 81922 183008 81978
rect 182688 81888 183008 81922
rect 213408 82350 213728 82384
rect 213408 82294 213478 82350
rect 213534 82294 213602 82350
rect 213658 82294 213728 82350
rect 213408 82226 213728 82294
rect 213408 82170 213478 82226
rect 213534 82170 213602 82226
rect 213658 82170 213728 82226
rect 213408 82102 213728 82170
rect 213408 82046 213478 82102
rect 213534 82046 213602 82102
rect 213658 82046 213728 82102
rect 213408 81978 213728 82046
rect 213408 81922 213478 81978
rect 213534 81922 213602 81978
rect 213658 81922 213728 81978
rect 213408 81888 213728 81922
rect 244128 82350 244448 82384
rect 244128 82294 244198 82350
rect 244254 82294 244322 82350
rect 244378 82294 244448 82350
rect 244128 82226 244448 82294
rect 244128 82170 244198 82226
rect 244254 82170 244322 82226
rect 244378 82170 244448 82226
rect 244128 82102 244448 82170
rect 244128 82046 244198 82102
rect 244254 82046 244322 82102
rect 244378 82046 244448 82102
rect 244128 81978 244448 82046
rect 244128 81922 244198 81978
rect 244254 81922 244322 81978
rect 244378 81922 244448 81978
rect 244128 81888 244448 81922
rect 75168 76350 75488 76384
rect 75168 76294 75238 76350
rect 75294 76294 75362 76350
rect 75418 76294 75488 76350
rect 75168 76226 75488 76294
rect 75168 76170 75238 76226
rect 75294 76170 75362 76226
rect 75418 76170 75488 76226
rect 75168 76102 75488 76170
rect 75168 76046 75238 76102
rect 75294 76046 75362 76102
rect 75418 76046 75488 76102
rect 75168 75978 75488 76046
rect 75168 75922 75238 75978
rect 75294 75922 75362 75978
rect 75418 75922 75488 75978
rect 75168 75888 75488 75922
rect 105888 76350 106208 76384
rect 105888 76294 105958 76350
rect 106014 76294 106082 76350
rect 106138 76294 106208 76350
rect 105888 76226 106208 76294
rect 105888 76170 105958 76226
rect 106014 76170 106082 76226
rect 106138 76170 106208 76226
rect 105888 76102 106208 76170
rect 105888 76046 105958 76102
rect 106014 76046 106082 76102
rect 106138 76046 106208 76102
rect 105888 75978 106208 76046
rect 105888 75922 105958 75978
rect 106014 75922 106082 75978
rect 106138 75922 106208 75978
rect 105888 75888 106208 75922
rect 136608 76350 136928 76384
rect 136608 76294 136678 76350
rect 136734 76294 136802 76350
rect 136858 76294 136928 76350
rect 136608 76226 136928 76294
rect 136608 76170 136678 76226
rect 136734 76170 136802 76226
rect 136858 76170 136928 76226
rect 136608 76102 136928 76170
rect 136608 76046 136678 76102
rect 136734 76046 136802 76102
rect 136858 76046 136928 76102
rect 136608 75978 136928 76046
rect 136608 75922 136678 75978
rect 136734 75922 136802 75978
rect 136858 75922 136928 75978
rect 136608 75888 136928 75922
rect 167328 76350 167648 76384
rect 167328 76294 167398 76350
rect 167454 76294 167522 76350
rect 167578 76294 167648 76350
rect 167328 76226 167648 76294
rect 167328 76170 167398 76226
rect 167454 76170 167522 76226
rect 167578 76170 167648 76226
rect 167328 76102 167648 76170
rect 167328 76046 167398 76102
rect 167454 76046 167522 76102
rect 167578 76046 167648 76102
rect 167328 75978 167648 76046
rect 167328 75922 167398 75978
rect 167454 75922 167522 75978
rect 167578 75922 167648 75978
rect 167328 75888 167648 75922
rect 198048 76350 198368 76384
rect 198048 76294 198118 76350
rect 198174 76294 198242 76350
rect 198298 76294 198368 76350
rect 198048 76226 198368 76294
rect 198048 76170 198118 76226
rect 198174 76170 198242 76226
rect 198298 76170 198368 76226
rect 198048 76102 198368 76170
rect 198048 76046 198118 76102
rect 198174 76046 198242 76102
rect 198298 76046 198368 76102
rect 198048 75978 198368 76046
rect 198048 75922 198118 75978
rect 198174 75922 198242 75978
rect 198298 75922 198368 75978
rect 198048 75888 198368 75922
rect 228768 76350 229088 76384
rect 228768 76294 228838 76350
rect 228894 76294 228962 76350
rect 229018 76294 229088 76350
rect 228768 76226 229088 76294
rect 228768 76170 228838 76226
rect 228894 76170 228962 76226
rect 229018 76170 229088 76226
rect 228768 76102 229088 76170
rect 228768 76046 228838 76102
rect 228894 76046 228962 76102
rect 229018 76046 229088 76102
rect 228768 75978 229088 76046
rect 228768 75922 228838 75978
rect 228894 75922 228962 75978
rect 229018 75922 229088 75978
rect 228768 75888 229088 75922
rect 259488 76350 259808 76384
rect 259488 76294 259558 76350
rect 259614 76294 259682 76350
rect 259738 76294 259808 76350
rect 259488 76226 259808 76294
rect 259488 76170 259558 76226
rect 259614 76170 259682 76226
rect 259738 76170 259808 76226
rect 259488 76102 259808 76170
rect 259488 76046 259558 76102
rect 259614 76046 259682 76102
rect 259738 76046 259808 76102
rect 259488 75978 259808 76046
rect 259488 75922 259558 75978
rect 259614 75922 259682 75978
rect 259738 75922 259808 75978
rect 259488 75888 259808 75922
rect 59808 64350 60128 64384
rect 59808 64294 59878 64350
rect 59934 64294 60002 64350
rect 60058 64294 60128 64350
rect 59808 64226 60128 64294
rect 59808 64170 59878 64226
rect 59934 64170 60002 64226
rect 60058 64170 60128 64226
rect 59808 64102 60128 64170
rect 59808 64046 59878 64102
rect 59934 64046 60002 64102
rect 60058 64046 60128 64102
rect 59808 63978 60128 64046
rect 59808 63922 59878 63978
rect 59934 63922 60002 63978
rect 60058 63922 60128 63978
rect 59808 63888 60128 63922
rect 90528 64350 90848 64384
rect 90528 64294 90598 64350
rect 90654 64294 90722 64350
rect 90778 64294 90848 64350
rect 90528 64226 90848 64294
rect 90528 64170 90598 64226
rect 90654 64170 90722 64226
rect 90778 64170 90848 64226
rect 90528 64102 90848 64170
rect 90528 64046 90598 64102
rect 90654 64046 90722 64102
rect 90778 64046 90848 64102
rect 90528 63978 90848 64046
rect 90528 63922 90598 63978
rect 90654 63922 90722 63978
rect 90778 63922 90848 63978
rect 90528 63888 90848 63922
rect 121248 64350 121568 64384
rect 121248 64294 121318 64350
rect 121374 64294 121442 64350
rect 121498 64294 121568 64350
rect 121248 64226 121568 64294
rect 121248 64170 121318 64226
rect 121374 64170 121442 64226
rect 121498 64170 121568 64226
rect 121248 64102 121568 64170
rect 121248 64046 121318 64102
rect 121374 64046 121442 64102
rect 121498 64046 121568 64102
rect 121248 63978 121568 64046
rect 121248 63922 121318 63978
rect 121374 63922 121442 63978
rect 121498 63922 121568 63978
rect 121248 63888 121568 63922
rect 151968 64350 152288 64384
rect 151968 64294 152038 64350
rect 152094 64294 152162 64350
rect 152218 64294 152288 64350
rect 151968 64226 152288 64294
rect 151968 64170 152038 64226
rect 152094 64170 152162 64226
rect 152218 64170 152288 64226
rect 151968 64102 152288 64170
rect 151968 64046 152038 64102
rect 152094 64046 152162 64102
rect 152218 64046 152288 64102
rect 151968 63978 152288 64046
rect 151968 63922 152038 63978
rect 152094 63922 152162 63978
rect 152218 63922 152288 63978
rect 151968 63888 152288 63922
rect 182688 64350 183008 64384
rect 182688 64294 182758 64350
rect 182814 64294 182882 64350
rect 182938 64294 183008 64350
rect 182688 64226 183008 64294
rect 182688 64170 182758 64226
rect 182814 64170 182882 64226
rect 182938 64170 183008 64226
rect 182688 64102 183008 64170
rect 182688 64046 182758 64102
rect 182814 64046 182882 64102
rect 182938 64046 183008 64102
rect 182688 63978 183008 64046
rect 182688 63922 182758 63978
rect 182814 63922 182882 63978
rect 182938 63922 183008 63978
rect 182688 63888 183008 63922
rect 213408 64350 213728 64384
rect 213408 64294 213478 64350
rect 213534 64294 213602 64350
rect 213658 64294 213728 64350
rect 213408 64226 213728 64294
rect 213408 64170 213478 64226
rect 213534 64170 213602 64226
rect 213658 64170 213728 64226
rect 213408 64102 213728 64170
rect 213408 64046 213478 64102
rect 213534 64046 213602 64102
rect 213658 64046 213728 64102
rect 213408 63978 213728 64046
rect 213408 63922 213478 63978
rect 213534 63922 213602 63978
rect 213658 63922 213728 63978
rect 213408 63888 213728 63922
rect 244128 64350 244448 64384
rect 244128 64294 244198 64350
rect 244254 64294 244322 64350
rect 244378 64294 244448 64350
rect 244128 64226 244448 64294
rect 244128 64170 244198 64226
rect 244254 64170 244322 64226
rect 244378 64170 244448 64226
rect 244128 64102 244448 64170
rect 244128 64046 244198 64102
rect 244254 64046 244322 64102
rect 244378 64046 244448 64102
rect 244128 63978 244448 64046
rect 244128 63922 244198 63978
rect 244254 63922 244322 63978
rect 244378 63922 244448 63978
rect 244128 63888 244448 63922
rect 75168 58350 75488 58384
rect 75168 58294 75238 58350
rect 75294 58294 75362 58350
rect 75418 58294 75488 58350
rect 75168 58226 75488 58294
rect 75168 58170 75238 58226
rect 75294 58170 75362 58226
rect 75418 58170 75488 58226
rect 75168 58102 75488 58170
rect 75168 58046 75238 58102
rect 75294 58046 75362 58102
rect 75418 58046 75488 58102
rect 75168 57978 75488 58046
rect 75168 57922 75238 57978
rect 75294 57922 75362 57978
rect 75418 57922 75488 57978
rect 75168 57888 75488 57922
rect 105888 58350 106208 58384
rect 105888 58294 105958 58350
rect 106014 58294 106082 58350
rect 106138 58294 106208 58350
rect 105888 58226 106208 58294
rect 105888 58170 105958 58226
rect 106014 58170 106082 58226
rect 106138 58170 106208 58226
rect 105888 58102 106208 58170
rect 105888 58046 105958 58102
rect 106014 58046 106082 58102
rect 106138 58046 106208 58102
rect 105888 57978 106208 58046
rect 105888 57922 105958 57978
rect 106014 57922 106082 57978
rect 106138 57922 106208 57978
rect 105888 57888 106208 57922
rect 136608 58350 136928 58384
rect 136608 58294 136678 58350
rect 136734 58294 136802 58350
rect 136858 58294 136928 58350
rect 136608 58226 136928 58294
rect 136608 58170 136678 58226
rect 136734 58170 136802 58226
rect 136858 58170 136928 58226
rect 136608 58102 136928 58170
rect 136608 58046 136678 58102
rect 136734 58046 136802 58102
rect 136858 58046 136928 58102
rect 136608 57978 136928 58046
rect 136608 57922 136678 57978
rect 136734 57922 136802 57978
rect 136858 57922 136928 57978
rect 136608 57888 136928 57922
rect 167328 58350 167648 58384
rect 167328 58294 167398 58350
rect 167454 58294 167522 58350
rect 167578 58294 167648 58350
rect 167328 58226 167648 58294
rect 167328 58170 167398 58226
rect 167454 58170 167522 58226
rect 167578 58170 167648 58226
rect 167328 58102 167648 58170
rect 167328 58046 167398 58102
rect 167454 58046 167522 58102
rect 167578 58046 167648 58102
rect 167328 57978 167648 58046
rect 167328 57922 167398 57978
rect 167454 57922 167522 57978
rect 167578 57922 167648 57978
rect 167328 57888 167648 57922
rect 198048 58350 198368 58384
rect 198048 58294 198118 58350
rect 198174 58294 198242 58350
rect 198298 58294 198368 58350
rect 198048 58226 198368 58294
rect 198048 58170 198118 58226
rect 198174 58170 198242 58226
rect 198298 58170 198368 58226
rect 198048 58102 198368 58170
rect 198048 58046 198118 58102
rect 198174 58046 198242 58102
rect 198298 58046 198368 58102
rect 198048 57978 198368 58046
rect 198048 57922 198118 57978
rect 198174 57922 198242 57978
rect 198298 57922 198368 57978
rect 198048 57888 198368 57922
rect 228768 58350 229088 58384
rect 228768 58294 228838 58350
rect 228894 58294 228962 58350
rect 229018 58294 229088 58350
rect 228768 58226 229088 58294
rect 228768 58170 228838 58226
rect 228894 58170 228962 58226
rect 229018 58170 229088 58226
rect 228768 58102 229088 58170
rect 228768 58046 228838 58102
rect 228894 58046 228962 58102
rect 229018 58046 229088 58102
rect 228768 57978 229088 58046
rect 228768 57922 228838 57978
rect 228894 57922 228962 57978
rect 229018 57922 229088 57978
rect 228768 57888 229088 57922
rect 259488 58350 259808 58384
rect 259488 58294 259558 58350
rect 259614 58294 259682 58350
rect 259738 58294 259808 58350
rect 259488 58226 259808 58294
rect 259488 58170 259558 58226
rect 259614 58170 259682 58226
rect 259738 58170 259808 58226
rect 259488 58102 259808 58170
rect 259488 58046 259558 58102
rect 259614 58046 259682 58102
rect 259738 58046 259808 58102
rect 259488 57978 259808 58046
rect 259488 57922 259558 57978
rect 259614 57922 259682 57978
rect 259738 57922 259808 57978
rect 259488 57888 259808 57922
rect 51996 4498 52052 4508
rect 66858 40350 67478 48802
rect 66858 40294 66954 40350
rect 67010 40294 67078 40350
rect 67134 40294 67202 40350
rect 67258 40294 67326 40350
rect 67382 40294 67478 40350
rect 66858 40226 67478 40294
rect 66858 40170 66954 40226
rect 67010 40170 67078 40226
rect 67134 40170 67202 40226
rect 67258 40170 67326 40226
rect 67382 40170 67478 40226
rect 66858 40102 67478 40170
rect 66858 40046 66954 40102
rect 67010 40046 67078 40102
rect 67134 40046 67202 40102
rect 67258 40046 67326 40102
rect 67382 40046 67478 40102
rect 66858 39978 67478 40046
rect 66858 39922 66954 39978
rect 67010 39922 67078 39978
rect 67134 39922 67202 39978
rect 67258 39922 67326 39978
rect 67382 39922 67478 39978
rect 66858 22350 67478 39922
rect 66858 22294 66954 22350
rect 67010 22294 67078 22350
rect 67134 22294 67202 22350
rect 67258 22294 67326 22350
rect 67382 22294 67478 22350
rect 66858 22226 67478 22294
rect 66858 22170 66954 22226
rect 67010 22170 67078 22226
rect 67134 22170 67202 22226
rect 67258 22170 67326 22226
rect 67382 22170 67478 22226
rect 66858 22102 67478 22170
rect 66858 22046 66954 22102
rect 67010 22046 67078 22102
rect 67134 22046 67202 22102
rect 67258 22046 67326 22102
rect 67382 22046 67478 22102
rect 66858 21978 67478 22046
rect 66858 21922 66954 21978
rect 67010 21922 67078 21978
rect 67134 21922 67202 21978
rect 67258 21922 67326 21978
rect 67382 21922 67478 21978
rect 51884 4386 51940 4396
rect 39858 -1176 39954 -1120
rect 40010 -1176 40078 -1120
rect 40134 -1176 40202 -1120
rect 40258 -1176 40326 -1120
rect 40382 -1176 40478 -1120
rect 39858 -1244 40478 -1176
rect 39858 -1300 39954 -1244
rect 40010 -1300 40078 -1244
rect 40134 -1300 40202 -1244
rect 40258 -1300 40326 -1244
rect 40382 -1300 40478 -1244
rect 39858 -1368 40478 -1300
rect 39858 -1424 39954 -1368
rect 40010 -1424 40078 -1368
rect 40134 -1424 40202 -1368
rect 40258 -1424 40326 -1368
rect 40382 -1424 40478 -1368
rect 39858 -1492 40478 -1424
rect 39858 -1548 39954 -1492
rect 40010 -1548 40078 -1492
rect 40134 -1548 40202 -1492
rect 40258 -1548 40326 -1492
rect 40382 -1548 40478 -1492
rect 39858 -1644 40478 -1548
rect 66858 4350 67478 21922
rect 66858 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 67478 4350
rect 66858 4226 67478 4294
rect 66858 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 67478 4226
rect 66858 4102 67478 4170
rect 66858 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 67478 4102
rect 66858 3978 67478 4046
rect 66858 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 67478 3978
rect 66858 -160 67478 3922
rect 66858 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 67478 -160
rect 66858 -284 67478 -216
rect 66858 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 67478 -284
rect 66858 -408 67478 -340
rect 66858 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 67478 -408
rect 66858 -532 67478 -464
rect 66858 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 67478 -532
rect 66858 -1644 67478 -588
rect 70578 46350 71198 48802
rect 70578 46294 70674 46350
rect 70730 46294 70798 46350
rect 70854 46294 70922 46350
rect 70978 46294 71046 46350
rect 71102 46294 71198 46350
rect 70578 46226 71198 46294
rect 70578 46170 70674 46226
rect 70730 46170 70798 46226
rect 70854 46170 70922 46226
rect 70978 46170 71046 46226
rect 71102 46170 71198 46226
rect 70578 46102 71198 46170
rect 70578 46046 70674 46102
rect 70730 46046 70798 46102
rect 70854 46046 70922 46102
rect 70978 46046 71046 46102
rect 71102 46046 71198 46102
rect 70578 45978 71198 46046
rect 70578 45922 70674 45978
rect 70730 45922 70798 45978
rect 70854 45922 70922 45978
rect 70978 45922 71046 45978
rect 71102 45922 71198 45978
rect 70578 28350 71198 45922
rect 70578 28294 70674 28350
rect 70730 28294 70798 28350
rect 70854 28294 70922 28350
rect 70978 28294 71046 28350
rect 71102 28294 71198 28350
rect 70578 28226 71198 28294
rect 70578 28170 70674 28226
rect 70730 28170 70798 28226
rect 70854 28170 70922 28226
rect 70978 28170 71046 28226
rect 71102 28170 71198 28226
rect 70578 28102 71198 28170
rect 70578 28046 70674 28102
rect 70730 28046 70798 28102
rect 70854 28046 70922 28102
rect 70978 28046 71046 28102
rect 71102 28046 71198 28102
rect 70578 27978 71198 28046
rect 70578 27922 70674 27978
rect 70730 27922 70798 27978
rect 70854 27922 70922 27978
rect 70978 27922 71046 27978
rect 71102 27922 71198 27978
rect 70578 10350 71198 27922
rect 70578 10294 70674 10350
rect 70730 10294 70798 10350
rect 70854 10294 70922 10350
rect 70978 10294 71046 10350
rect 71102 10294 71198 10350
rect 70578 10226 71198 10294
rect 70578 10170 70674 10226
rect 70730 10170 70798 10226
rect 70854 10170 70922 10226
rect 70978 10170 71046 10226
rect 71102 10170 71198 10226
rect 70578 10102 71198 10170
rect 70578 10046 70674 10102
rect 70730 10046 70798 10102
rect 70854 10046 70922 10102
rect 70978 10046 71046 10102
rect 71102 10046 71198 10102
rect 70578 9978 71198 10046
rect 70578 9922 70674 9978
rect 70730 9922 70798 9978
rect 70854 9922 70922 9978
rect 70978 9922 71046 9978
rect 71102 9922 71198 9978
rect 70578 -1120 71198 9922
rect 70578 -1176 70674 -1120
rect 70730 -1176 70798 -1120
rect 70854 -1176 70922 -1120
rect 70978 -1176 71046 -1120
rect 71102 -1176 71198 -1120
rect 70578 -1244 71198 -1176
rect 70578 -1300 70674 -1244
rect 70730 -1300 70798 -1244
rect 70854 -1300 70922 -1244
rect 70978 -1300 71046 -1244
rect 71102 -1300 71198 -1244
rect 70578 -1368 71198 -1300
rect 70578 -1424 70674 -1368
rect 70730 -1424 70798 -1368
rect 70854 -1424 70922 -1368
rect 70978 -1424 71046 -1368
rect 71102 -1424 71198 -1368
rect 70578 -1492 71198 -1424
rect 70578 -1548 70674 -1492
rect 70730 -1548 70798 -1492
rect 70854 -1548 70922 -1492
rect 70978 -1548 71046 -1492
rect 71102 -1548 71198 -1492
rect 70578 -1644 71198 -1548
rect 97578 40350 98198 48802
rect 97578 40294 97674 40350
rect 97730 40294 97798 40350
rect 97854 40294 97922 40350
rect 97978 40294 98046 40350
rect 98102 40294 98198 40350
rect 97578 40226 98198 40294
rect 97578 40170 97674 40226
rect 97730 40170 97798 40226
rect 97854 40170 97922 40226
rect 97978 40170 98046 40226
rect 98102 40170 98198 40226
rect 97578 40102 98198 40170
rect 97578 40046 97674 40102
rect 97730 40046 97798 40102
rect 97854 40046 97922 40102
rect 97978 40046 98046 40102
rect 98102 40046 98198 40102
rect 97578 39978 98198 40046
rect 97578 39922 97674 39978
rect 97730 39922 97798 39978
rect 97854 39922 97922 39978
rect 97978 39922 98046 39978
rect 98102 39922 98198 39978
rect 97578 22350 98198 39922
rect 97578 22294 97674 22350
rect 97730 22294 97798 22350
rect 97854 22294 97922 22350
rect 97978 22294 98046 22350
rect 98102 22294 98198 22350
rect 97578 22226 98198 22294
rect 97578 22170 97674 22226
rect 97730 22170 97798 22226
rect 97854 22170 97922 22226
rect 97978 22170 98046 22226
rect 98102 22170 98198 22226
rect 97578 22102 98198 22170
rect 97578 22046 97674 22102
rect 97730 22046 97798 22102
rect 97854 22046 97922 22102
rect 97978 22046 98046 22102
rect 98102 22046 98198 22102
rect 97578 21978 98198 22046
rect 97578 21922 97674 21978
rect 97730 21922 97798 21978
rect 97854 21922 97922 21978
rect 97978 21922 98046 21978
rect 98102 21922 98198 21978
rect 97578 4350 98198 21922
rect 97578 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 98198 4350
rect 97578 4226 98198 4294
rect 97578 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 98198 4226
rect 97578 4102 98198 4170
rect 97578 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 98198 4102
rect 97578 3978 98198 4046
rect 97578 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 98198 3978
rect 97578 -160 98198 3922
rect 97578 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 98198 -160
rect 97578 -284 98198 -216
rect 97578 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 98198 -284
rect 97578 -408 98198 -340
rect 97578 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 98198 -408
rect 97578 -532 98198 -464
rect 97578 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 98198 -532
rect 97578 -1644 98198 -588
rect 101298 46350 101918 48802
rect 101298 46294 101394 46350
rect 101450 46294 101518 46350
rect 101574 46294 101642 46350
rect 101698 46294 101766 46350
rect 101822 46294 101918 46350
rect 101298 46226 101918 46294
rect 101298 46170 101394 46226
rect 101450 46170 101518 46226
rect 101574 46170 101642 46226
rect 101698 46170 101766 46226
rect 101822 46170 101918 46226
rect 101298 46102 101918 46170
rect 101298 46046 101394 46102
rect 101450 46046 101518 46102
rect 101574 46046 101642 46102
rect 101698 46046 101766 46102
rect 101822 46046 101918 46102
rect 101298 45978 101918 46046
rect 101298 45922 101394 45978
rect 101450 45922 101518 45978
rect 101574 45922 101642 45978
rect 101698 45922 101766 45978
rect 101822 45922 101918 45978
rect 101298 28350 101918 45922
rect 101298 28294 101394 28350
rect 101450 28294 101518 28350
rect 101574 28294 101642 28350
rect 101698 28294 101766 28350
rect 101822 28294 101918 28350
rect 101298 28226 101918 28294
rect 101298 28170 101394 28226
rect 101450 28170 101518 28226
rect 101574 28170 101642 28226
rect 101698 28170 101766 28226
rect 101822 28170 101918 28226
rect 101298 28102 101918 28170
rect 101298 28046 101394 28102
rect 101450 28046 101518 28102
rect 101574 28046 101642 28102
rect 101698 28046 101766 28102
rect 101822 28046 101918 28102
rect 101298 27978 101918 28046
rect 101298 27922 101394 27978
rect 101450 27922 101518 27978
rect 101574 27922 101642 27978
rect 101698 27922 101766 27978
rect 101822 27922 101918 27978
rect 101298 10350 101918 27922
rect 101298 10294 101394 10350
rect 101450 10294 101518 10350
rect 101574 10294 101642 10350
rect 101698 10294 101766 10350
rect 101822 10294 101918 10350
rect 101298 10226 101918 10294
rect 101298 10170 101394 10226
rect 101450 10170 101518 10226
rect 101574 10170 101642 10226
rect 101698 10170 101766 10226
rect 101822 10170 101918 10226
rect 101298 10102 101918 10170
rect 101298 10046 101394 10102
rect 101450 10046 101518 10102
rect 101574 10046 101642 10102
rect 101698 10046 101766 10102
rect 101822 10046 101918 10102
rect 101298 9978 101918 10046
rect 101298 9922 101394 9978
rect 101450 9922 101518 9978
rect 101574 9922 101642 9978
rect 101698 9922 101766 9978
rect 101822 9922 101918 9978
rect 101298 -1120 101918 9922
rect 101298 -1176 101394 -1120
rect 101450 -1176 101518 -1120
rect 101574 -1176 101642 -1120
rect 101698 -1176 101766 -1120
rect 101822 -1176 101918 -1120
rect 101298 -1244 101918 -1176
rect 101298 -1300 101394 -1244
rect 101450 -1300 101518 -1244
rect 101574 -1300 101642 -1244
rect 101698 -1300 101766 -1244
rect 101822 -1300 101918 -1244
rect 101298 -1368 101918 -1300
rect 101298 -1424 101394 -1368
rect 101450 -1424 101518 -1368
rect 101574 -1424 101642 -1368
rect 101698 -1424 101766 -1368
rect 101822 -1424 101918 -1368
rect 101298 -1492 101918 -1424
rect 101298 -1548 101394 -1492
rect 101450 -1548 101518 -1492
rect 101574 -1548 101642 -1492
rect 101698 -1548 101766 -1492
rect 101822 -1548 101918 -1492
rect 101298 -1644 101918 -1548
rect 128298 40350 128918 48802
rect 128298 40294 128394 40350
rect 128450 40294 128518 40350
rect 128574 40294 128642 40350
rect 128698 40294 128766 40350
rect 128822 40294 128918 40350
rect 128298 40226 128918 40294
rect 128298 40170 128394 40226
rect 128450 40170 128518 40226
rect 128574 40170 128642 40226
rect 128698 40170 128766 40226
rect 128822 40170 128918 40226
rect 128298 40102 128918 40170
rect 128298 40046 128394 40102
rect 128450 40046 128518 40102
rect 128574 40046 128642 40102
rect 128698 40046 128766 40102
rect 128822 40046 128918 40102
rect 128298 39978 128918 40046
rect 128298 39922 128394 39978
rect 128450 39922 128518 39978
rect 128574 39922 128642 39978
rect 128698 39922 128766 39978
rect 128822 39922 128918 39978
rect 128298 22350 128918 39922
rect 128298 22294 128394 22350
rect 128450 22294 128518 22350
rect 128574 22294 128642 22350
rect 128698 22294 128766 22350
rect 128822 22294 128918 22350
rect 128298 22226 128918 22294
rect 128298 22170 128394 22226
rect 128450 22170 128518 22226
rect 128574 22170 128642 22226
rect 128698 22170 128766 22226
rect 128822 22170 128918 22226
rect 128298 22102 128918 22170
rect 128298 22046 128394 22102
rect 128450 22046 128518 22102
rect 128574 22046 128642 22102
rect 128698 22046 128766 22102
rect 128822 22046 128918 22102
rect 128298 21978 128918 22046
rect 128298 21922 128394 21978
rect 128450 21922 128518 21978
rect 128574 21922 128642 21978
rect 128698 21922 128766 21978
rect 128822 21922 128918 21978
rect 128298 4350 128918 21922
rect 128298 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 128918 4350
rect 128298 4226 128918 4294
rect 128298 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 128918 4226
rect 128298 4102 128918 4170
rect 128298 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 128918 4102
rect 128298 3978 128918 4046
rect 128298 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 128918 3978
rect 128298 -160 128918 3922
rect 128298 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 128918 -160
rect 128298 -284 128918 -216
rect 128298 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 128918 -284
rect 128298 -408 128918 -340
rect 128298 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 128918 -408
rect 128298 -532 128918 -464
rect 128298 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 128918 -532
rect 128298 -1644 128918 -588
rect 132018 46350 132638 48802
rect 132018 46294 132114 46350
rect 132170 46294 132238 46350
rect 132294 46294 132362 46350
rect 132418 46294 132486 46350
rect 132542 46294 132638 46350
rect 132018 46226 132638 46294
rect 132018 46170 132114 46226
rect 132170 46170 132238 46226
rect 132294 46170 132362 46226
rect 132418 46170 132486 46226
rect 132542 46170 132638 46226
rect 132018 46102 132638 46170
rect 132018 46046 132114 46102
rect 132170 46046 132238 46102
rect 132294 46046 132362 46102
rect 132418 46046 132486 46102
rect 132542 46046 132638 46102
rect 132018 45978 132638 46046
rect 132018 45922 132114 45978
rect 132170 45922 132238 45978
rect 132294 45922 132362 45978
rect 132418 45922 132486 45978
rect 132542 45922 132638 45978
rect 132018 28350 132638 45922
rect 132018 28294 132114 28350
rect 132170 28294 132238 28350
rect 132294 28294 132362 28350
rect 132418 28294 132486 28350
rect 132542 28294 132638 28350
rect 132018 28226 132638 28294
rect 132018 28170 132114 28226
rect 132170 28170 132238 28226
rect 132294 28170 132362 28226
rect 132418 28170 132486 28226
rect 132542 28170 132638 28226
rect 132018 28102 132638 28170
rect 132018 28046 132114 28102
rect 132170 28046 132238 28102
rect 132294 28046 132362 28102
rect 132418 28046 132486 28102
rect 132542 28046 132638 28102
rect 132018 27978 132638 28046
rect 132018 27922 132114 27978
rect 132170 27922 132238 27978
rect 132294 27922 132362 27978
rect 132418 27922 132486 27978
rect 132542 27922 132638 27978
rect 132018 10350 132638 27922
rect 132018 10294 132114 10350
rect 132170 10294 132238 10350
rect 132294 10294 132362 10350
rect 132418 10294 132486 10350
rect 132542 10294 132638 10350
rect 132018 10226 132638 10294
rect 132018 10170 132114 10226
rect 132170 10170 132238 10226
rect 132294 10170 132362 10226
rect 132418 10170 132486 10226
rect 132542 10170 132638 10226
rect 132018 10102 132638 10170
rect 132018 10046 132114 10102
rect 132170 10046 132238 10102
rect 132294 10046 132362 10102
rect 132418 10046 132486 10102
rect 132542 10046 132638 10102
rect 132018 9978 132638 10046
rect 132018 9922 132114 9978
rect 132170 9922 132238 9978
rect 132294 9922 132362 9978
rect 132418 9922 132486 9978
rect 132542 9922 132638 9978
rect 132018 -1120 132638 9922
rect 132018 -1176 132114 -1120
rect 132170 -1176 132238 -1120
rect 132294 -1176 132362 -1120
rect 132418 -1176 132486 -1120
rect 132542 -1176 132638 -1120
rect 132018 -1244 132638 -1176
rect 132018 -1300 132114 -1244
rect 132170 -1300 132238 -1244
rect 132294 -1300 132362 -1244
rect 132418 -1300 132486 -1244
rect 132542 -1300 132638 -1244
rect 132018 -1368 132638 -1300
rect 132018 -1424 132114 -1368
rect 132170 -1424 132238 -1368
rect 132294 -1424 132362 -1368
rect 132418 -1424 132486 -1368
rect 132542 -1424 132638 -1368
rect 132018 -1492 132638 -1424
rect 132018 -1548 132114 -1492
rect 132170 -1548 132238 -1492
rect 132294 -1548 132362 -1492
rect 132418 -1548 132486 -1492
rect 132542 -1548 132638 -1492
rect 132018 -1644 132638 -1548
rect 159018 40350 159638 48802
rect 159018 40294 159114 40350
rect 159170 40294 159238 40350
rect 159294 40294 159362 40350
rect 159418 40294 159486 40350
rect 159542 40294 159638 40350
rect 159018 40226 159638 40294
rect 159018 40170 159114 40226
rect 159170 40170 159238 40226
rect 159294 40170 159362 40226
rect 159418 40170 159486 40226
rect 159542 40170 159638 40226
rect 159018 40102 159638 40170
rect 159018 40046 159114 40102
rect 159170 40046 159238 40102
rect 159294 40046 159362 40102
rect 159418 40046 159486 40102
rect 159542 40046 159638 40102
rect 159018 39978 159638 40046
rect 159018 39922 159114 39978
rect 159170 39922 159238 39978
rect 159294 39922 159362 39978
rect 159418 39922 159486 39978
rect 159542 39922 159638 39978
rect 159018 22350 159638 39922
rect 159018 22294 159114 22350
rect 159170 22294 159238 22350
rect 159294 22294 159362 22350
rect 159418 22294 159486 22350
rect 159542 22294 159638 22350
rect 159018 22226 159638 22294
rect 159018 22170 159114 22226
rect 159170 22170 159238 22226
rect 159294 22170 159362 22226
rect 159418 22170 159486 22226
rect 159542 22170 159638 22226
rect 159018 22102 159638 22170
rect 159018 22046 159114 22102
rect 159170 22046 159238 22102
rect 159294 22046 159362 22102
rect 159418 22046 159486 22102
rect 159542 22046 159638 22102
rect 159018 21978 159638 22046
rect 159018 21922 159114 21978
rect 159170 21922 159238 21978
rect 159294 21922 159362 21978
rect 159418 21922 159486 21978
rect 159542 21922 159638 21978
rect 159018 4350 159638 21922
rect 159018 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 159638 4350
rect 159018 4226 159638 4294
rect 159018 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 159638 4226
rect 159018 4102 159638 4170
rect 159018 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 159638 4102
rect 159018 3978 159638 4046
rect 159018 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 159638 3978
rect 159018 -160 159638 3922
rect 159018 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 159638 -160
rect 159018 -284 159638 -216
rect 159018 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 159638 -284
rect 159018 -408 159638 -340
rect 159018 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 159638 -408
rect 159018 -532 159638 -464
rect 159018 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 159638 -532
rect 159018 -1644 159638 -588
rect 162738 46350 163358 48802
rect 162738 46294 162834 46350
rect 162890 46294 162958 46350
rect 163014 46294 163082 46350
rect 163138 46294 163206 46350
rect 163262 46294 163358 46350
rect 162738 46226 163358 46294
rect 162738 46170 162834 46226
rect 162890 46170 162958 46226
rect 163014 46170 163082 46226
rect 163138 46170 163206 46226
rect 163262 46170 163358 46226
rect 162738 46102 163358 46170
rect 162738 46046 162834 46102
rect 162890 46046 162958 46102
rect 163014 46046 163082 46102
rect 163138 46046 163206 46102
rect 163262 46046 163358 46102
rect 162738 45978 163358 46046
rect 162738 45922 162834 45978
rect 162890 45922 162958 45978
rect 163014 45922 163082 45978
rect 163138 45922 163206 45978
rect 163262 45922 163358 45978
rect 162738 28350 163358 45922
rect 162738 28294 162834 28350
rect 162890 28294 162958 28350
rect 163014 28294 163082 28350
rect 163138 28294 163206 28350
rect 163262 28294 163358 28350
rect 162738 28226 163358 28294
rect 162738 28170 162834 28226
rect 162890 28170 162958 28226
rect 163014 28170 163082 28226
rect 163138 28170 163206 28226
rect 163262 28170 163358 28226
rect 162738 28102 163358 28170
rect 162738 28046 162834 28102
rect 162890 28046 162958 28102
rect 163014 28046 163082 28102
rect 163138 28046 163206 28102
rect 163262 28046 163358 28102
rect 162738 27978 163358 28046
rect 162738 27922 162834 27978
rect 162890 27922 162958 27978
rect 163014 27922 163082 27978
rect 163138 27922 163206 27978
rect 163262 27922 163358 27978
rect 162738 10350 163358 27922
rect 162738 10294 162834 10350
rect 162890 10294 162958 10350
rect 163014 10294 163082 10350
rect 163138 10294 163206 10350
rect 163262 10294 163358 10350
rect 162738 10226 163358 10294
rect 162738 10170 162834 10226
rect 162890 10170 162958 10226
rect 163014 10170 163082 10226
rect 163138 10170 163206 10226
rect 163262 10170 163358 10226
rect 162738 10102 163358 10170
rect 162738 10046 162834 10102
rect 162890 10046 162958 10102
rect 163014 10046 163082 10102
rect 163138 10046 163206 10102
rect 163262 10046 163358 10102
rect 162738 9978 163358 10046
rect 162738 9922 162834 9978
rect 162890 9922 162958 9978
rect 163014 9922 163082 9978
rect 163138 9922 163206 9978
rect 163262 9922 163358 9978
rect 162738 -1120 163358 9922
rect 162738 -1176 162834 -1120
rect 162890 -1176 162958 -1120
rect 163014 -1176 163082 -1120
rect 163138 -1176 163206 -1120
rect 163262 -1176 163358 -1120
rect 162738 -1244 163358 -1176
rect 162738 -1300 162834 -1244
rect 162890 -1300 162958 -1244
rect 163014 -1300 163082 -1244
rect 163138 -1300 163206 -1244
rect 163262 -1300 163358 -1244
rect 162738 -1368 163358 -1300
rect 162738 -1424 162834 -1368
rect 162890 -1424 162958 -1368
rect 163014 -1424 163082 -1368
rect 163138 -1424 163206 -1368
rect 163262 -1424 163358 -1368
rect 162738 -1492 163358 -1424
rect 162738 -1548 162834 -1492
rect 162890 -1548 162958 -1492
rect 163014 -1548 163082 -1492
rect 163138 -1548 163206 -1492
rect 163262 -1548 163358 -1492
rect 162738 -1644 163358 -1548
rect 189738 40350 190358 48802
rect 189738 40294 189834 40350
rect 189890 40294 189958 40350
rect 190014 40294 190082 40350
rect 190138 40294 190206 40350
rect 190262 40294 190358 40350
rect 189738 40226 190358 40294
rect 189738 40170 189834 40226
rect 189890 40170 189958 40226
rect 190014 40170 190082 40226
rect 190138 40170 190206 40226
rect 190262 40170 190358 40226
rect 189738 40102 190358 40170
rect 189738 40046 189834 40102
rect 189890 40046 189958 40102
rect 190014 40046 190082 40102
rect 190138 40046 190206 40102
rect 190262 40046 190358 40102
rect 189738 39978 190358 40046
rect 189738 39922 189834 39978
rect 189890 39922 189958 39978
rect 190014 39922 190082 39978
rect 190138 39922 190206 39978
rect 190262 39922 190358 39978
rect 189738 22350 190358 39922
rect 189738 22294 189834 22350
rect 189890 22294 189958 22350
rect 190014 22294 190082 22350
rect 190138 22294 190206 22350
rect 190262 22294 190358 22350
rect 189738 22226 190358 22294
rect 189738 22170 189834 22226
rect 189890 22170 189958 22226
rect 190014 22170 190082 22226
rect 190138 22170 190206 22226
rect 190262 22170 190358 22226
rect 189738 22102 190358 22170
rect 189738 22046 189834 22102
rect 189890 22046 189958 22102
rect 190014 22046 190082 22102
rect 190138 22046 190206 22102
rect 190262 22046 190358 22102
rect 189738 21978 190358 22046
rect 189738 21922 189834 21978
rect 189890 21922 189958 21978
rect 190014 21922 190082 21978
rect 190138 21922 190206 21978
rect 190262 21922 190358 21978
rect 189738 4350 190358 21922
rect 189738 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 190358 4350
rect 189738 4226 190358 4294
rect 189738 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 190358 4226
rect 189738 4102 190358 4170
rect 189738 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 190358 4102
rect 189738 3978 190358 4046
rect 189738 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 190358 3978
rect 189738 -160 190358 3922
rect 189738 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 190358 -160
rect 189738 -284 190358 -216
rect 189738 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 190358 -284
rect 189738 -408 190358 -340
rect 189738 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 190358 -408
rect 189738 -532 190358 -464
rect 189738 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 190358 -532
rect 189738 -1644 190358 -588
rect 193458 46350 194078 48802
rect 193458 46294 193554 46350
rect 193610 46294 193678 46350
rect 193734 46294 193802 46350
rect 193858 46294 193926 46350
rect 193982 46294 194078 46350
rect 193458 46226 194078 46294
rect 193458 46170 193554 46226
rect 193610 46170 193678 46226
rect 193734 46170 193802 46226
rect 193858 46170 193926 46226
rect 193982 46170 194078 46226
rect 193458 46102 194078 46170
rect 193458 46046 193554 46102
rect 193610 46046 193678 46102
rect 193734 46046 193802 46102
rect 193858 46046 193926 46102
rect 193982 46046 194078 46102
rect 193458 45978 194078 46046
rect 193458 45922 193554 45978
rect 193610 45922 193678 45978
rect 193734 45922 193802 45978
rect 193858 45922 193926 45978
rect 193982 45922 194078 45978
rect 193458 28350 194078 45922
rect 193458 28294 193554 28350
rect 193610 28294 193678 28350
rect 193734 28294 193802 28350
rect 193858 28294 193926 28350
rect 193982 28294 194078 28350
rect 193458 28226 194078 28294
rect 193458 28170 193554 28226
rect 193610 28170 193678 28226
rect 193734 28170 193802 28226
rect 193858 28170 193926 28226
rect 193982 28170 194078 28226
rect 193458 28102 194078 28170
rect 193458 28046 193554 28102
rect 193610 28046 193678 28102
rect 193734 28046 193802 28102
rect 193858 28046 193926 28102
rect 193982 28046 194078 28102
rect 193458 27978 194078 28046
rect 193458 27922 193554 27978
rect 193610 27922 193678 27978
rect 193734 27922 193802 27978
rect 193858 27922 193926 27978
rect 193982 27922 194078 27978
rect 193458 10350 194078 27922
rect 193458 10294 193554 10350
rect 193610 10294 193678 10350
rect 193734 10294 193802 10350
rect 193858 10294 193926 10350
rect 193982 10294 194078 10350
rect 193458 10226 194078 10294
rect 193458 10170 193554 10226
rect 193610 10170 193678 10226
rect 193734 10170 193802 10226
rect 193858 10170 193926 10226
rect 193982 10170 194078 10226
rect 193458 10102 194078 10170
rect 193458 10046 193554 10102
rect 193610 10046 193678 10102
rect 193734 10046 193802 10102
rect 193858 10046 193926 10102
rect 193982 10046 194078 10102
rect 193458 9978 194078 10046
rect 193458 9922 193554 9978
rect 193610 9922 193678 9978
rect 193734 9922 193802 9978
rect 193858 9922 193926 9978
rect 193982 9922 194078 9978
rect 193458 -1120 194078 9922
rect 193458 -1176 193554 -1120
rect 193610 -1176 193678 -1120
rect 193734 -1176 193802 -1120
rect 193858 -1176 193926 -1120
rect 193982 -1176 194078 -1120
rect 193458 -1244 194078 -1176
rect 193458 -1300 193554 -1244
rect 193610 -1300 193678 -1244
rect 193734 -1300 193802 -1244
rect 193858 -1300 193926 -1244
rect 193982 -1300 194078 -1244
rect 193458 -1368 194078 -1300
rect 193458 -1424 193554 -1368
rect 193610 -1424 193678 -1368
rect 193734 -1424 193802 -1368
rect 193858 -1424 193926 -1368
rect 193982 -1424 194078 -1368
rect 193458 -1492 194078 -1424
rect 193458 -1548 193554 -1492
rect 193610 -1548 193678 -1492
rect 193734 -1548 193802 -1492
rect 193858 -1548 193926 -1492
rect 193982 -1548 194078 -1492
rect 193458 -1644 194078 -1548
rect 220458 40350 221078 48802
rect 220458 40294 220554 40350
rect 220610 40294 220678 40350
rect 220734 40294 220802 40350
rect 220858 40294 220926 40350
rect 220982 40294 221078 40350
rect 220458 40226 221078 40294
rect 220458 40170 220554 40226
rect 220610 40170 220678 40226
rect 220734 40170 220802 40226
rect 220858 40170 220926 40226
rect 220982 40170 221078 40226
rect 220458 40102 221078 40170
rect 220458 40046 220554 40102
rect 220610 40046 220678 40102
rect 220734 40046 220802 40102
rect 220858 40046 220926 40102
rect 220982 40046 221078 40102
rect 220458 39978 221078 40046
rect 220458 39922 220554 39978
rect 220610 39922 220678 39978
rect 220734 39922 220802 39978
rect 220858 39922 220926 39978
rect 220982 39922 221078 39978
rect 220458 22350 221078 39922
rect 220458 22294 220554 22350
rect 220610 22294 220678 22350
rect 220734 22294 220802 22350
rect 220858 22294 220926 22350
rect 220982 22294 221078 22350
rect 220458 22226 221078 22294
rect 220458 22170 220554 22226
rect 220610 22170 220678 22226
rect 220734 22170 220802 22226
rect 220858 22170 220926 22226
rect 220982 22170 221078 22226
rect 220458 22102 221078 22170
rect 220458 22046 220554 22102
rect 220610 22046 220678 22102
rect 220734 22046 220802 22102
rect 220858 22046 220926 22102
rect 220982 22046 221078 22102
rect 220458 21978 221078 22046
rect 220458 21922 220554 21978
rect 220610 21922 220678 21978
rect 220734 21922 220802 21978
rect 220858 21922 220926 21978
rect 220982 21922 221078 21978
rect 220458 4350 221078 21922
rect 220458 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 221078 4350
rect 220458 4226 221078 4294
rect 220458 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 221078 4226
rect 220458 4102 221078 4170
rect 220458 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 221078 4102
rect 220458 3978 221078 4046
rect 220458 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 221078 3978
rect 220458 -160 221078 3922
rect 220458 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 221078 -160
rect 220458 -284 221078 -216
rect 220458 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 221078 -284
rect 220458 -408 221078 -340
rect 220458 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 221078 -408
rect 220458 -532 221078 -464
rect 220458 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 221078 -532
rect 220458 -1644 221078 -588
rect 224178 46350 224798 48802
rect 224178 46294 224274 46350
rect 224330 46294 224398 46350
rect 224454 46294 224522 46350
rect 224578 46294 224646 46350
rect 224702 46294 224798 46350
rect 224178 46226 224798 46294
rect 224178 46170 224274 46226
rect 224330 46170 224398 46226
rect 224454 46170 224522 46226
rect 224578 46170 224646 46226
rect 224702 46170 224798 46226
rect 224178 46102 224798 46170
rect 224178 46046 224274 46102
rect 224330 46046 224398 46102
rect 224454 46046 224522 46102
rect 224578 46046 224646 46102
rect 224702 46046 224798 46102
rect 224178 45978 224798 46046
rect 224178 45922 224274 45978
rect 224330 45922 224398 45978
rect 224454 45922 224522 45978
rect 224578 45922 224646 45978
rect 224702 45922 224798 45978
rect 224178 28350 224798 45922
rect 224178 28294 224274 28350
rect 224330 28294 224398 28350
rect 224454 28294 224522 28350
rect 224578 28294 224646 28350
rect 224702 28294 224798 28350
rect 224178 28226 224798 28294
rect 224178 28170 224274 28226
rect 224330 28170 224398 28226
rect 224454 28170 224522 28226
rect 224578 28170 224646 28226
rect 224702 28170 224798 28226
rect 224178 28102 224798 28170
rect 224178 28046 224274 28102
rect 224330 28046 224398 28102
rect 224454 28046 224522 28102
rect 224578 28046 224646 28102
rect 224702 28046 224798 28102
rect 224178 27978 224798 28046
rect 224178 27922 224274 27978
rect 224330 27922 224398 27978
rect 224454 27922 224522 27978
rect 224578 27922 224646 27978
rect 224702 27922 224798 27978
rect 224178 10350 224798 27922
rect 224178 10294 224274 10350
rect 224330 10294 224398 10350
rect 224454 10294 224522 10350
rect 224578 10294 224646 10350
rect 224702 10294 224798 10350
rect 224178 10226 224798 10294
rect 224178 10170 224274 10226
rect 224330 10170 224398 10226
rect 224454 10170 224522 10226
rect 224578 10170 224646 10226
rect 224702 10170 224798 10226
rect 224178 10102 224798 10170
rect 224178 10046 224274 10102
rect 224330 10046 224398 10102
rect 224454 10046 224522 10102
rect 224578 10046 224646 10102
rect 224702 10046 224798 10102
rect 224178 9978 224798 10046
rect 224178 9922 224274 9978
rect 224330 9922 224398 9978
rect 224454 9922 224522 9978
rect 224578 9922 224646 9978
rect 224702 9922 224798 9978
rect 224178 -1120 224798 9922
rect 224178 -1176 224274 -1120
rect 224330 -1176 224398 -1120
rect 224454 -1176 224522 -1120
rect 224578 -1176 224646 -1120
rect 224702 -1176 224798 -1120
rect 224178 -1244 224798 -1176
rect 224178 -1300 224274 -1244
rect 224330 -1300 224398 -1244
rect 224454 -1300 224522 -1244
rect 224578 -1300 224646 -1244
rect 224702 -1300 224798 -1244
rect 224178 -1368 224798 -1300
rect 224178 -1424 224274 -1368
rect 224330 -1424 224398 -1368
rect 224454 -1424 224522 -1368
rect 224578 -1424 224646 -1368
rect 224702 -1424 224798 -1368
rect 224178 -1492 224798 -1424
rect 224178 -1548 224274 -1492
rect 224330 -1548 224398 -1492
rect 224454 -1548 224522 -1492
rect 224578 -1548 224646 -1492
rect 224702 -1548 224798 -1492
rect 224178 -1644 224798 -1548
rect 251178 40350 251798 48802
rect 251178 40294 251274 40350
rect 251330 40294 251398 40350
rect 251454 40294 251522 40350
rect 251578 40294 251646 40350
rect 251702 40294 251798 40350
rect 251178 40226 251798 40294
rect 251178 40170 251274 40226
rect 251330 40170 251398 40226
rect 251454 40170 251522 40226
rect 251578 40170 251646 40226
rect 251702 40170 251798 40226
rect 251178 40102 251798 40170
rect 251178 40046 251274 40102
rect 251330 40046 251398 40102
rect 251454 40046 251522 40102
rect 251578 40046 251646 40102
rect 251702 40046 251798 40102
rect 251178 39978 251798 40046
rect 251178 39922 251274 39978
rect 251330 39922 251398 39978
rect 251454 39922 251522 39978
rect 251578 39922 251646 39978
rect 251702 39922 251798 39978
rect 251178 22350 251798 39922
rect 251178 22294 251274 22350
rect 251330 22294 251398 22350
rect 251454 22294 251522 22350
rect 251578 22294 251646 22350
rect 251702 22294 251798 22350
rect 251178 22226 251798 22294
rect 251178 22170 251274 22226
rect 251330 22170 251398 22226
rect 251454 22170 251522 22226
rect 251578 22170 251646 22226
rect 251702 22170 251798 22226
rect 251178 22102 251798 22170
rect 251178 22046 251274 22102
rect 251330 22046 251398 22102
rect 251454 22046 251522 22102
rect 251578 22046 251646 22102
rect 251702 22046 251798 22102
rect 251178 21978 251798 22046
rect 251178 21922 251274 21978
rect 251330 21922 251398 21978
rect 251454 21922 251522 21978
rect 251578 21922 251646 21978
rect 251702 21922 251798 21978
rect 251178 4350 251798 21922
rect 251178 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 251798 4350
rect 251178 4226 251798 4294
rect 251178 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 251798 4226
rect 251178 4102 251798 4170
rect 251178 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 251798 4102
rect 251178 3978 251798 4046
rect 251178 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 251798 3978
rect 251178 -160 251798 3922
rect 251178 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 251798 -160
rect 251178 -284 251798 -216
rect 251178 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 251798 -284
rect 251178 -408 251798 -340
rect 251178 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 251798 -408
rect 251178 -532 251798 -464
rect 251178 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 251798 -532
rect 251178 -1644 251798 -588
rect 254898 46350 255518 48802
rect 267148 47908 267204 249340
rect 267372 246372 267428 246382
rect 267372 220108 267428 246316
rect 268716 246178 268772 246188
rect 268716 245364 268772 246122
rect 268716 245298 268772 245308
rect 267260 220052 267428 220108
rect 267260 48580 267316 220052
rect 269276 148820 269332 257292
rect 281898 256350 282518 257490
rect 281898 256294 281994 256350
rect 282050 256294 282118 256350
rect 282174 256294 282242 256350
rect 282298 256294 282366 256350
rect 282422 256294 282518 256350
rect 273868 256228 273924 256238
rect 270508 252838 270564 252848
rect 269612 252478 269668 252488
rect 269500 252118 269556 252128
rect 269388 214340 269444 214350
rect 269388 172116 269444 214284
rect 269388 172050 269444 172060
rect 269276 148754 269332 148764
rect 267260 48514 267316 48524
rect 267148 47842 267204 47852
rect 254898 46294 254994 46350
rect 255050 46294 255118 46350
rect 255174 46294 255242 46350
rect 255298 46294 255366 46350
rect 255422 46294 255518 46350
rect 254898 46226 255518 46294
rect 254898 46170 254994 46226
rect 255050 46170 255118 46226
rect 255174 46170 255242 46226
rect 255298 46170 255366 46226
rect 255422 46170 255518 46226
rect 254898 46102 255518 46170
rect 254898 46046 254994 46102
rect 255050 46046 255118 46102
rect 255174 46046 255242 46102
rect 255298 46046 255366 46102
rect 255422 46046 255518 46102
rect 254898 45978 255518 46046
rect 254898 45922 254994 45978
rect 255050 45922 255118 45978
rect 255174 45922 255242 45978
rect 255298 45922 255366 45978
rect 255422 45922 255518 45978
rect 254898 28350 255518 45922
rect 269500 33012 269556 252062
rect 269612 34692 269668 252422
rect 269724 217812 269780 217822
rect 269724 160468 269780 217756
rect 269836 211092 269892 211102
rect 269836 201572 269892 211036
rect 269836 201506 269892 201516
rect 269724 160402 269780 160412
rect 270508 36148 270564 252782
rect 270620 234388 270676 234398
rect 270620 157556 270676 234332
rect 270732 216580 270788 216590
rect 270732 169204 270788 216524
rect 272412 211316 272468 211326
rect 272412 209860 272468 211260
rect 272412 209794 272468 209804
rect 272748 210756 272804 210766
rect 272636 209412 272692 209422
rect 272524 209076 272580 209086
rect 272524 208348 272580 209020
rect 272412 208292 272580 208348
rect 272412 189588 272468 208292
rect 272636 196588 272692 209356
rect 272524 196532 272692 196588
rect 272524 192500 272580 196532
rect 272524 192434 272580 192444
rect 272412 189522 272468 189532
rect 272748 183764 272804 210700
rect 272860 209524 272916 209534
rect 272860 186676 272916 209468
rect 273196 209300 273252 209310
rect 273084 209188 273140 209198
rect 273084 195412 273140 209132
rect 273196 198324 273252 209244
rect 273196 198258 273252 198268
rect 273084 195346 273140 195356
rect 272860 186610 272916 186620
rect 272748 183698 272804 183708
rect 270732 169138 270788 169148
rect 273868 163380 273924 256172
rect 281898 256226 282518 256294
rect 281898 256170 281994 256226
rect 282050 256170 282118 256226
rect 282174 256170 282242 256226
rect 282298 256170 282366 256226
rect 282422 256170 282518 256226
rect 281898 256102 282518 256170
rect 281898 256046 281994 256102
rect 282050 256046 282118 256102
rect 282174 256046 282242 256102
rect 282298 256046 282366 256102
rect 282422 256046 282518 256102
rect 281898 255978 282518 256046
rect 281898 255922 281994 255978
rect 282050 255922 282118 255978
rect 282174 255922 282242 255978
rect 282298 255922 282366 255978
rect 282422 255922 282518 255978
rect 273980 254660 274036 254670
rect 273980 166292 274036 254604
rect 275548 252658 275604 252668
rect 274652 249418 274708 249428
rect 274204 216356 274260 216366
rect 273980 166226 274036 166236
rect 274092 213220 274148 213230
rect 273868 163314 273924 163324
rect 270620 157490 270676 157500
rect 274092 154644 274148 213164
rect 274204 175028 274260 216300
rect 274204 174962 274260 174972
rect 274652 156324 274708 249362
rect 274652 156258 274708 156268
rect 274092 154578 274148 154588
rect 273756 154084 273812 154094
rect 273756 152938 273812 154028
rect 273756 136164 273812 152882
rect 273756 136098 273812 136108
rect 270508 36082 270564 36092
rect 275548 34916 275604 252602
rect 275660 252298 275716 252308
rect 275660 48132 275716 252242
rect 281898 238350 282518 255922
rect 281898 238294 281994 238350
rect 282050 238294 282118 238350
rect 282174 238294 282242 238350
rect 282298 238294 282366 238350
rect 282422 238294 282518 238350
rect 281898 238226 282518 238294
rect 281898 238170 281994 238226
rect 282050 238170 282118 238226
rect 282174 238170 282242 238226
rect 282298 238170 282366 238226
rect 282422 238170 282518 238226
rect 281898 238102 282518 238170
rect 281898 238046 281994 238102
rect 282050 238046 282118 238102
rect 282174 238046 282242 238102
rect 282298 238046 282366 238102
rect 282422 238046 282518 238102
rect 281898 237978 282518 238046
rect 281898 237922 281994 237978
rect 282050 237922 282118 237978
rect 282174 237922 282242 237978
rect 282298 237922 282366 237978
rect 282422 237922 282518 237978
rect 281898 220350 282518 237922
rect 281898 220294 281994 220350
rect 282050 220294 282118 220350
rect 282174 220294 282242 220350
rect 282298 220294 282366 220350
rect 282422 220294 282518 220350
rect 281898 220226 282518 220294
rect 281898 220170 281994 220226
rect 282050 220170 282118 220226
rect 282174 220170 282242 220226
rect 282298 220170 282366 220226
rect 282422 220170 282518 220226
rect 281898 220102 282518 220170
rect 281898 220046 281994 220102
rect 282050 220046 282118 220102
rect 282174 220046 282242 220102
rect 282298 220046 282366 220102
rect 282422 220046 282518 220102
rect 281898 219978 282518 220046
rect 281898 219922 281994 219978
rect 282050 219922 282118 219978
rect 282174 219922 282242 219978
rect 282298 219922 282366 219978
rect 282422 219922 282518 219978
rect 275772 212996 275828 213006
rect 275772 177940 275828 212940
rect 275772 177874 275828 177884
rect 281898 202350 282518 219922
rect 281898 202294 281994 202350
rect 282050 202294 282118 202350
rect 282174 202294 282242 202350
rect 282298 202294 282366 202350
rect 282422 202294 282518 202350
rect 281898 202226 282518 202294
rect 281898 202170 281994 202226
rect 282050 202170 282118 202226
rect 282174 202170 282242 202226
rect 282298 202170 282366 202226
rect 282422 202170 282518 202226
rect 281898 202102 282518 202170
rect 281898 202046 281994 202102
rect 282050 202046 282118 202102
rect 282174 202046 282242 202102
rect 282298 202046 282366 202102
rect 282422 202046 282518 202102
rect 281898 201978 282518 202046
rect 281898 201922 281994 201978
rect 282050 201922 282118 201978
rect 282174 201922 282242 201978
rect 282298 201922 282366 201978
rect 282422 201922 282518 201978
rect 281898 184350 282518 201922
rect 281898 184294 281994 184350
rect 282050 184294 282118 184350
rect 282174 184294 282242 184350
rect 282298 184294 282366 184350
rect 282422 184294 282518 184350
rect 281898 184226 282518 184294
rect 281898 184170 281994 184226
rect 282050 184170 282118 184226
rect 282174 184170 282242 184226
rect 282298 184170 282366 184226
rect 282422 184170 282518 184226
rect 281898 184102 282518 184170
rect 281898 184046 281994 184102
rect 282050 184046 282118 184102
rect 282174 184046 282242 184102
rect 282298 184046 282366 184102
rect 282422 184046 282518 184102
rect 281898 183978 282518 184046
rect 281898 183922 281994 183978
rect 282050 183922 282118 183978
rect 282174 183922 282242 183978
rect 282298 183922 282366 183978
rect 282422 183922 282518 183978
rect 275660 48066 275716 48076
rect 281898 166350 282518 183922
rect 281898 166294 281994 166350
rect 282050 166294 282118 166350
rect 282174 166294 282242 166350
rect 282298 166294 282366 166350
rect 282422 166294 282518 166350
rect 281898 166226 282518 166294
rect 281898 166170 281994 166226
rect 282050 166170 282118 166226
rect 282174 166170 282242 166226
rect 282298 166170 282366 166226
rect 282422 166170 282518 166226
rect 281898 166102 282518 166170
rect 281898 166046 281994 166102
rect 282050 166046 282118 166102
rect 282174 166046 282242 166102
rect 282298 166046 282366 166102
rect 282422 166046 282518 166102
rect 281898 165978 282518 166046
rect 281898 165922 281994 165978
rect 282050 165922 282118 165978
rect 282174 165922 282242 165978
rect 282298 165922 282366 165978
rect 282422 165922 282518 165978
rect 281898 148350 282518 165922
rect 281898 148294 281994 148350
rect 282050 148294 282118 148350
rect 282174 148294 282242 148350
rect 282298 148294 282366 148350
rect 282422 148294 282518 148350
rect 281898 148226 282518 148294
rect 281898 148170 281994 148226
rect 282050 148170 282118 148226
rect 282174 148170 282242 148226
rect 282298 148170 282366 148226
rect 282422 148170 282518 148226
rect 281898 148102 282518 148170
rect 281898 148046 281994 148102
rect 282050 148046 282118 148102
rect 282174 148046 282242 148102
rect 282298 148046 282366 148102
rect 282422 148046 282518 148102
rect 281898 147978 282518 148046
rect 281898 147922 281994 147978
rect 282050 147922 282118 147978
rect 282174 147922 282242 147978
rect 282298 147922 282366 147978
rect 282422 147922 282518 147978
rect 281898 130350 282518 147922
rect 281898 130294 281994 130350
rect 282050 130294 282118 130350
rect 282174 130294 282242 130350
rect 282298 130294 282366 130350
rect 282422 130294 282518 130350
rect 281898 130226 282518 130294
rect 281898 130170 281994 130226
rect 282050 130170 282118 130226
rect 282174 130170 282242 130226
rect 282298 130170 282366 130226
rect 282422 130170 282518 130226
rect 281898 130102 282518 130170
rect 281898 130046 281994 130102
rect 282050 130046 282118 130102
rect 282174 130046 282242 130102
rect 282298 130046 282366 130102
rect 282422 130046 282518 130102
rect 281898 129978 282518 130046
rect 281898 129922 281994 129978
rect 282050 129922 282118 129978
rect 282174 129922 282242 129978
rect 282298 129922 282366 129978
rect 282422 129922 282518 129978
rect 281898 112350 282518 129922
rect 281898 112294 281994 112350
rect 282050 112294 282118 112350
rect 282174 112294 282242 112350
rect 282298 112294 282366 112350
rect 282422 112294 282518 112350
rect 281898 112226 282518 112294
rect 281898 112170 281994 112226
rect 282050 112170 282118 112226
rect 282174 112170 282242 112226
rect 282298 112170 282366 112226
rect 282422 112170 282518 112226
rect 281898 112102 282518 112170
rect 281898 112046 281994 112102
rect 282050 112046 282118 112102
rect 282174 112046 282242 112102
rect 282298 112046 282366 112102
rect 282422 112046 282518 112102
rect 281898 111978 282518 112046
rect 281898 111922 281994 111978
rect 282050 111922 282118 111978
rect 282174 111922 282242 111978
rect 282298 111922 282366 111978
rect 282422 111922 282518 111978
rect 281898 94350 282518 111922
rect 281898 94294 281994 94350
rect 282050 94294 282118 94350
rect 282174 94294 282242 94350
rect 282298 94294 282366 94350
rect 282422 94294 282518 94350
rect 281898 94226 282518 94294
rect 281898 94170 281994 94226
rect 282050 94170 282118 94226
rect 282174 94170 282242 94226
rect 282298 94170 282366 94226
rect 282422 94170 282518 94226
rect 281898 94102 282518 94170
rect 281898 94046 281994 94102
rect 282050 94046 282118 94102
rect 282174 94046 282242 94102
rect 282298 94046 282366 94102
rect 282422 94046 282518 94102
rect 281898 93978 282518 94046
rect 281898 93922 281994 93978
rect 282050 93922 282118 93978
rect 282174 93922 282242 93978
rect 282298 93922 282366 93978
rect 282422 93922 282518 93978
rect 281898 76350 282518 93922
rect 281898 76294 281994 76350
rect 282050 76294 282118 76350
rect 282174 76294 282242 76350
rect 282298 76294 282366 76350
rect 282422 76294 282518 76350
rect 281898 76226 282518 76294
rect 281898 76170 281994 76226
rect 282050 76170 282118 76226
rect 282174 76170 282242 76226
rect 282298 76170 282366 76226
rect 282422 76170 282518 76226
rect 281898 76102 282518 76170
rect 281898 76046 281994 76102
rect 282050 76046 282118 76102
rect 282174 76046 282242 76102
rect 282298 76046 282366 76102
rect 282422 76046 282518 76102
rect 281898 75978 282518 76046
rect 281898 75922 281994 75978
rect 282050 75922 282118 75978
rect 282174 75922 282242 75978
rect 282298 75922 282366 75978
rect 282422 75922 282518 75978
rect 281898 58350 282518 75922
rect 281898 58294 281994 58350
rect 282050 58294 282118 58350
rect 282174 58294 282242 58350
rect 282298 58294 282366 58350
rect 282422 58294 282518 58350
rect 281898 58226 282518 58294
rect 281898 58170 281994 58226
rect 282050 58170 282118 58226
rect 282174 58170 282242 58226
rect 282298 58170 282366 58226
rect 282422 58170 282518 58226
rect 281898 58102 282518 58170
rect 281898 58046 281994 58102
rect 282050 58046 282118 58102
rect 282174 58046 282242 58102
rect 282298 58046 282366 58102
rect 282422 58046 282518 58102
rect 281898 57978 282518 58046
rect 281898 57922 281994 57978
rect 282050 57922 282118 57978
rect 282174 57922 282242 57978
rect 282298 57922 282366 57978
rect 282422 57922 282518 57978
rect 275548 34850 275604 34860
rect 281898 40350 282518 57922
rect 281898 40294 281994 40350
rect 282050 40294 282118 40350
rect 282174 40294 282242 40350
rect 282298 40294 282366 40350
rect 282422 40294 282518 40350
rect 281898 40226 282518 40294
rect 281898 40170 281994 40226
rect 282050 40170 282118 40226
rect 282174 40170 282242 40226
rect 282298 40170 282366 40226
rect 282422 40170 282518 40226
rect 281898 40102 282518 40170
rect 281898 40046 281994 40102
rect 282050 40046 282118 40102
rect 282174 40046 282242 40102
rect 282298 40046 282366 40102
rect 282422 40046 282518 40102
rect 281898 39978 282518 40046
rect 281898 39922 281994 39978
rect 282050 39922 282118 39978
rect 282174 39922 282242 39978
rect 282298 39922 282366 39978
rect 282422 39922 282518 39978
rect 269612 34626 269668 34636
rect 269500 32946 269556 32956
rect 254898 28294 254994 28350
rect 255050 28294 255118 28350
rect 255174 28294 255242 28350
rect 255298 28294 255366 28350
rect 255422 28294 255518 28350
rect 254898 28226 255518 28294
rect 254898 28170 254994 28226
rect 255050 28170 255118 28226
rect 255174 28170 255242 28226
rect 255298 28170 255366 28226
rect 255422 28170 255518 28226
rect 254898 28102 255518 28170
rect 254898 28046 254994 28102
rect 255050 28046 255118 28102
rect 255174 28046 255242 28102
rect 255298 28046 255366 28102
rect 255422 28046 255518 28102
rect 254898 27978 255518 28046
rect 254898 27922 254994 27978
rect 255050 27922 255118 27978
rect 255174 27922 255242 27978
rect 255298 27922 255366 27978
rect 255422 27922 255518 27978
rect 254898 10350 255518 27922
rect 254898 10294 254994 10350
rect 255050 10294 255118 10350
rect 255174 10294 255242 10350
rect 255298 10294 255366 10350
rect 255422 10294 255518 10350
rect 254898 10226 255518 10294
rect 254898 10170 254994 10226
rect 255050 10170 255118 10226
rect 255174 10170 255242 10226
rect 255298 10170 255366 10226
rect 255422 10170 255518 10226
rect 254898 10102 255518 10170
rect 254898 10046 254994 10102
rect 255050 10046 255118 10102
rect 255174 10046 255242 10102
rect 255298 10046 255366 10102
rect 255422 10046 255518 10102
rect 254898 9978 255518 10046
rect 254898 9922 254994 9978
rect 255050 9922 255118 9978
rect 255174 9922 255242 9978
rect 255298 9922 255366 9978
rect 255422 9922 255518 9978
rect 254898 -1120 255518 9922
rect 254898 -1176 254994 -1120
rect 255050 -1176 255118 -1120
rect 255174 -1176 255242 -1120
rect 255298 -1176 255366 -1120
rect 255422 -1176 255518 -1120
rect 254898 -1244 255518 -1176
rect 254898 -1300 254994 -1244
rect 255050 -1300 255118 -1244
rect 255174 -1300 255242 -1244
rect 255298 -1300 255366 -1244
rect 255422 -1300 255518 -1244
rect 254898 -1368 255518 -1300
rect 254898 -1424 254994 -1368
rect 255050 -1424 255118 -1368
rect 255174 -1424 255242 -1368
rect 255298 -1424 255366 -1368
rect 255422 -1424 255518 -1368
rect 254898 -1492 255518 -1424
rect 254898 -1548 254994 -1492
rect 255050 -1548 255118 -1492
rect 255174 -1548 255242 -1492
rect 255298 -1548 255366 -1492
rect 255422 -1548 255518 -1492
rect 254898 -1644 255518 -1548
rect 281898 22350 282518 39922
rect 281898 22294 281994 22350
rect 282050 22294 282118 22350
rect 282174 22294 282242 22350
rect 282298 22294 282366 22350
rect 282422 22294 282518 22350
rect 281898 22226 282518 22294
rect 281898 22170 281994 22226
rect 282050 22170 282118 22226
rect 282174 22170 282242 22226
rect 282298 22170 282366 22226
rect 282422 22170 282518 22226
rect 281898 22102 282518 22170
rect 281898 22046 281994 22102
rect 282050 22046 282118 22102
rect 282174 22046 282242 22102
rect 282298 22046 282366 22102
rect 282422 22046 282518 22102
rect 281898 21978 282518 22046
rect 281898 21922 281994 21978
rect 282050 21922 282118 21978
rect 282174 21922 282242 21978
rect 282298 21922 282366 21978
rect 282422 21922 282518 21978
rect 281898 4350 282518 21922
rect 281898 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 282518 4350
rect 281898 4226 282518 4294
rect 281898 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 282518 4226
rect 281898 4102 282518 4170
rect 281898 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 282518 4102
rect 281898 3978 282518 4046
rect 281898 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 282518 3978
rect 281898 -160 282518 3922
rect 281898 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 282518 -160
rect 281898 -284 282518 -216
rect 281898 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 282518 -284
rect 281898 -408 282518 -340
rect 281898 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 282518 -408
rect 281898 -532 282518 -464
rect 281898 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 282518 -532
rect 281898 -1644 282518 -588
rect 285618 244350 286238 257490
rect 312618 256350 313238 257490
rect 312618 256294 312714 256350
rect 312770 256294 312838 256350
rect 312894 256294 312962 256350
rect 313018 256294 313086 256350
rect 313142 256294 313238 256350
rect 312618 256226 313238 256294
rect 312618 256170 312714 256226
rect 312770 256170 312838 256226
rect 312894 256170 312962 256226
rect 313018 256170 313086 256226
rect 313142 256170 313238 256226
rect 312618 256102 313238 256170
rect 312618 256046 312714 256102
rect 312770 256046 312838 256102
rect 312894 256046 312962 256102
rect 313018 256046 313086 256102
rect 313142 256046 313238 256102
rect 312618 255978 313238 256046
rect 312618 255922 312714 255978
rect 312770 255922 312838 255978
rect 312894 255922 312962 255978
rect 313018 255922 313086 255978
rect 313142 255922 313238 255978
rect 285618 244294 285714 244350
rect 285770 244294 285838 244350
rect 285894 244294 285962 244350
rect 286018 244294 286086 244350
rect 286142 244294 286238 244350
rect 285618 244226 286238 244294
rect 285618 244170 285714 244226
rect 285770 244170 285838 244226
rect 285894 244170 285962 244226
rect 286018 244170 286086 244226
rect 286142 244170 286238 244226
rect 285618 244102 286238 244170
rect 285618 244046 285714 244102
rect 285770 244046 285838 244102
rect 285894 244046 285962 244102
rect 286018 244046 286086 244102
rect 286142 244046 286238 244102
rect 285618 243978 286238 244046
rect 285618 243922 285714 243978
rect 285770 243922 285838 243978
rect 285894 243922 285962 243978
rect 286018 243922 286086 243978
rect 286142 243922 286238 243978
rect 285618 226350 286238 243922
rect 285618 226294 285714 226350
rect 285770 226294 285838 226350
rect 285894 226294 285962 226350
rect 286018 226294 286086 226350
rect 286142 226294 286238 226350
rect 285618 226226 286238 226294
rect 285618 226170 285714 226226
rect 285770 226170 285838 226226
rect 285894 226170 285962 226226
rect 286018 226170 286086 226226
rect 286142 226170 286238 226226
rect 285618 226102 286238 226170
rect 285618 226046 285714 226102
rect 285770 226046 285838 226102
rect 285894 226046 285962 226102
rect 286018 226046 286086 226102
rect 286142 226046 286238 226102
rect 285618 225978 286238 226046
rect 285618 225922 285714 225978
rect 285770 225922 285838 225978
rect 285894 225922 285962 225978
rect 286018 225922 286086 225978
rect 286142 225922 286238 225978
rect 285618 208350 286238 225922
rect 285618 208294 285714 208350
rect 285770 208294 285838 208350
rect 285894 208294 285962 208350
rect 286018 208294 286086 208350
rect 286142 208294 286238 208350
rect 285618 208226 286238 208294
rect 285618 208170 285714 208226
rect 285770 208170 285838 208226
rect 285894 208170 285962 208226
rect 286018 208170 286086 208226
rect 286142 208170 286238 208226
rect 285618 208102 286238 208170
rect 285618 208046 285714 208102
rect 285770 208046 285838 208102
rect 285894 208046 285962 208102
rect 286018 208046 286086 208102
rect 286142 208046 286238 208102
rect 285618 207978 286238 208046
rect 285618 207922 285714 207978
rect 285770 207922 285838 207978
rect 285894 207922 285962 207978
rect 286018 207922 286086 207978
rect 286142 207922 286238 207978
rect 285618 190350 286238 207922
rect 285618 190294 285714 190350
rect 285770 190294 285838 190350
rect 285894 190294 285962 190350
rect 286018 190294 286086 190350
rect 286142 190294 286238 190350
rect 285618 190226 286238 190294
rect 285618 190170 285714 190226
rect 285770 190170 285838 190226
rect 285894 190170 285962 190226
rect 286018 190170 286086 190226
rect 286142 190170 286238 190226
rect 285618 190102 286238 190170
rect 285618 190046 285714 190102
rect 285770 190046 285838 190102
rect 285894 190046 285962 190102
rect 286018 190046 286086 190102
rect 286142 190046 286238 190102
rect 285618 189978 286238 190046
rect 285618 189922 285714 189978
rect 285770 189922 285838 189978
rect 285894 189922 285962 189978
rect 286018 189922 286086 189978
rect 286142 189922 286238 189978
rect 285618 172350 286238 189922
rect 285618 172294 285714 172350
rect 285770 172294 285838 172350
rect 285894 172294 285962 172350
rect 286018 172294 286086 172350
rect 286142 172294 286238 172350
rect 285618 172226 286238 172294
rect 285618 172170 285714 172226
rect 285770 172170 285838 172226
rect 285894 172170 285962 172226
rect 286018 172170 286086 172226
rect 286142 172170 286238 172226
rect 285618 172102 286238 172170
rect 285618 172046 285714 172102
rect 285770 172046 285838 172102
rect 285894 172046 285962 172102
rect 286018 172046 286086 172102
rect 286142 172046 286238 172102
rect 285618 171978 286238 172046
rect 285618 171922 285714 171978
rect 285770 171922 285838 171978
rect 285894 171922 285962 171978
rect 286018 171922 286086 171978
rect 286142 171922 286238 171978
rect 285618 154350 286238 171922
rect 285618 154294 285714 154350
rect 285770 154294 285838 154350
rect 285894 154294 285962 154350
rect 286018 154294 286086 154350
rect 286142 154294 286238 154350
rect 285618 154226 286238 154294
rect 285618 154170 285714 154226
rect 285770 154170 285838 154226
rect 285894 154170 285962 154226
rect 286018 154170 286086 154226
rect 286142 154170 286238 154226
rect 285618 154102 286238 154170
rect 285618 154046 285714 154102
rect 285770 154046 285838 154102
rect 285894 154046 285962 154102
rect 286018 154046 286086 154102
rect 286142 154046 286238 154102
rect 285618 153978 286238 154046
rect 285618 153922 285714 153978
rect 285770 153922 285838 153978
rect 285894 153922 285962 153978
rect 286018 153922 286086 153978
rect 286142 153922 286238 153978
rect 285618 136350 286238 153922
rect 285618 136294 285714 136350
rect 285770 136294 285838 136350
rect 285894 136294 285962 136350
rect 286018 136294 286086 136350
rect 286142 136294 286238 136350
rect 285618 136226 286238 136294
rect 285618 136170 285714 136226
rect 285770 136170 285838 136226
rect 285894 136170 285962 136226
rect 286018 136170 286086 136226
rect 286142 136170 286238 136226
rect 285618 136102 286238 136170
rect 285618 136046 285714 136102
rect 285770 136046 285838 136102
rect 285894 136046 285962 136102
rect 286018 136046 286086 136102
rect 286142 136046 286238 136102
rect 285618 135978 286238 136046
rect 285618 135922 285714 135978
rect 285770 135922 285838 135978
rect 285894 135922 285962 135978
rect 286018 135922 286086 135978
rect 286142 135922 286238 135978
rect 285618 118350 286238 135922
rect 285618 118294 285714 118350
rect 285770 118294 285838 118350
rect 285894 118294 285962 118350
rect 286018 118294 286086 118350
rect 286142 118294 286238 118350
rect 285618 118226 286238 118294
rect 285618 118170 285714 118226
rect 285770 118170 285838 118226
rect 285894 118170 285962 118226
rect 286018 118170 286086 118226
rect 286142 118170 286238 118226
rect 285618 118102 286238 118170
rect 285618 118046 285714 118102
rect 285770 118046 285838 118102
rect 285894 118046 285962 118102
rect 286018 118046 286086 118102
rect 286142 118046 286238 118102
rect 285618 117978 286238 118046
rect 285618 117922 285714 117978
rect 285770 117922 285838 117978
rect 285894 117922 285962 117978
rect 286018 117922 286086 117978
rect 286142 117922 286238 117978
rect 285618 100350 286238 117922
rect 285618 100294 285714 100350
rect 285770 100294 285838 100350
rect 285894 100294 285962 100350
rect 286018 100294 286086 100350
rect 286142 100294 286238 100350
rect 285618 100226 286238 100294
rect 285618 100170 285714 100226
rect 285770 100170 285838 100226
rect 285894 100170 285962 100226
rect 286018 100170 286086 100226
rect 286142 100170 286238 100226
rect 285618 100102 286238 100170
rect 285618 100046 285714 100102
rect 285770 100046 285838 100102
rect 285894 100046 285962 100102
rect 286018 100046 286086 100102
rect 286142 100046 286238 100102
rect 285618 99978 286238 100046
rect 285618 99922 285714 99978
rect 285770 99922 285838 99978
rect 285894 99922 285962 99978
rect 286018 99922 286086 99978
rect 286142 99922 286238 99978
rect 285618 82350 286238 99922
rect 285618 82294 285714 82350
rect 285770 82294 285838 82350
rect 285894 82294 285962 82350
rect 286018 82294 286086 82350
rect 286142 82294 286238 82350
rect 285618 82226 286238 82294
rect 285618 82170 285714 82226
rect 285770 82170 285838 82226
rect 285894 82170 285962 82226
rect 286018 82170 286086 82226
rect 286142 82170 286238 82226
rect 285618 82102 286238 82170
rect 285618 82046 285714 82102
rect 285770 82046 285838 82102
rect 285894 82046 285962 82102
rect 286018 82046 286086 82102
rect 286142 82046 286238 82102
rect 285618 81978 286238 82046
rect 285618 81922 285714 81978
rect 285770 81922 285838 81978
rect 285894 81922 285962 81978
rect 286018 81922 286086 81978
rect 286142 81922 286238 81978
rect 285618 64350 286238 81922
rect 285618 64294 285714 64350
rect 285770 64294 285838 64350
rect 285894 64294 285962 64350
rect 286018 64294 286086 64350
rect 286142 64294 286238 64350
rect 285618 64226 286238 64294
rect 285618 64170 285714 64226
rect 285770 64170 285838 64226
rect 285894 64170 285962 64226
rect 286018 64170 286086 64226
rect 286142 64170 286238 64226
rect 285618 64102 286238 64170
rect 285618 64046 285714 64102
rect 285770 64046 285838 64102
rect 285894 64046 285962 64102
rect 286018 64046 286086 64102
rect 286142 64046 286238 64102
rect 285618 63978 286238 64046
rect 285618 63922 285714 63978
rect 285770 63922 285838 63978
rect 285894 63922 285962 63978
rect 286018 63922 286086 63978
rect 286142 63922 286238 63978
rect 285618 46350 286238 63922
rect 285618 46294 285714 46350
rect 285770 46294 285838 46350
rect 285894 46294 285962 46350
rect 286018 46294 286086 46350
rect 286142 46294 286238 46350
rect 285618 46226 286238 46294
rect 285618 46170 285714 46226
rect 285770 46170 285838 46226
rect 285894 46170 285962 46226
rect 286018 46170 286086 46226
rect 286142 46170 286238 46226
rect 285618 46102 286238 46170
rect 285618 46046 285714 46102
rect 285770 46046 285838 46102
rect 285894 46046 285962 46102
rect 286018 46046 286086 46102
rect 286142 46046 286238 46102
rect 285618 45978 286238 46046
rect 285618 45922 285714 45978
rect 285770 45922 285838 45978
rect 285894 45922 285962 45978
rect 286018 45922 286086 45978
rect 286142 45922 286238 45978
rect 285618 28350 286238 45922
rect 285618 28294 285714 28350
rect 285770 28294 285838 28350
rect 285894 28294 285962 28350
rect 286018 28294 286086 28350
rect 286142 28294 286238 28350
rect 285618 28226 286238 28294
rect 285618 28170 285714 28226
rect 285770 28170 285838 28226
rect 285894 28170 285962 28226
rect 286018 28170 286086 28226
rect 286142 28170 286238 28226
rect 285618 28102 286238 28170
rect 285618 28046 285714 28102
rect 285770 28046 285838 28102
rect 285894 28046 285962 28102
rect 286018 28046 286086 28102
rect 286142 28046 286238 28102
rect 285618 27978 286238 28046
rect 285618 27922 285714 27978
rect 285770 27922 285838 27978
rect 285894 27922 285962 27978
rect 286018 27922 286086 27978
rect 286142 27922 286238 27978
rect 285618 10350 286238 27922
rect 285618 10294 285714 10350
rect 285770 10294 285838 10350
rect 285894 10294 285962 10350
rect 286018 10294 286086 10350
rect 286142 10294 286238 10350
rect 285618 10226 286238 10294
rect 285618 10170 285714 10226
rect 285770 10170 285838 10226
rect 285894 10170 285962 10226
rect 286018 10170 286086 10226
rect 286142 10170 286238 10226
rect 285618 10102 286238 10170
rect 285618 10046 285714 10102
rect 285770 10046 285838 10102
rect 285894 10046 285962 10102
rect 286018 10046 286086 10102
rect 286142 10046 286238 10102
rect 285618 9978 286238 10046
rect 285618 9922 285714 9978
rect 285770 9922 285838 9978
rect 285894 9922 285962 9978
rect 286018 9922 286086 9978
rect 286142 9922 286238 9978
rect 285618 -1120 286238 9922
rect 291452 252084 291508 252094
rect 291452 6020 291508 252028
rect 312618 238350 313238 255922
rect 312618 238294 312714 238350
rect 312770 238294 312838 238350
rect 312894 238294 312962 238350
rect 313018 238294 313086 238350
rect 313142 238294 313238 238350
rect 312618 238226 313238 238294
rect 312618 238170 312714 238226
rect 312770 238170 312838 238226
rect 312894 238170 312962 238226
rect 313018 238170 313086 238226
rect 313142 238170 313238 238226
rect 312618 238102 313238 238170
rect 312618 238046 312714 238102
rect 312770 238046 312838 238102
rect 312894 238046 312962 238102
rect 313018 238046 313086 238102
rect 313142 238046 313238 238102
rect 312618 237978 313238 238046
rect 312618 237922 312714 237978
rect 312770 237922 312838 237978
rect 312894 237922 312962 237978
rect 313018 237922 313086 237978
rect 313142 237922 313238 237978
rect 312618 220350 313238 237922
rect 312618 220294 312714 220350
rect 312770 220294 312838 220350
rect 312894 220294 312962 220350
rect 313018 220294 313086 220350
rect 313142 220294 313238 220350
rect 312618 220226 313238 220294
rect 312618 220170 312714 220226
rect 312770 220170 312838 220226
rect 312894 220170 312962 220226
rect 313018 220170 313086 220226
rect 313142 220170 313238 220226
rect 312618 220102 313238 220170
rect 312618 220046 312714 220102
rect 312770 220046 312838 220102
rect 312894 220046 312962 220102
rect 313018 220046 313086 220102
rect 313142 220046 313238 220102
rect 312618 219978 313238 220046
rect 312618 219922 312714 219978
rect 312770 219922 312838 219978
rect 312894 219922 312962 219978
rect 313018 219922 313086 219978
rect 313142 219922 313238 219978
rect 307468 212884 307524 212894
rect 291564 211078 291620 211088
rect 291564 154308 291620 211022
rect 291564 105140 291620 154252
rect 296492 210898 296548 210908
rect 296492 156660 296548 210842
rect 296492 108052 296548 156604
rect 296492 107986 296548 107996
rect 291564 105074 291620 105084
rect 299500 82147 299820 82204
rect 299500 82091 299528 82147
rect 299584 82091 299632 82147
rect 299688 82091 299736 82147
rect 299792 82091 299820 82147
rect 299500 82043 299820 82091
rect 299500 81987 299528 82043
rect 299584 81987 299632 82043
rect 299688 81987 299736 82043
rect 299792 81987 299820 82043
rect 299500 81939 299820 81987
rect 299500 81883 299528 81939
rect 299584 81883 299632 81939
rect 299688 81883 299736 81939
rect 299792 81883 299820 81939
rect 299500 81826 299820 81883
rect 295342 76350 295662 76384
rect 295342 76294 295412 76350
rect 295468 76294 295536 76350
rect 295592 76294 295662 76350
rect 295342 76226 295662 76294
rect 295342 76170 295412 76226
rect 295468 76170 295536 76226
rect 295592 76170 295662 76226
rect 295342 76102 295662 76170
rect 295342 76046 295412 76102
rect 295468 76046 295536 76102
rect 295592 76046 295662 76102
rect 295342 75978 295662 76046
rect 295342 75922 295412 75978
rect 295468 75922 295536 75978
rect 295592 75922 295662 75978
rect 295342 75888 295662 75922
rect 303658 76350 303978 76384
rect 303658 76294 303728 76350
rect 303784 76294 303852 76350
rect 303908 76294 303978 76350
rect 303658 76226 303978 76294
rect 303658 76170 303728 76226
rect 303784 76170 303852 76226
rect 303908 76170 303978 76226
rect 303658 76102 303978 76170
rect 303658 76046 303728 76102
rect 303784 76046 303852 76102
rect 303908 76046 303978 76102
rect 303658 75978 303978 76046
rect 303658 75922 303728 75978
rect 303784 75922 303852 75978
rect 303908 75922 303978 75978
rect 303658 75888 303978 75922
rect 299500 64350 299820 64384
rect 299500 64294 299570 64350
rect 299626 64294 299694 64350
rect 299750 64294 299820 64350
rect 299500 64226 299820 64294
rect 299500 64170 299570 64226
rect 299626 64170 299694 64226
rect 299750 64170 299820 64226
rect 299500 64102 299820 64170
rect 299500 64046 299570 64102
rect 299626 64046 299694 64102
rect 299750 64046 299820 64102
rect 299500 63978 299820 64046
rect 299500 63922 299570 63978
rect 299626 63922 299694 63978
rect 299750 63922 299820 63978
rect 299500 63888 299820 63922
rect 295342 58350 295662 58384
rect 295342 58294 295412 58350
rect 295468 58294 295536 58350
rect 295592 58294 295662 58350
rect 295342 58226 295662 58294
rect 295342 58170 295412 58226
rect 295468 58170 295536 58226
rect 295592 58170 295662 58226
rect 295342 58102 295662 58170
rect 295342 58046 295412 58102
rect 295468 58046 295536 58102
rect 295592 58046 295662 58102
rect 295342 57978 295662 58046
rect 295342 57922 295412 57978
rect 295468 57922 295536 57978
rect 295592 57922 295662 57978
rect 295342 57888 295662 57922
rect 303658 58350 303978 58384
rect 303658 58294 303728 58350
rect 303784 58294 303852 58350
rect 303908 58294 303978 58350
rect 303658 58226 303978 58294
rect 303658 58170 303728 58226
rect 303784 58170 303852 58226
rect 303908 58170 303978 58226
rect 303658 58102 303978 58170
rect 303658 58046 303728 58102
rect 303784 58046 303852 58102
rect 303908 58046 303978 58102
rect 303658 57978 303978 58046
rect 303658 57922 303728 57978
rect 303784 57922 303852 57978
rect 303908 57922 303978 57978
rect 303658 57888 303978 57922
rect 307468 50260 307524 212828
rect 312618 202350 313238 219922
rect 316338 244350 316958 257490
rect 316338 244294 316434 244350
rect 316490 244294 316558 244350
rect 316614 244294 316682 244350
rect 316738 244294 316806 244350
rect 316862 244294 316958 244350
rect 316338 244226 316958 244294
rect 316338 244170 316434 244226
rect 316490 244170 316558 244226
rect 316614 244170 316682 244226
rect 316738 244170 316806 244226
rect 316862 244170 316958 244226
rect 316338 244102 316958 244170
rect 316338 244046 316434 244102
rect 316490 244046 316558 244102
rect 316614 244046 316682 244102
rect 316738 244046 316806 244102
rect 316862 244046 316958 244102
rect 316338 243978 316958 244046
rect 316338 243922 316434 243978
rect 316490 243922 316558 243978
rect 316614 243922 316682 243978
rect 316738 243922 316806 243978
rect 316862 243922 316958 243978
rect 316338 226350 316958 243922
rect 316338 226294 316434 226350
rect 316490 226294 316558 226350
rect 316614 226294 316682 226350
rect 316738 226294 316806 226350
rect 316862 226294 316958 226350
rect 316338 226226 316958 226294
rect 316338 226170 316434 226226
rect 316490 226170 316558 226226
rect 316614 226170 316682 226226
rect 316738 226170 316806 226226
rect 316862 226170 316958 226226
rect 316338 226102 316958 226170
rect 316338 226046 316434 226102
rect 316490 226046 316558 226102
rect 316614 226046 316682 226102
rect 316738 226046 316806 226102
rect 316862 226046 316958 226102
rect 316338 225978 316958 226046
rect 316338 225922 316434 225978
rect 316490 225922 316558 225978
rect 316614 225922 316682 225978
rect 316738 225922 316806 225978
rect 316862 225922 316958 225978
rect 312618 202294 312714 202350
rect 312770 202294 312838 202350
rect 312894 202294 312962 202350
rect 313018 202294 313086 202350
rect 313142 202294 313238 202350
rect 312618 202226 313238 202294
rect 312618 202170 312714 202226
rect 312770 202170 312838 202226
rect 312894 202170 312962 202226
rect 313018 202170 313086 202226
rect 313142 202170 313238 202226
rect 312618 202102 313238 202170
rect 312618 202046 312714 202102
rect 312770 202046 312838 202102
rect 312894 202046 312962 202102
rect 313018 202046 313086 202102
rect 313142 202046 313238 202102
rect 312618 201978 313238 202046
rect 312618 201922 312714 201978
rect 312770 201922 312838 201978
rect 312894 201922 312962 201978
rect 313018 201922 313086 201978
rect 313142 201922 313238 201978
rect 312618 184350 313238 201922
rect 312618 184294 312714 184350
rect 312770 184294 312838 184350
rect 312894 184294 312962 184350
rect 313018 184294 313086 184350
rect 313142 184294 313238 184350
rect 312618 184226 313238 184294
rect 312618 184170 312714 184226
rect 312770 184170 312838 184226
rect 312894 184170 312962 184226
rect 313018 184170 313086 184226
rect 313142 184170 313238 184226
rect 312618 184102 313238 184170
rect 312618 184046 312714 184102
rect 312770 184046 312838 184102
rect 312894 184046 312962 184102
rect 313018 184046 313086 184102
rect 313142 184046 313238 184102
rect 312618 183978 313238 184046
rect 312618 183922 312714 183978
rect 312770 183922 312838 183978
rect 312894 183922 312962 183978
rect 313018 183922 313086 183978
rect 313142 183922 313238 183978
rect 312618 166350 313238 183922
rect 312618 166294 312714 166350
rect 312770 166294 312838 166350
rect 312894 166294 312962 166350
rect 313018 166294 313086 166350
rect 313142 166294 313238 166350
rect 312618 166226 313238 166294
rect 312618 166170 312714 166226
rect 312770 166170 312838 166226
rect 312894 166170 312962 166226
rect 313018 166170 313086 166226
rect 313142 166170 313238 166226
rect 312618 166102 313238 166170
rect 312618 166046 312714 166102
rect 312770 166046 312838 166102
rect 312894 166046 312962 166102
rect 313018 166046 313086 166102
rect 313142 166046 313238 166102
rect 312618 165978 313238 166046
rect 312618 165922 312714 165978
rect 312770 165922 312838 165978
rect 312894 165922 312962 165978
rect 313018 165922 313086 165978
rect 313142 165922 313238 165978
rect 312618 148350 313238 165922
rect 314188 212772 314244 212782
rect 312618 148294 312714 148350
rect 312770 148294 312838 148350
rect 312894 148294 312962 148350
rect 313018 148294 313086 148350
rect 313142 148294 313238 148350
rect 312618 148226 313238 148294
rect 312618 148170 312714 148226
rect 312770 148170 312838 148226
rect 312894 148170 312962 148226
rect 313018 148170 313086 148226
rect 313142 148170 313238 148226
rect 312618 148102 313238 148170
rect 312618 148046 312714 148102
rect 312770 148046 312838 148102
rect 312894 148046 312962 148102
rect 313018 148046 313086 148102
rect 313142 148046 313238 148102
rect 312618 147978 313238 148046
rect 312618 147922 312714 147978
rect 312770 147922 312838 147978
rect 312894 147922 312962 147978
rect 313018 147922 313086 147978
rect 313142 147922 313238 147978
rect 312618 130350 313238 147922
rect 312618 130294 312714 130350
rect 312770 130294 312838 130350
rect 312894 130294 312962 130350
rect 313018 130294 313086 130350
rect 313142 130294 313238 130350
rect 312618 130226 313238 130294
rect 312618 130170 312714 130226
rect 312770 130170 312838 130226
rect 312894 130170 312962 130226
rect 313018 130170 313086 130226
rect 313142 130170 313238 130226
rect 312618 130102 313238 130170
rect 312618 130046 312714 130102
rect 312770 130046 312838 130102
rect 312894 130046 312962 130102
rect 313018 130046 313086 130102
rect 313142 130046 313238 130102
rect 312618 129978 313238 130046
rect 312618 129922 312714 129978
rect 312770 129922 312838 129978
rect 312894 129922 312962 129978
rect 313018 129922 313086 129978
rect 313142 129922 313238 129978
rect 312618 112350 313238 129922
rect 313404 153658 313460 153668
rect 313404 116788 313460 153602
rect 313404 116722 313460 116732
rect 312618 112294 312714 112350
rect 312770 112294 312838 112350
rect 312894 112294 312962 112350
rect 313018 112294 313086 112350
rect 313142 112294 313238 112350
rect 312618 112226 313238 112294
rect 312618 112170 312714 112226
rect 312770 112170 312838 112226
rect 312894 112170 312962 112226
rect 313018 112170 313086 112226
rect 313142 112170 313238 112226
rect 312618 112102 313238 112170
rect 312618 112046 312714 112102
rect 312770 112046 312838 112102
rect 312894 112046 312962 112102
rect 313018 112046 313086 112102
rect 313142 112046 313238 112102
rect 312618 111978 313238 112046
rect 312618 111922 312714 111978
rect 312770 111922 312838 111978
rect 312894 111922 312962 111978
rect 313018 111922 313086 111978
rect 313142 111922 313238 111978
rect 312618 94350 313238 111922
rect 312618 94294 312714 94350
rect 312770 94294 312838 94350
rect 312894 94294 312962 94350
rect 313018 94294 313086 94350
rect 313142 94294 313238 94350
rect 312618 94226 313238 94294
rect 312618 94170 312714 94226
rect 312770 94170 312838 94226
rect 312894 94170 312962 94226
rect 313018 94170 313086 94226
rect 313142 94170 313238 94226
rect 312618 94102 313238 94170
rect 312618 94046 312714 94102
rect 312770 94046 312838 94102
rect 312894 94046 312962 94102
rect 313018 94046 313086 94102
rect 313142 94046 313238 94102
rect 312618 93978 313238 94046
rect 312618 93922 312714 93978
rect 312770 93922 312838 93978
rect 312894 93922 312962 93978
rect 313018 93922 313086 93978
rect 313142 93922 313238 93978
rect 307816 82147 308136 82204
rect 307816 82091 307844 82147
rect 307900 82091 307948 82147
rect 308004 82091 308052 82147
rect 308108 82091 308136 82147
rect 307816 82043 308136 82091
rect 307816 81987 307844 82043
rect 307900 81987 307948 82043
rect 308004 81987 308052 82043
rect 308108 81987 308136 82043
rect 307816 81939 308136 81987
rect 307816 81883 307844 81939
rect 307900 81883 307948 81939
rect 308004 81883 308052 81939
rect 308108 81883 308136 81939
rect 307816 81826 308136 81883
rect 311974 76350 312294 76384
rect 311974 76294 312044 76350
rect 312100 76294 312168 76350
rect 312224 76294 312294 76350
rect 311974 76226 312294 76294
rect 311974 76170 312044 76226
rect 312100 76170 312168 76226
rect 312224 76170 312294 76226
rect 311974 76102 312294 76170
rect 311974 76046 312044 76102
rect 312100 76046 312168 76102
rect 312224 76046 312294 76102
rect 311974 75978 312294 76046
rect 311974 75922 312044 75978
rect 312100 75922 312168 75978
rect 312224 75922 312294 75978
rect 311974 75888 312294 75922
rect 312618 76350 313238 93922
rect 312618 76294 312714 76350
rect 312770 76294 312838 76350
rect 312894 76294 312962 76350
rect 313018 76294 313086 76350
rect 313142 76294 313238 76350
rect 312618 76226 313238 76294
rect 312618 76170 312714 76226
rect 312770 76170 312838 76226
rect 312894 76170 312962 76226
rect 313018 76170 313086 76226
rect 313142 76170 313238 76226
rect 312618 76102 313238 76170
rect 312618 76046 312714 76102
rect 312770 76046 312838 76102
rect 312894 76046 312962 76102
rect 313018 76046 313086 76102
rect 313142 76046 313238 76102
rect 312618 75978 313238 76046
rect 312618 75922 312714 75978
rect 312770 75922 312838 75978
rect 312894 75922 312962 75978
rect 313018 75922 313086 75978
rect 313142 75922 313238 75978
rect 307816 64350 308136 64384
rect 307816 64294 307886 64350
rect 307942 64294 308010 64350
rect 308066 64294 308136 64350
rect 307816 64226 308136 64294
rect 307816 64170 307886 64226
rect 307942 64170 308010 64226
rect 308066 64170 308136 64226
rect 307816 64102 308136 64170
rect 307816 64046 307886 64102
rect 307942 64046 308010 64102
rect 308066 64046 308136 64102
rect 307816 63978 308136 64046
rect 307816 63922 307886 63978
rect 307942 63922 308010 63978
rect 308066 63922 308136 63978
rect 307816 63888 308136 63922
rect 311974 58350 312294 58384
rect 311974 58294 312044 58350
rect 312100 58294 312168 58350
rect 312224 58294 312294 58350
rect 311974 58226 312294 58294
rect 311974 58170 312044 58226
rect 312100 58170 312168 58226
rect 312224 58170 312294 58226
rect 311974 58102 312294 58170
rect 311974 58046 312044 58102
rect 312100 58046 312168 58102
rect 312224 58046 312294 58102
rect 311974 57978 312294 58046
rect 311974 57922 312044 57978
rect 312100 57922 312168 57978
rect 312224 57922 312294 57978
rect 311974 57888 312294 57922
rect 312618 58350 313238 75922
rect 312618 58294 312714 58350
rect 312770 58294 312838 58350
rect 312894 58294 312962 58350
rect 313018 58294 313086 58350
rect 313142 58294 313238 58350
rect 312618 58226 313238 58294
rect 312618 58170 312714 58226
rect 312770 58170 312838 58226
rect 312894 58170 312962 58226
rect 313018 58170 313086 58226
rect 313142 58170 313238 58226
rect 312618 58102 313238 58170
rect 312618 58046 312714 58102
rect 312770 58046 312838 58102
rect 312894 58046 312962 58102
rect 313018 58046 313086 58102
rect 313142 58046 313238 58102
rect 312618 57978 313238 58046
rect 312618 57922 312714 57978
rect 312770 57922 312838 57978
rect 312894 57922 312962 57978
rect 313018 57922 313086 57978
rect 313142 57922 313238 57978
rect 307468 50194 307524 50204
rect 291452 5954 291508 5964
rect 312618 40350 313238 57922
rect 314188 50260 314244 212716
rect 316338 208350 316958 225922
rect 343338 256350 343958 257490
rect 343338 256294 343434 256350
rect 343490 256294 343558 256350
rect 343614 256294 343682 256350
rect 343738 256294 343806 256350
rect 343862 256294 343958 256350
rect 343338 256226 343958 256294
rect 343338 256170 343434 256226
rect 343490 256170 343558 256226
rect 343614 256170 343682 256226
rect 343738 256170 343806 256226
rect 343862 256170 343958 256226
rect 343338 256102 343958 256170
rect 343338 256046 343434 256102
rect 343490 256046 343558 256102
rect 343614 256046 343682 256102
rect 343738 256046 343806 256102
rect 343862 256046 343958 256102
rect 343338 255978 343958 256046
rect 343338 255922 343434 255978
rect 343490 255922 343558 255978
rect 343614 255922 343682 255978
rect 343738 255922 343806 255978
rect 343862 255922 343958 255978
rect 343338 238350 343958 255922
rect 343338 238294 343434 238350
rect 343490 238294 343558 238350
rect 343614 238294 343682 238350
rect 343738 238294 343806 238350
rect 343862 238294 343958 238350
rect 343338 238226 343958 238294
rect 343338 238170 343434 238226
rect 343490 238170 343558 238226
rect 343614 238170 343682 238226
rect 343738 238170 343806 238226
rect 343862 238170 343958 238226
rect 343338 238102 343958 238170
rect 343338 238046 343434 238102
rect 343490 238046 343558 238102
rect 343614 238046 343682 238102
rect 343738 238046 343806 238102
rect 343862 238046 343958 238102
rect 343338 237978 343958 238046
rect 343338 237922 343434 237978
rect 343490 237922 343558 237978
rect 343614 237922 343682 237978
rect 343738 237922 343806 237978
rect 343862 237922 343958 237978
rect 343338 220350 343958 237922
rect 343338 220294 343434 220350
rect 343490 220294 343558 220350
rect 343614 220294 343682 220350
rect 343738 220294 343806 220350
rect 343862 220294 343958 220350
rect 343338 220226 343958 220294
rect 343338 220170 343434 220226
rect 343490 220170 343558 220226
rect 343614 220170 343682 220226
rect 343738 220170 343806 220226
rect 343862 220170 343958 220226
rect 343338 220102 343958 220170
rect 343338 220046 343434 220102
rect 343490 220046 343558 220102
rect 343614 220046 343682 220102
rect 343738 220046 343806 220102
rect 343862 220046 343958 220102
rect 343338 219978 343958 220046
rect 343338 219922 343434 219978
rect 343490 219922 343558 219978
rect 343614 219922 343682 219978
rect 343738 219922 343806 219978
rect 343862 219922 343958 219978
rect 316338 208294 316434 208350
rect 316490 208294 316558 208350
rect 316614 208294 316682 208350
rect 316738 208294 316806 208350
rect 316862 208294 316958 208350
rect 316338 208226 316958 208294
rect 316338 208170 316434 208226
rect 316490 208170 316558 208226
rect 316614 208170 316682 208226
rect 316738 208170 316806 208226
rect 316862 208170 316958 208226
rect 316338 208102 316958 208170
rect 316338 208046 316434 208102
rect 316490 208046 316558 208102
rect 316614 208046 316682 208102
rect 316738 208046 316806 208102
rect 316862 208046 316958 208102
rect 316338 207978 316958 208046
rect 316338 207922 316434 207978
rect 316490 207922 316558 207978
rect 316614 207922 316682 207978
rect 316738 207922 316806 207978
rect 316862 207922 316958 207978
rect 316338 190350 316958 207922
rect 316338 190294 316434 190350
rect 316490 190294 316558 190350
rect 316614 190294 316682 190350
rect 316738 190294 316806 190350
rect 316862 190294 316958 190350
rect 316338 190226 316958 190294
rect 316338 190170 316434 190226
rect 316490 190170 316558 190226
rect 316614 190170 316682 190226
rect 316738 190170 316806 190226
rect 316862 190170 316958 190226
rect 316338 190102 316958 190170
rect 316338 190046 316434 190102
rect 316490 190046 316558 190102
rect 316614 190046 316682 190102
rect 316738 190046 316806 190102
rect 316862 190046 316958 190102
rect 316338 189978 316958 190046
rect 316338 189922 316434 189978
rect 316490 189922 316558 189978
rect 316614 189922 316682 189978
rect 316738 189922 316806 189978
rect 316862 189922 316958 189978
rect 316338 172350 316958 189922
rect 316338 172294 316434 172350
rect 316490 172294 316558 172350
rect 316614 172294 316682 172350
rect 316738 172294 316806 172350
rect 316862 172294 316958 172350
rect 316338 172226 316958 172294
rect 316338 172170 316434 172226
rect 316490 172170 316558 172226
rect 316614 172170 316682 172226
rect 316738 172170 316806 172226
rect 316862 172170 316958 172226
rect 316338 172102 316958 172170
rect 316338 172046 316434 172102
rect 316490 172046 316558 172102
rect 316614 172046 316682 172102
rect 316738 172046 316806 172102
rect 316862 172046 316958 172102
rect 316338 171978 316958 172046
rect 316338 171922 316434 171978
rect 316490 171922 316558 171978
rect 316614 171922 316682 171978
rect 316738 171922 316806 171978
rect 316862 171922 316958 171978
rect 316338 154350 316958 171922
rect 316338 154294 316434 154350
rect 316490 154294 316558 154350
rect 316614 154294 316682 154350
rect 316738 154294 316806 154350
rect 316862 154294 316958 154350
rect 316338 154226 316958 154294
rect 316338 154170 316434 154226
rect 316490 154170 316558 154226
rect 316614 154170 316682 154226
rect 316738 154170 316806 154226
rect 316862 154170 316958 154226
rect 316338 154102 316958 154170
rect 316338 154046 316434 154102
rect 316490 154046 316558 154102
rect 316614 154046 316682 154102
rect 316738 154046 316806 154102
rect 316862 154046 316958 154102
rect 316338 153978 316958 154046
rect 316338 153922 316434 153978
rect 316490 153922 316558 153978
rect 316614 153922 316682 153978
rect 316738 153922 316806 153978
rect 316862 153922 316958 153978
rect 316338 136350 316958 153922
rect 316338 136294 316434 136350
rect 316490 136294 316558 136350
rect 316614 136294 316682 136350
rect 316738 136294 316806 136350
rect 316862 136294 316958 136350
rect 316338 136226 316958 136294
rect 316338 136170 316434 136226
rect 316490 136170 316558 136226
rect 316614 136170 316682 136226
rect 316738 136170 316806 136226
rect 316862 136170 316958 136226
rect 316338 136102 316958 136170
rect 316338 136046 316434 136102
rect 316490 136046 316558 136102
rect 316614 136046 316682 136102
rect 316738 136046 316806 136102
rect 316862 136046 316958 136102
rect 316338 135978 316958 136046
rect 316338 135922 316434 135978
rect 316490 135922 316558 135978
rect 316614 135922 316682 135978
rect 316738 135922 316806 135978
rect 316862 135922 316958 135978
rect 316338 118350 316958 135922
rect 316338 118294 316434 118350
rect 316490 118294 316558 118350
rect 316614 118294 316682 118350
rect 316738 118294 316806 118350
rect 316862 118294 316958 118350
rect 316338 118226 316958 118294
rect 316338 118170 316434 118226
rect 316490 118170 316558 118226
rect 316614 118170 316682 118226
rect 316738 118170 316806 118226
rect 316862 118170 316958 118226
rect 316338 118102 316958 118170
rect 316338 118046 316434 118102
rect 316490 118046 316558 118102
rect 316614 118046 316682 118102
rect 316738 118046 316806 118102
rect 316862 118046 316958 118102
rect 316338 117978 316958 118046
rect 316338 117922 316434 117978
rect 316490 117922 316558 117978
rect 316614 117922 316682 117978
rect 316738 117922 316806 117978
rect 316862 117922 316958 117978
rect 316338 100350 316958 117922
rect 316338 100294 316434 100350
rect 316490 100294 316558 100350
rect 316614 100294 316682 100350
rect 316738 100294 316806 100350
rect 316862 100294 316958 100350
rect 316338 100226 316958 100294
rect 316338 100170 316434 100226
rect 316490 100170 316558 100226
rect 316614 100170 316682 100226
rect 316738 100170 316806 100226
rect 316862 100170 316958 100226
rect 316338 100102 316958 100170
rect 316338 100046 316434 100102
rect 316490 100046 316558 100102
rect 316614 100046 316682 100102
rect 316738 100046 316806 100102
rect 316862 100046 316958 100102
rect 316338 99978 316958 100046
rect 316338 99922 316434 99978
rect 316490 99922 316558 99978
rect 316614 99922 316682 99978
rect 316738 99922 316806 99978
rect 316862 99922 316958 99978
rect 316338 84316 316958 99922
rect 320908 212660 320964 212670
rect 316132 82147 316452 82204
rect 316132 82091 316160 82147
rect 316216 82091 316264 82147
rect 316320 82091 316368 82147
rect 316424 82091 316452 82147
rect 316132 82043 316452 82091
rect 316132 81987 316160 82043
rect 316216 81987 316264 82043
rect 316320 81987 316368 82043
rect 316424 81987 316452 82043
rect 316132 81939 316452 81987
rect 316132 81883 316160 81939
rect 316216 81883 316264 81939
rect 316320 81883 316368 81939
rect 316424 81883 316452 81939
rect 316132 81826 316452 81883
rect 320290 76350 320610 76384
rect 320290 76294 320360 76350
rect 320416 76294 320484 76350
rect 320540 76294 320610 76350
rect 320290 76226 320610 76294
rect 320290 76170 320360 76226
rect 320416 76170 320484 76226
rect 320540 76170 320610 76226
rect 320290 76102 320610 76170
rect 320290 76046 320360 76102
rect 320416 76046 320484 76102
rect 320540 76046 320610 76102
rect 320290 75978 320610 76046
rect 320290 75922 320360 75978
rect 320416 75922 320484 75978
rect 320540 75922 320610 75978
rect 320290 75888 320610 75922
rect 316132 64350 316452 64384
rect 316132 64294 316202 64350
rect 316258 64294 316326 64350
rect 316382 64294 316452 64350
rect 316132 64226 316452 64294
rect 316132 64170 316202 64226
rect 316258 64170 316326 64226
rect 316382 64170 316452 64226
rect 316132 64102 316452 64170
rect 316132 64046 316202 64102
rect 316258 64046 316326 64102
rect 316382 64046 316452 64102
rect 316132 63978 316452 64046
rect 316132 63922 316202 63978
rect 316258 63922 316326 63978
rect 316382 63922 316452 63978
rect 316132 63888 316452 63922
rect 320290 58350 320610 58384
rect 320290 58294 320360 58350
rect 320416 58294 320484 58350
rect 320540 58294 320610 58350
rect 320290 58226 320610 58294
rect 320290 58170 320360 58226
rect 320416 58170 320484 58226
rect 320540 58170 320610 58226
rect 320290 58102 320610 58170
rect 320290 58046 320360 58102
rect 320416 58046 320484 58102
rect 320540 58046 320610 58102
rect 320290 57978 320610 58046
rect 320290 57922 320360 57978
rect 320416 57922 320484 57978
rect 320540 57922 320610 57978
rect 320290 57888 320610 57922
rect 314188 50194 314244 50204
rect 312618 40294 312714 40350
rect 312770 40294 312838 40350
rect 312894 40294 312962 40350
rect 313018 40294 313086 40350
rect 313142 40294 313238 40350
rect 312618 40226 313238 40294
rect 312618 40170 312714 40226
rect 312770 40170 312838 40226
rect 312894 40170 312962 40226
rect 313018 40170 313086 40226
rect 313142 40170 313238 40226
rect 312618 40102 313238 40170
rect 312618 40046 312714 40102
rect 312770 40046 312838 40102
rect 312894 40046 312962 40102
rect 313018 40046 313086 40102
rect 313142 40046 313238 40102
rect 312618 39978 313238 40046
rect 312618 39922 312714 39978
rect 312770 39922 312838 39978
rect 312894 39922 312962 39978
rect 313018 39922 313086 39978
rect 313142 39922 313238 39978
rect 312618 22350 313238 39922
rect 312618 22294 312714 22350
rect 312770 22294 312838 22350
rect 312894 22294 312962 22350
rect 313018 22294 313086 22350
rect 313142 22294 313238 22350
rect 312618 22226 313238 22294
rect 312618 22170 312714 22226
rect 312770 22170 312838 22226
rect 312894 22170 312962 22226
rect 313018 22170 313086 22226
rect 313142 22170 313238 22226
rect 312618 22102 313238 22170
rect 312618 22046 312714 22102
rect 312770 22046 312838 22102
rect 312894 22046 312962 22102
rect 313018 22046 313086 22102
rect 313142 22046 313238 22102
rect 312618 21978 313238 22046
rect 312618 21922 312714 21978
rect 312770 21922 312838 21978
rect 312894 21922 312962 21978
rect 313018 21922 313086 21978
rect 313142 21922 313238 21978
rect 285618 -1176 285714 -1120
rect 285770 -1176 285838 -1120
rect 285894 -1176 285962 -1120
rect 286018 -1176 286086 -1120
rect 286142 -1176 286238 -1120
rect 285618 -1244 286238 -1176
rect 285618 -1300 285714 -1244
rect 285770 -1300 285838 -1244
rect 285894 -1300 285962 -1244
rect 286018 -1300 286086 -1244
rect 286142 -1300 286238 -1244
rect 285618 -1368 286238 -1300
rect 285618 -1424 285714 -1368
rect 285770 -1424 285838 -1368
rect 285894 -1424 285962 -1368
rect 286018 -1424 286086 -1368
rect 286142 -1424 286238 -1368
rect 285618 -1492 286238 -1424
rect 285618 -1548 285714 -1492
rect 285770 -1548 285838 -1492
rect 285894 -1548 285962 -1492
rect 286018 -1548 286086 -1492
rect 286142 -1548 286238 -1492
rect 285618 -1644 286238 -1548
rect 312618 4350 313238 21922
rect 312618 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 313238 4350
rect 312618 4226 313238 4294
rect 312618 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 313238 4226
rect 312618 4102 313238 4170
rect 312618 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 313238 4102
rect 312618 3978 313238 4046
rect 312618 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 313238 3978
rect 312618 -160 313238 3922
rect 312618 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 313238 -160
rect 312618 -284 313238 -216
rect 312618 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 313238 -284
rect 312618 -408 313238 -340
rect 312618 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 313238 -408
rect 312618 -532 313238 -464
rect 312618 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 313238 -532
rect 312618 -1644 313238 -588
rect 316338 46350 316958 50964
rect 320908 50260 320964 212604
rect 343338 202350 343958 219922
rect 343338 202294 343434 202350
rect 343490 202294 343558 202350
rect 343614 202294 343682 202350
rect 343738 202294 343806 202350
rect 343862 202294 343958 202350
rect 343338 202226 343958 202294
rect 343338 202170 343434 202226
rect 343490 202170 343558 202226
rect 343614 202170 343682 202226
rect 343738 202170 343806 202226
rect 343862 202170 343958 202226
rect 343338 202102 343958 202170
rect 343338 202046 343434 202102
rect 343490 202046 343558 202102
rect 343614 202046 343682 202102
rect 343738 202046 343806 202102
rect 343862 202046 343958 202102
rect 343338 201978 343958 202046
rect 343338 201922 343434 201978
rect 343490 201922 343558 201978
rect 343614 201922 343682 201978
rect 343738 201922 343806 201978
rect 343862 201922 343958 201978
rect 343338 184350 343958 201922
rect 343338 184294 343434 184350
rect 343490 184294 343558 184350
rect 343614 184294 343682 184350
rect 343738 184294 343806 184350
rect 343862 184294 343958 184350
rect 343338 184226 343958 184294
rect 343338 184170 343434 184226
rect 343490 184170 343558 184226
rect 343614 184170 343682 184226
rect 343738 184170 343806 184226
rect 343862 184170 343958 184226
rect 343338 184102 343958 184170
rect 343338 184046 343434 184102
rect 343490 184046 343558 184102
rect 343614 184046 343682 184102
rect 343738 184046 343806 184102
rect 343862 184046 343958 184102
rect 343338 183978 343958 184046
rect 343338 183922 343434 183978
rect 343490 183922 343558 183978
rect 343614 183922 343682 183978
rect 343738 183922 343806 183978
rect 343862 183922 343958 183978
rect 343338 166350 343958 183922
rect 343338 166294 343434 166350
rect 343490 166294 343558 166350
rect 343614 166294 343682 166350
rect 343738 166294 343806 166350
rect 343862 166294 343958 166350
rect 343338 166226 343958 166294
rect 343338 166170 343434 166226
rect 343490 166170 343558 166226
rect 343614 166170 343682 166226
rect 343738 166170 343806 166226
rect 343862 166170 343958 166226
rect 343338 166102 343958 166170
rect 343338 166046 343434 166102
rect 343490 166046 343558 166102
rect 343614 166046 343682 166102
rect 343738 166046 343806 166102
rect 343862 166046 343958 166102
rect 343338 165978 343958 166046
rect 343338 165922 343434 165978
rect 343490 165922 343558 165978
rect 343614 165922 343682 165978
rect 343738 165922 343806 165978
rect 343862 165922 343958 165978
rect 343338 148350 343958 165922
rect 343338 148294 343434 148350
rect 343490 148294 343558 148350
rect 343614 148294 343682 148350
rect 343738 148294 343806 148350
rect 343862 148294 343958 148350
rect 343338 148226 343958 148294
rect 343338 148170 343434 148226
rect 343490 148170 343558 148226
rect 343614 148170 343682 148226
rect 343738 148170 343806 148226
rect 343862 148170 343958 148226
rect 343338 148102 343958 148170
rect 343338 148046 343434 148102
rect 343490 148046 343558 148102
rect 343614 148046 343682 148102
rect 343738 148046 343806 148102
rect 343862 148046 343958 148102
rect 343338 147978 343958 148046
rect 343338 147922 343434 147978
rect 343490 147922 343558 147978
rect 343614 147922 343682 147978
rect 343738 147922 343806 147978
rect 343862 147922 343958 147978
rect 343338 130350 343958 147922
rect 343338 130294 343434 130350
rect 343490 130294 343558 130350
rect 343614 130294 343682 130350
rect 343738 130294 343806 130350
rect 343862 130294 343958 130350
rect 343338 130226 343958 130294
rect 343338 130170 343434 130226
rect 343490 130170 343558 130226
rect 343614 130170 343682 130226
rect 343738 130170 343806 130226
rect 343862 130170 343958 130226
rect 343338 130102 343958 130170
rect 343338 130046 343434 130102
rect 343490 130046 343558 130102
rect 343614 130046 343682 130102
rect 343738 130046 343806 130102
rect 343862 130046 343958 130102
rect 343338 129978 343958 130046
rect 343338 129922 343434 129978
rect 343490 129922 343558 129978
rect 343614 129922 343682 129978
rect 343738 129922 343806 129978
rect 343862 129922 343958 129978
rect 343338 112350 343958 129922
rect 343338 112294 343434 112350
rect 343490 112294 343558 112350
rect 343614 112294 343682 112350
rect 343738 112294 343806 112350
rect 343862 112294 343958 112350
rect 343338 112226 343958 112294
rect 343338 112170 343434 112226
rect 343490 112170 343558 112226
rect 343614 112170 343682 112226
rect 343738 112170 343806 112226
rect 343862 112170 343958 112226
rect 343338 112102 343958 112170
rect 343338 112046 343434 112102
rect 343490 112046 343558 112102
rect 343614 112046 343682 112102
rect 343738 112046 343806 112102
rect 343862 112046 343958 112102
rect 343338 111978 343958 112046
rect 343338 111922 343434 111978
rect 343490 111922 343558 111978
rect 343614 111922 343682 111978
rect 343738 111922 343806 111978
rect 343862 111922 343958 111978
rect 343338 94350 343958 111922
rect 343338 94294 343434 94350
rect 343490 94294 343558 94350
rect 343614 94294 343682 94350
rect 343738 94294 343806 94350
rect 343862 94294 343958 94350
rect 343338 94226 343958 94294
rect 343338 94170 343434 94226
rect 343490 94170 343558 94226
rect 343614 94170 343682 94226
rect 343738 94170 343806 94226
rect 343862 94170 343958 94226
rect 343338 94102 343958 94170
rect 343338 94046 343434 94102
rect 343490 94046 343558 94102
rect 343614 94046 343682 94102
rect 343738 94046 343806 94102
rect 343862 94046 343958 94102
rect 343338 93978 343958 94046
rect 343338 93922 343434 93978
rect 343490 93922 343558 93978
rect 343614 93922 343682 93978
rect 343738 93922 343806 93978
rect 343862 93922 343958 93978
rect 324448 82147 324768 82204
rect 324448 82091 324476 82147
rect 324532 82091 324580 82147
rect 324636 82091 324684 82147
rect 324740 82091 324768 82147
rect 324448 82043 324768 82091
rect 324448 81987 324476 82043
rect 324532 81987 324580 82043
rect 324636 81987 324684 82043
rect 324740 81987 324768 82043
rect 324448 81939 324768 81987
rect 324448 81883 324476 81939
rect 324532 81883 324580 81939
rect 324636 81883 324684 81939
rect 324740 81883 324768 81939
rect 324448 81826 324768 81883
rect 343338 76350 343958 93922
rect 343338 76294 343434 76350
rect 343490 76294 343558 76350
rect 343614 76294 343682 76350
rect 343738 76294 343806 76350
rect 343862 76294 343958 76350
rect 343338 76226 343958 76294
rect 343338 76170 343434 76226
rect 343490 76170 343558 76226
rect 343614 76170 343682 76226
rect 343738 76170 343806 76226
rect 343862 76170 343958 76226
rect 343338 76102 343958 76170
rect 343338 76046 343434 76102
rect 343490 76046 343558 76102
rect 343614 76046 343682 76102
rect 343738 76046 343806 76102
rect 343862 76046 343958 76102
rect 343338 75978 343958 76046
rect 343338 75922 343434 75978
rect 343490 75922 343558 75978
rect 343614 75922 343682 75978
rect 343738 75922 343806 75978
rect 343862 75922 343958 75978
rect 324448 64350 324768 64384
rect 324448 64294 324518 64350
rect 324574 64294 324642 64350
rect 324698 64294 324768 64350
rect 324448 64226 324768 64294
rect 324448 64170 324518 64226
rect 324574 64170 324642 64226
rect 324698 64170 324768 64226
rect 324448 64102 324768 64170
rect 324448 64046 324518 64102
rect 324574 64046 324642 64102
rect 324698 64046 324768 64102
rect 324448 63978 324768 64046
rect 324448 63922 324518 63978
rect 324574 63922 324642 63978
rect 324698 63922 324768 63978
rect 324448 63888 324768 63922
rect 320908 50194 320964 50204
rect 343338 58350 343958 75922
rect 343338 58294 343434 58350
rect 343490 58294 343558 58350
rect 343614 58294 343682 58350
rect 343738 58294 343806 58350
rect 343862 58294 343958 58350
rect 343338 58226 343958 58294
rect 343338 58170 343434 58226
rect 343490 58170 343558 58226
rect 343614 58170 343682 58226
rect 343738 58170 343806 58226
rect 343862 58170 343958 58226
rect 343338 58102 343958 58170
rect 343338 58046 343434 58102
rect 343490 58046 343558 58102
rect 343614 58046 343682 58102
rect 343738 58046 343806 58102
rect 343862 58046 343958 58102
rect 343338 57978 343958 58046
rect 343338 57922 343434 57978
rect 343490 57922 343558 57978
rect 343614 57922 343682 57978
rect 343738 57922 343806 57978
rect 343862 57922 343958 57978
rect 316338 46294 316434 46350
rect 316490 46294 316558 46350
rect 316614 46294 316682 46350
rect 316738 46294 316806 46350
rect 316862 46294 316958 46350
rect 316338 46226 316958 46294
rect 316338 46170 316434 46226
rect 316490 46170 316558 46226
rect 316614 46170 316682 46226
rect 316738 46170 316806 46226
rect 316862 46170 316958 46226
rect 316338 46102 316958 46170
rect 316338 46046 316434 46102
rect 316490 46046 316558 46102
rect 316614 46046 316682 46102
rect 316738 46046 316806 46102
rect 316862 46046 316958 46102
rect 316338 45978 316958 46046
rect 316338 45922 316434 45978
rect 316490 45922 316558 45978
rect 316614 45922 316682 45978
rect 316738 45922 316806 45978
rect 316862 45922 316958 45978
rect 316338 28350 316958 45922
rect 316338 28294 316434 28350
rect 316490 28294 316558 28350
rect 316614 28294 316682 28350
rect 316738 28294 316806 28350
rect 316862 28294 316958 28350
rect 316338 28226 316958 28294
rect 316338 28170 316434 28226
rect 316490 28170 316558 28226
rect 316614 28170 316682 28226
rect 316738 28170 316806 28226
rect 316862 28170 316958 28226
rect 316338 28102 316958 28170
rect 316338 28046 316434 28102
rect 316490 28046 316558 28102
rect 316614 28046 316682 28102
rect 316738 28046 316806 28102
rect 316862 28046 316958 28102
rect 316338 27978 316958 28046
rect 316338 27922 316434 27978
rect 316490 27922 316558 27978
rect 316614 27922 316682 27978
rect 316738 27922 316806 27978
rect 316862 27922 316958 27978
rect 316338 10350 316958 27922
rect 316338 10294 316434 10350
rect 316490 10294 316558 10350
rect 316614 10294 316682 10350
rect 316738 10294 316806 10350
rect 316862 10294 316958 10350
rect 316338 10226 316958 10294
rect 316338 10170 316434 10226
rect 316490 10170 316558 10226
rect 316614 10170 316682 10226
rect 316738 10170 316806 10226
rect 316862 10170 316958 10226
rect 316338 10102 316958 10170
rect 316338 10046 316434 10102
rect 316490 10046 316558 10102
rect 316614 10046 316682 10102
rect 316738 10046 316806 10102
rect 316862 10046 316958 10102
rect 316338 9978 316958 10046
rect 316338 9922 316434 9978
rect 316490 9922 316558 9978
rect 316614 9922 316682 9978
rect 316738 9922 316806 9978
rect 316862 9922 316958 9978
rect 316338 -1120 316958 9922
rect 316338 -1176 316434 -1120
rect 316490 -1176 316558 -1120
rect 316614 -1176 316682 -1120
rect 316738 -1176 316806 -1120
rect 316862 -1176 316958 -1120
rect 316338 -1244 316958 -1176
rect 316338 -1300 316434 -1244
rect 316490 -1300 316558 -1244
rect 316614 -1300 316682 -1244
rect 316738 -1300 316806 -1244
rect 316862 -1300 316958 -1244
rect 316338 -1368 316958 -1300
rect 316338 -1424 316434 -1368
rect 316490 -1424 316558 -1368
rect 316614 -1424 316682 -1368
rect 316738 -1424 316806 -1368
rect 316862 -1424 316958 -1368
rect 316338 -1492 316958 -1424
rect 316338 -1548 316434 -1492
rect 316490 -1548 316558 -1492
rect 316614 -1548 316682 -1492
rect 316738 -1548 316806 -1492
rect 316862 -1548 316958 -1492
rect 316338 -1644 316958 -1548
rect 343338 40350 343958 57922
rect 343338 40294 343434 40350
rect 343490 40294 343558 40350
rect 343614 40294 343682 40350
rect 343738 40294 343806 40350
rect 343862 40294 343958 40350
rect 343338 40226 343958 40294
rect 343338 40170 343434 40226
rect 343490 40170 343558 40226
rect 343614 40170 343682 40226
rect 343738 40170 343806 40226
rect 343862 40170 343958 40226
rect 343338 40102 343958 40170
rect 343338 40046 343434 40102
rect 343490 40046 343558 40102
rect 343614 40046 343682 40102
rect 343738 40046 343806 40102
rect 343862 40046 343958 40102
rect 343338 39978 343958 40046
rect 343338 39922 343434 39978
rect 343490 39922 343558 39978
rect 343614 39922 343682 39978
rect 343738 39922 343806 39978
rect 343862 39922 343958 39978
rect 343338 22350 343958 39922
rect 343338 22294 343434 22350
rect 343490 22294 343558 22350
rect 343614 22294 343682 22350
rect 343738 22294 343806 22350
rect 343862 22294 343958 22350
rect 343338 22226 343958 22294
rect 343338 22170 343434 22226
rect 343490 22170 343558 22226
rect 343614 22170 343682 22226
rect 343738 22170 343806 22226
rect 343862 22170 343958 22226
rect 343338 22102 343958 22170
rect 343338 22046 343434 22102
rect 343490 22046 343558 22102
rect 343614 22046 343682 22102
rect 343738 22046 343806 22102
rect 343862 22046 343958 22102
rect 343338 21978 343958 22046
rect 343338 21922 343434 21978
rect 343490 21922 343558 21978
rect 343614 21922 343682 21978
rect 343738 21922 343806 21978
rect 343862 21922 343958 21978
rect 343338 4350 343958 21922
rect 343338 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 343958 4350
rect 343338 4226 343958 4294
rect 343338 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 343958 4226
rect 343338 4102 343958 4170
rect 343338 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 343958 4102
rect 343338 3978 343958 4046
rect 343338 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 343958 3978
rect 343338 -160 343958 3922
rect 343338 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 343958 -160
rect 343338 -284 343958 -216
rect 343338 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 343958 -284
rect 343338 -408 343958 -340
rect 343338 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 343958 -408
rect 343338 -532 343958 -464
rect 343338 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 343958 -532
rect 343338 -1644 343958 -588
rect 347058 244350 347678 257490
rect 347058 244294 347154 244350
rect 347210 244294 347278 244350
rect 347334 244294 347402 244350
rect 347458 244294 347526 244350
rect 347582 244294 347678 244350
rect 347058 244226 347678 244294
rect 347058 244170 347154 244226
rect 347210 244170 347278 244226
rect 347334 244170 347402 244226
rect 347458 244170 347526 244226
rect 347582 244170 347678 244226
rect 347058 244102 347678 244170
rect 347058 244046 347154 244102
rect 347210 244046 347278 244102
rect 347334 244046 347402 244102
rect 347458 244046 347526 244102
rect 347582 244046 347678 244102
rect 347058 243978 347678 244046
rect 347058 243922 347154 243978
rect 347210 243922 347278 243978
rect 347334 243922 347402 243978
rect 347458 243922 347526 243978
rect 347582 243922 347678 243978
rect 347058 226350 347678 243922
rect 347058 226294 347154 226350
rect 347210 226294 347278 226350
rect 347334 226294 347402 226350
rect 347458 226294 347526 226350
rect 347582 226294 347678 226350
rect 347058 226226 347678 226294
rect 347058 226170 347154 226226
rect 347210 226170 347278 226226
rect 347334 226170 347402 226226
rect 347458 226170 347526 226226
rect 347582 226170 347678 226226
rect 347058 226102 347678 226170
rect 347058 226046 347154 226102
rect 347210 226046 347278 226102
rect 347334 226046 347402 226102
rect 347458 226046 347526 226102
rect 347582 226046 347678 226102
rect 347058 225978 347678 226046
rect 347058 225922 347154 225978
rect 347210 225922 347278 225978
rect 347334 225922 347402 225978
rect 347458 225922 347526 225978
rect 347582 225922 347678 225978
rect 347058 208350 347678 225922
rect 347058 208294 347154 208350
rect 347210 208294 347278 208350
rect 347334 208294 347402 208350
rect 347458 208294 347526 208350
rect 347582 208294 347678 208350
rect 347058 208226 347678 208294
rect 347058 208170 347154 208226
rect 347210 208170 347278 208226
rect 347334 208170 347402 208226
rect 347458 208170 347526 208226
rect 347582 208170 347678 208226
rect 347058 208102 347678 208170
rect 347058 208046 347154 208102
rect 347210 208046 347278 208102
rect 347334 208046 347402 208102
rect 347458 208046 347526 208102
rect 347582 208046 347678 208102
rect 347058 207978 347678 208046
rect 347058 207922 347154 207978
rect 347210 207922 347278 207978
rect 347334 207922 347402 207978
rect 347458 207922 347526 207978
rect 347582 207922 347678 207978
rect 347058 190350 347678 207922
rect 347058 190294 347154 190350
rect 347210 190294 347278 190350
rect 347334 190294 347402 190350
rect 347458 190294 347526 190350
rect 347582 190294 347678 190350
rect 347058 190226 347678 190294
rect 347058 190170 347154 190226
rect 347210 190170 347278 190226
rect 347334 190170 347402 190226
rect 347458 190170 347526 190226
rect 347582 190170 347678 190226
rect 347058 190102 347678 190170
rect 347058 190046 347154 190102
rect 347210 190046 347278 190102
rect 347334 190046 347402 190102
rect 347458 190046 347526 190102
rect 347582 190046 347678 190102
rect 347058 189978 347678 190046
rect 347058 189922 347154 189978
rect 347210 189922 347278 189978
rect 347334 189922 347402 189978
rect 347458 189922 347526 189978
rect 347582 189922 347678 189978
rect 347058 172350 347678 189922
rect 347058 172294 347154 172350
rect 347210 172294 347278 172350
rect 347334 172294 347402 172350
rect 347458 172294 347526 172350
rect 347582 172294 347678 172350
rect 347058 172226 347678 172294
rect 347058 172170 347154 172226
rect 347210 172170 347278 172226
rect 347334 172170 347402 172226
rect 347458 172170 347526 172226
rect 347582 172170 347678 172226
rect 347058 172102 347678 172170
rect 347058 172046 347154 172102
rect 347210 172046 347278 172102
rect 347334 172046 347402 172102
rect 347458 172046 347526 172102
rect 347582 172046 347678 172102
rect 347058 171978 347678 172046
rect 347058 171922 347154 171978
rect 347210 171922 347278 171978
rect 347334 171922 347402 171978
rect 347458 171922 347526 171978
rect 347582 171922 347678 171978
rect 347058 154350 347678 171922
rect 347058 154294 347154 154350
rect 347210 154294 347278 154350
rect 347334 154294 347402 154350
rect 347458 154294 347526 154350
rect 347582 154294 347678 154350
rect 347058 154226 347678 154294
rect 347058 154170 347154 154226
rect 347210 154170 347278 154226
rect 347334 154170 347402 154226
rect 347458 154170 347526 154226
rect 347582 154170 347678 154226
rect 347058 154102 347678 154170
rect 347058 154046 347154 154102
rect 347210 154046 347278 154102
rect 347334 154046 347402 154102
rect 347458 154046 347526 154102
rect 347582 154046 347678 154102
rect 347058 153978 347678 154046
rect 347058 153922 347154 153978
rect 347210 153922 347278 153978
rect 347334 153922 347402 153978
rect 347458 153922 347526 153978
rect 347582 153922 347678 153978
rect 347058 136350 347678 153922
rect 347058 136294 347154 136350
rect 347210 136294 347278 136350
rect 347334 136294 347402 136350
rect 347458 136294 347526 136350
rect 347582 136294 347678 136350
rect 347058 136226 347678 136294
rect 347058 136170 347154 136226
rect 347210 136170 347278 136226
rect 347334 136170 347402 136226
rect 347458 136170 347526 136226
rect 347582 136170 347678 136226
rect 347058 136102 347678 136170
rect 347058 136046 347154 136102
rect 347210 136046 347278 136102
rect 347334 136046 347402 136102
rect 347458 136046 347526 136102
rect 347582 136046 347678 136102
rect 347058 135978 347678 136046
rect 347058 135922 347154 135978
rect 347210 135922 347278 135978
rect 347334 135922 347402 135978
rect 347458 135922 347526 135978
rect 347582 135922 347678 135978
rect 347058 118350 347678 135922
rect 347058 118294 347154 118350
rect 347210 118294 347278 118350
rect 347334 118294 347402 118350
rect 347458 118294 347526 118350
rect 347582 118294 347678 118350
rect 347058 118226 347678 118294
rect 347058 118170 347154 118226
rect 347210 118170 347278 118226
rect 347334 118170 347402 118226
rect 347458 118170 347526 118226
rect 347582 118170 347678 118226
rect 347058 118102 347678 118170
rect 347058 118046 347154 118102
rect 347210 118046 347278 118102
rect 347334 118046 347402 118102
rect 347458 118046 347526 118102
rect 347582 118046 347678 118102
rect 347058 117978 347678 118046
rect 347058 117922 347154 117978
rect 347210 117922 347278 117978
rect 347334 117922 347402 117978
rect 347458 117922 347526 117978
rect 347582 117922 347678 117978
rect 347058 100350 347678 117922
rect 347058 100294 347154 100350
rect 347210 100294 347278 100350
rect 347334 100294 347402 100350
rect 347458 100294 347526 100350
rect 347582 100294 347678 100350
rect 347058 100226 347678 100294
rect 347058 100170 347154 100226
rect 347210 100170 347278 100226
rect 347334 100170 347402 100226
rect 347458 100170 347526 100226
rect 347582 100170 347678 100226
rect 347058 100102 347678 100170
rect 347058 100046 347154 100102
rect 347210 100046 347278 100102
rect 347334 100046 347402 100102
rect 347458 100046 347526 100102
rect 347582 100046 347678 100102
rect 347058 99978 347678 100046
rect 347058 99922 347154 99978
rect 347210 99922 347278 99978
rect 347334 99922 347402 99978
rect 347458 99922 347526 99978
rect 347582 99922 347678 99978
rect 347058 82350 347678 99922
rect 347058 82294 347154 82350
rect 347210 82294 347278 82350
rect 347334 82294 347402 82350
rect 347458 82294 347526 82350
rect 347582 82294 347678 82350
rect 347058 82226 347678 82294
rect 347058 82170 347154 82226
rect 347210 82170 347278 82226
rect 347334 82170 347402 82226
rect 347458 82170 347526 82226
rect 347582 82170 347678 82226
rect 347058 82102 347678 82170
rect 347058 82046 347154 82102
rect 347210 82046 347278 82102
rect 347334 82046 347402 82102
rect 347458 82046 347526 82102
rect 347582 82046 347678 82102
rect 347058 81978 347678 82046
rect 347058 81922 347154 81978
rect 347210 81922 347278 81978
rect 347334 81922 347402 81978
rect 347458 81922 347526 81978
rect 347582 81922 347678 81978
rect 347058 64350 347678 81922
rect 347058 64294 347154 64350
rect 347210 64294 347278 64350
rect 347334 64294 347402 64350
rect 347458 64294 347526 64350
rect 347582 64294 347678 64350
rect 347058 64226 347678 64294
rect 347058 64170 347154 64226
rect 347210 64170 347278 64226
rect 347334 64170 347402 64226
rect 347458 64170 347526 64226
rect 347582 64170 347678 64226
rect 347058 64102 347678 64170
rect 347058 64046 347154 64102
rect 347210 64046 347278 64102
rect 347334 64046 347402 64102
rect 347458 64046 347526 64102
rect 347582 64046 347678 64102
rect 347058 63978 347678 64046
rect 347058 63922 347154 63978
rect 347210 63922 347278 63978
rect 347334 63922 347402 63978
rect 347458 63922 347526 63978
rect 347582 63922 347678 63978
rect 347058 46350 347678 63922
rect 347058 46294 347154 46350
rect 347210 46294 347278 46350
rect 347334 46294 347402 46350
rect 347458 46294 347526 46350
rect 347582 46294 347678 46350
rect 347058 46226 347678 46294
rect 347058 46170 347154 46226
rect 347210 46170 347278 46226
rect 347334 46170 347402 46226
rect 347458 46170 347526 46226
rect 347582 46170 347678 46226
rect 347058 46102 347678 46170
rect 347058 46046 347154 46102
rect 347210 46046 347278 46102
rect 347334 46046 347402 46102
rect 347458 46046 347526 46102
rect 347582 46046 347678 46102
rect 347058 45978 347678 46046
rect 347058 45922 347154 45978
rect 347210 45922 347278 45978
rect 347334 45922 347402 45978
rect 347458 45922 347526 45978
rect 347582 45922 347678 45978
rect 347058 28350 347678 45922
rect 347058 28294 347154 28350
rect 347210 28294 347278 28350
rect 347334 28294 347402 28350
rect 347458 28294 347526 28350
rect 347582 28294 347678 28350
rect 347058 28226 347678 28294
rect 347058 28170 347154 28226
rect 347210 28170 347278 28226
rect 347334 28170 347402 28226
rect 347458 28170 347526 28226
rect 347582 28170 347678 28226
rect 347058 28102 347678 28170
rect 347058 28046 347154 28102
rect 347210 28046 347278 28102
rect 347334 28046 347402 28102
rect 347458 28046 347526 28102
rect 347582 28046 347678 28102
rect 347058 27978 347678 28046
rect 347058 27922 347154 27978
rect 347210 27922 347278 27978
rect 347334 27922 347402 27978
rect 347458 27922 347526 27978
rect 347582 27922 347678 27978
rect 347058 10350 347678 27922
rect 347058 10294 347154 10350
rect 347210 10294 347278 10350
rect 347334 10294 347402 10350
rect 347458 10294 347526 10350
rect 347582 10294 347678 10350
rect 347058 10226 347678 10294
rect 347058 10170 347154 10226
rect 347210 10170 347278 10226
rect 347334 10170 347402 10226
rect 347458 10170 347526 10226
rect 347582 10170 347678 10226
rect 347058 10102 347678 10170
rect 347058 10046 347154 10102
rect 347210 10046 347278 10102
rect 347334 10046 347402 10102
rect 347458 10046 347526 10102
rect 347582 10046 347678 10102
rect 347058 9978 347678 10046
rect 347058 9922 347154 9978
rect 347210 9922 347278 9978
rect 347334 9922 347402 9978
rect 347458 9922 347526 9978
rect 347582 9922 347678 9978
rect 347058 -1120 347678 9922
rect 348572 257348 348628 257358
rect 348572 4788 348628 257292
rect 358652 41188 358708 257822
rect 362012 256004 362068 256014
rect 358652 41122 358708 41132
rect 358764 253198 358820 253208
rect 358764 38164 358820 253142
rect 358988 253018 359044 253028
rect 358988 41412 359044 252962
rect 359212 252838 359268 252848
rect 359212 44660 359268 252782
rect 359212 44594 359268 44604
rect 358988 41346 359044 41356
rect 362012 41300 362068 255948
rect 362124 255892 362180 255902
rect 362124 49588 362180 255836
rect 367052 154420 367108 154430
rect 367052 153972 367108 154364
rect 367052 153906 367108 153916
rect 371308 154196 371364 154206
rect 371308 153748 371364 154140
rect 372316 154196 372372 386092
rect 372316 154130 372372 154140
rect 372428 386036 372484 386046
rect 371308 153682 371364 153692
rect 372428 153658 372484 385980
rect 372988 154084 373044 393148
rect 375452 388108 375508 407596
rect 375228 388052 375508 388108
rect 375676 402836 375732 402846
rect 373100 385678 373156 385688
rect 373100 160692 373156 385622
rect 375228 376348 375284 388052
rect 375564 385924 375620 385934
rect 375228 376292 375508 376348
rect 375228 288372 375284 288382
rect 373772 288298 373828 288308
rect 373772 253316 373828 288242
rect 375228 288298 375284 288316
rect 375228 288232 375284 288242
rect 373772 253250 373828 253260
rect 373884 286138 373940 286148
rect 373884 253198 373940 286082
rect 375228 286138 375284 286170
rect 375228 286066 375284 286076
rect 375228 265972 375284 265982
rect 375228 257878 375284 265916
rect 375228 257812 375284 257822
rect 373884 253132 373940 253142
rect 374058 256350 374678 257490
rect 374058 256294 374154 256350
rect 374210 256294 374278 256350
rect 374334 256294 374402 256350
rect 374458 256294 374526 256350
rect 374582 256294 374678 256350
rect 374058 256226 374678 256294
rect 374058 256170 374154 256226
rect 374210 256170 374278 256226
rect 374334 256170 374402 256226
rect 374458 256170 374526 256226
rect 374582 256170 374678 256226
rect 374058 256102 374678 256170
rect 374058 256046 374154 256102
rect 374210 256046 374278 256102
rect 374334 256046 374402 256102
rect 374458 256046 374526 256102
rect 374582 256046 374678 256102
rect 374058 255978 374678 256046
rect 374058 255922 374154 255978
rect 374210 255922 374278 255978
rect 374334 255922 374402 255978
rect 374458 255922 374526 255978
rect 374582 255922 374678 255978
rect 373100 160626 373156 160636
rect 374058 238350 374678 255922
rect 374058 238294 374154 238350
rect 374210 238294 374278 238350
rect 374334 238294 374402 238350
rect 374458 238294 374526 238350
rect 374582 238294 374678 238350
rect 374058 238226 374678 238294
rect 374058 238170 374154 238226
rect 374210 238170 374278 238226
rect 374334 238170 374402 238226
rect 374458 238170 374526 238226
rect 374582 238170 374678 238226
rect 374058 238102 374678 238170
rect 374058 238046 374154 238102
rect 374210 238046 374278 238102
rect 374334 238046 374402 238102
rect 374458 238046 374526 238102
rect 374582 238046 374678 238102
rect 374058 237978 374678 238046
rect 374058 237922 374154 237978
rect 374210 237922 374278 237978
rect 374334 237922 374402 237978
rect 374458 237922 374526 237978
rect 374582 237922 374678 237978
rect 374058 220350 374678 237922
rect 374058 220294 374154 220350
rect 374210 220294 374278 220350
rect 374334 220294 374402 220350
rect 374458 220294 374526 220350
rect 374582 220294 374678 220350
rect 374058 220226 374678 220294
rect 374058 220170 374154 220226
rect 374210 220170 374278 220226
rect 374334 220170 374402 220226
rect 374458 220170 374526 220226
rect 374582 220170 374678 220226
rect 374058 220102 374678 220170
rect 374058 220046 374154 220102
rect 374210 220046 374278 220102
rect 374334 220046 374402 220102
rect 374458 220046 374526 220102
rect 374582 220046 374678 220102
rect 374058 219978 374678 220046
rect 374058 219922 374154 219978
rect 374210 219922 374278 219978
rect 374334 219922 374402 219978
rect 374458 219922 374526 219978
rect 374582 219922 374678 219978
rect 374058 202350 374678 219922
rect 374058 202294 374154 202350
rect 374210 202294 374278 202350
rect 374334 202294 374402 202350
rect 374458 202294 374526 202350
rect 374582 202294 374678 202350
rect 374058 202226 374678 202294
rect 374058 202170 374154 202226
rect 374210 202170 374278 202226
rect 374334 202170 374402 202226
rect 374458 202170 374526 202226
rect 374582 202170 374678 202226
rect 374058 202102 374678 202170
rect 374058 202046 374154 202102
rect 374210 202046 374278 202102
rect 374334 202046 374402 202102
rect 374458 202046 374526 202102
rect 374582 202046 374678 202102
rect 374058 201978 374678 202046
rect 374058 201922 374154 201978
rect 374210 201922 374278 201978
rect 374334 201922 374402 201978
rect 374458 201922 374526 201978
rect 374582 201922 374678 201978
rect 374058 184350 374678 201922
rect 374058 184294 374154 184350
rect 374210 184294 374278 184350
rect 374334 184294 374402 184350
rect 374458 184294 374526 184350
rect 374582 184294 374678 184350
rect 374058 184226 374678 184294
rect 374058 184170 374154 184226
rect 374210 184170 374278 184226
rect 374334 184170 374402 184226
rect 374458 184170 374526 184226
rect 374582 184170 374678 184226
rect 374058 184102 374678 184170
rect 374058 184046 374154 184102
rect 374210 184046 374278 184102
rect 374334 184046 374402 184102
rect 374458 184046 374526 184102
rect 374582 184046 374678 184102
rect 374058 183978 374678 184046
rect 374058 183922 374154 183978
rect 374210 183922 374278 183978
rect 374334 183922 374402 183978
rect 374458 183922 374526 183978
rect 374582 183922 374678 183978
rect 374058 166350 374678 183922
rect 374058 166294 374154 166350
rect 374210 166294 374278 166350
rect 374334 166294 374402 166350
rect 374458 166294 374526 166350
rect 374582 166294 374678 166350
rect 374058 166226 374678 166294
rect 374058 166170 374154 166226
rect 374210 166170 374278 166226
rect 374334 166170 374402 166226
rect 374458 166170 374526 166226
rect 374582 166170 374678 166226
rect 374058 166102 374678 166170
rect 374058 166046 374154 166102
rect 374210 166046 374278 166102
rect 374334 166046 374402 166102
rect 374458 166046 374526 166102
rect 374582 166046 374678 166102
rect 374058 165978 374678 166046
rect 374058 165922 374154 165978
rect 374210 165922 374278 165978
rect 374334 165922 374402 165978
rect 374458 165922 374526 165978
rect 374582 165922 374678 165978
rect 372988 154018 373044 154028
rect 372428 153592 372484 153602
rect 374058 148350 374678 165922
rect 375452 153972 375508 376292
rect 375564 160804 375620 385868
rect 375676 319732 375732 402780
rect 375676 319666 375732 319676
rect 376348 314132 376404 408940
rect 377778 406350 378398 408578
rect 377778 406294 377874 406350
rect 377930 406294 377998 406350
rect 378054 406294 378122 406350
rect 378178 406294 378246 406350
rect 378302 406294 378398 406350
rect 377778 406226 378398 406294
rect 377778 406170 377874 406226
rect 377930 406170 377998 406226
rect 378054 406170 378122 406226
rect 378178 406170 378246 406226
rect 378302 406170 378398 406226
rect 377778 406102 378398 406170
rect 377778 406046 377874 406102
rect 377930 406046 377998 406102
rect 378054 406046 378122 406102
rect 378178 406046 378246 406102
rect 378302 406046 378398 406102
rect 377778 405978 378398 406046
rect 377778 405922 377874 405978
rect 377930 405922 377998 405978
rect 378054 405922 378122 405978
rect 378178 405922 378246 405978
rect 378302 405922 378398 405978
rect 376460 404292 376516 404302
rect 376460 317492 376516 404236
rect 376460 317426 376516 317436
rect 376572 396340 376628 396350
rect 376572 315252 376628 396284
rect 376572 315186 376628 315196
rect 377778 388350 378398 405922
rect 377778 388294 377874 388350
rect 377930 388294 377998 388350
rect 378054 388294 378122 388350
rect 378178 388294 378246 388350
rect 378302 388294 378398 388350
rect 377778 388226 378398 388294
rect 377778 388170 377874 388226
rect 377930 388170 377998 388226
rect 378054 388170 378122 388226
rect 378178 388170 378246 388226
rect 378302 388170 378398 388226
rect 377778 388102 378398 388170
rect 377778 388046 377874 388102
rect 377930 388046 377998 388102
rect 378054 388046 378122 388102
rect 378178 388046 378246 388102
rect 378302 388046 378398 388102
rect 377778 387978 378398 388046
rect 377778 387922 377874 387978
rect 377930 387922 377998 387978
rect 378054 387922 378122 387978
rect 378178 387922 378246 387978
rect 378302 387922 378398 387978
rect 377778 370350 378398 387922
rect 377778 370294 377874 370350
rect 377930 370294 377998 370350
rect 378054 370294 378122 370350
rect 378178 370294 378246 370350
rect 378302 370294 378398 370350
rect 377778 370226 378398 370294
rect 377778 370170 377874 370226
rect 377930 370170 377998 370226
rect 378054 370170 378122 370226
rect 378178 370170 378246 370226
rect 378302 370170 378398 370226
rect 377778 370102 378398 370170
rect 377778 370046 377874 370102
rect 377930 370046 377998 370102
rect 378054 370046 378122 370102
rect 378178 370046 378246 370102
rect 378302 370046 378398 370102
rect 377778 369978 378398 370046
rect 377778 369922 377874 369978
rect 377930 369922 377998 369978
rect 378054 369922 378122 369978
rect 378178 369922 378246 369978
rect 378302 369922 378398 369978
rect 377778 352350 378398 369922
rect 377778 352294 377874 352350
rect 377930 352294 377998 352350
rect 378054 352294 378122 352350
rect 378178 352294 378246 352350
rect 378302 352294 378398 352350
rect 377778 352226 378398 352294
rect 377778 352170 377874 352226
rect 377930 352170 377998 352226
rect 378054 352170 378122 352226
rect 378178 352170 378246 352226
rect 378302 352170 378398 352226
rect 377778 352102 378398 352170
rect 377778 352046 377874 352102
rect 377930 352046 377998 352102
rect 378054 352046 378122 352102
rect 378178 352046 378246 352102
rect 378302 352046 378398 352102
rect 377778 351978 378398 352046
rect 377778 351922 377874 351978
rect 377930 351922 377998 351978
rect 378054 351922 378122 351978
rect 378178 351922 378246 351978
rect 378302 351922 378398 351978
rect 377778 334350 378398 351922
rect 377778 334294 377874 334350
rect 377930 334294 377998 334350
rect 378054 334294 378122 334350
rect 378178 334294 378246 334350
rect 378302 334294 378398 334350
rect 377778 334226 378398 334294
rect 377778 334170 377874 334226
rect 377930 334170 377998 334226
rect 378054 334170 378122 334226
rect 378178 334170 378246 334226
rect 378302 334170 378398 334226
rect 377778 334102 378398 334170
rect 377778 334046 377874 334102
rect 377930 334046 377998 334102
rect 378054 334046 378122 334102
rect 378178 334046 378246 334102
rect 378302 334046 378398 334102
rect 377778 333978 378398 334046
rect 377778 333922 377874 333978
rect 377930 333922 377998 333978
rect 378054 333922 378122 333978
rect 378178 333922 378246 333978
rect 378302 333922 378398 333978
rect 377778 316350 378398 333922
rect 378476 405972 378532 405982
rect 378476 316708 378532 405916
rect 404778 400350 405398 408578
rect 404778 400294 404874 400350
rect 404930 400294 404998 400350
rect 405054 400294 405122 400350
rect 405178 400294 405246 400350
rect 405302 400294 405398 400350
rect 404778 400226 405398 400294
rect 404778 400170 404874 400226
rect 404930 400170 404998 400226
rect 405054 400170 405122 400226
rect 405178 400170 405246 400226
rect 405302 400170 405398 400226
rect 404778 400102 405398 400170
rect 404778 400046 404874 400102
rect 404930 400046 404998 400102
rect 405054 400046 405122 400102
rect 405178 400046 405246 400102
rect 405302 400046 405398 400102
rect 404778 399978 405398 400046
rect 404778 399922 404874 399978
rect 404930 399922 404998 399978
rect 405054 399922 405122 399978
rect 405178 399922 405246 399978
rect 405302 399922 405398 399978
rect 378700 399364 378756 399374
rect 378476 316642 378532 316652
rect 378588 396228 378644 396238
rect 377778 316294 377874 316350
rect 377930 316294 377998 316350
rect 378054 316294 378122 316350
rect 378178 316294 378246 316350
rect 378302 316294 378398 316350
rect 377778 316226 378398 316294
rect 377778 316170 377874 316226
rect 377930 316170 377998 316226
rect 378054 316170 378122 316226
rect 378178 316170 378246 316226
rect 378302 316170 378398 316226
rect 377778 316102 378398 316170
rect 377778 316046 377874 316102
rect 377930 316046 377998 316102
rect 378054 316046 378122 316102
rect 378178 316046 378246 316102
rect 378302 316046 378398 316102
rect 377778 315978 378398 316046
rect 377778 315922 377874 315978
rect 377930 315922 377998 315978
rect 378054 315922 378122 315978
rect 378178 315922 378246 315978
rect 378302 315922 378398 315978
rect 376348 314066 376404 314076
rect 376348 298452 376404 298462
rect 375676 283892 375732 283902
rect 375676 253018 375732 283836
rect 375788 271572 375844 271582
rect 375788 256004 375844 271516
rect 375788 255938 375844 255948
rect 375900 270452 375956 270462
rect 375900 255892 375956 270396
rect 375900 255826 375956 255836
rect 376124 261492 376180 261502
rect 375676 252952 375732 252962
rect 376124 232708 376180 261436
rect 376124 232642 376180 232652
rect 376236 259252 376292 259262
rect 376236 212548 376292 259196
rect 376348 229348 376404 298396
rect 377778 298350 378398 315922
rect 378588 313460 378644 396172
rect 378700 318388 378756 399308
rect 378812 397908 378868 397918
rect 378812 320068 378868 397852
rect 378924 396452 378980 396462
rect 378924 382452 378980 396396
rect 378924 382386 378980 382396
rect 383964 388738 384020 388748
rect 378924 370132 378980 370142
rect 378924 368788 378980 370076
rect 378924 368722 378980 368732
rect 379596 364532 379652 364542
rect 379596 362068 379652 364476
rect 379596 362002 379652 362012
rect 379596 361172 379652 361182
rect 379596 358708 379652 361116
rect 379596 358642 379652 358652
rect 379596 352212 379652 352222
rect 379596 350308 379652 352156
rect 379596 350242 379652 350252
rect 378812 320002 378868 320012
rect 380492 330932 380548 330942
rect 378700 318322 378756 318332
rect 378812 317492 378868 317502
rect 378812 315140 378868 317436
rect 378812 315074 378868 315084
rect 378588 313012 378644 313404
rect 378588 312946 378644 312956
rect 379484 306292 379540 306302
rect 379372 305172 379428 305182
rect 379260 304052 379316 304062
rect 379036 302932 379092 302942
rect 378924 301812 378980 301822
rect 377778 298294 377874 298350
rect 377930 298294 377998 298350
rect 378054 298294 378122 298350
rect 378178 298294 378246 298350
rect 378302 298294 378398 298350
rect 377778 298226 378398 298294
rect 377778 298170 377874 298226
rect 377930 298170 377998 298226
rect 378054 298170 378122 298226
rect 378178 298170 378246 298226
rect 378302 298170 378398 298226
rect 377778 298102 378398 298170
rect 377778 298046 377874 298102
rect 377930 298046 377998 298102
rect 378054 298046 378122 298102
rect 378178 298046 378246 298102
rect 378302 298046 378398 298102
rect 377778 297978 378398 298046
rect 377778 297922 377874 297978
rect 377930 297922 377998 297978
rect 378054 297922 378122 297978
rect 378178 297922 378246 297978
rect 378302 297922 378398 297978
rect 376460 281652 376516 281662
rect 376460 252838 376516 281596
rect 376460 252772 376516 252782
rect 377778 280350 378398 297922
rect 377778 280294 377874 280350
rect 377930 280294 377998 280350
rect 378054 280294 378122 280350
rect 378178 280294 378246 280350
rect 378302 280294 378398 280350
rect 377778 280226 378398 280294
rect 377778 280170 377874 280226
rect 377930 280170 377998 280226
rect 378054 280170 378122 280226
rect 378178 280170 378246 280226
rect 378302 280170 378398 280226
rect 377778 280102 378398 280170
rect 377778 280046 377874 280102
rect 377930 280046 377998 280102
rect 378054 280046 378122 280102
rect 378178 280046 378246 280102
rect 378302 280046 378398 280102
rect 377778 279978 378398 280046
rect 377778 279922 377874 279978
rect 377930 279922 377998 279978
rect 378054 279922 378122 279978
rect 378178 279922 378246 279978
rect 378302 279922 378398 279978
rect 377778 262350 378398 279922
rect 378812 299572 378868 299582
rect 378588 267092 378644 267102
rect 377778 262294 377874 262350
rect 377930 262294 377998 262350
rect 378054 262294 378122 262350
rect 378178 262294 378246 262350
rect 378302 262294 378398 262350
rect 377778 262226 378398 262294
rect 377778 262170 377874 262226
rect 377930 262170 377998 262226
rect 378054 262170 378122 262226
rect 378178 262170 378246 262226
rect 378302 262170 378398 262226
rect 377778 262102 378398 262170
rect 377778 262046 377874 262102
rect 377930 262046 377998 262102
rect 378054 262046 378122 262102
rect 378178 262046 378246 262102
rect 378302 262046 378398 262102
rect 377778 261978 378398 262046
rect 377778 261922 377874 261978
rect 377930 261922 377998 261978
rect 378054 261922 378122 261978
rect 378178 261922 378246 261978
rect 378302 261922 378398 261978
rect 376348 229282 376404 229292
rect 377778 244350 378398 261922
rect 377778 244294 377874 244350
rect 377930 244294 377998 244350
rect 378054 244294 378122 244350
rect 378178 244294 378246 244350
rect 378302 244294 378398 244350
rect 377778 244226 378398 244294
rect 377778 244170 377874 244226
rect 377930 244170 377998 244226
rect 378054 244170 378122 244226
rect 378178 244170 378246 244226
rect 378302 244170 378398 244226
rect 377778 244102 378398 244170
rect 377778 244046 377874 244102
rect 377930 244046 377998 244102
rect 378054 244046 378122 244102
rect 378178 244046 378246 244102
rect 378302 244046 378398 244102
rect 377778 243978 378398 244046
rect 377778 243922 377874 243978
rect 377930 243922 377998 243978
rect 378054 243922 378122 243978
rect 378178 243922 378246 243978
rect 378302 243922 378398 243978
rect 376236 212482 376292 212492
rect 377778 226350 378398 243922
rect 378476 262612 378532 262622
rect 378476 231028 378532 262556
rect 378588 248388 378644 267036
rect 378700 264852 378756 264862
rect 378700 248612 378756 264796
rect 378812 260484 378868 299516
rect 378924 265524 378980 301756
rect 379036 268772 379092 302876
rect 379036 268706 379092 268716
rect 379148 300692 379204 300702
rect 378924 265458 378980 265468
rect 379148 263844 379204 300636
rect 379260 270452 379316 303996
rect 379372 271918 379428 305116
rect 379484 273924 379540 306236
rect 379484 273858 379540 273868
rect 380268 273924 380324 273934
rect 379372 271862 379876 271918
rect 379260 270386 379316 270396
rect 379820 270564 379876 271862
rect 379148 263778 379204 263788
rect 379708 265524 379764 265534
rect 378812 255108 378868 260428
rect 378812 255042 378868 255052
rect 378924 263732 378980 263742
rect 378700 248546 378756 248556
rect 378588 248322 378644 248332
rect 378924 247716 378980 263676
rect 379708 256340 379764 265468
rect 379708 256274 379764 256284
rect 379820 250292 379876 270508
rect 380044 270452 380100 270462
rect 380044 268884 380100 270396
rect 379932 268772 379988 268782
rect 379932 267204 379988 268716
rect 379932 255780 379988 267148
rect 380044 257460 380100 268828
rect 380044 257394 380100 257404
rect 380156 263844 380212 263854
rect 379932 255714 379988 255724
rect 380156 254772 380212 263788
rect 380156 254706 380212 254716
rect 380268 251972 380324 273868
rect 380268 251906 380324 251916
rect 379820 250226 379876 250236
rect 378924 247650 378980 247660
rect 378476 230962 378532 230972
rect 377778 226294 377874 226350
rect 377930 226294 377998 226350
rect 378054 226294 378122 226350
rect 378178 226294 378246 226350
rect 378302 226294 378398 226350
rect 377778 226226 378398 226294
rect 377778 226170 377874 226226
rect 377930 226170 377998 226226
rect 378054 226170 378122 226226
rect 378178 226170 378246 226226
rect 378302 226170 378398 226226
rect 377778 226102 378398 226170
rect 377778 226046 377874 226102
rect 377930 226046 377998 226102
rect 378054 226046 378122 226102
rect 378178 226046 378246 226102
rect 378302 226046 378398 226102
rect 377778 225978 378398 226046
rect 377778 225922 377874 225978
rect 377930 225922 377998 225978
rect 378054 225922 378122 225978
rect 378178 225922 378246 225978
rect 378302 225922 378398 225978
rect 375564 160738 375620 160748
rect 377778 208350 378398 225922
rect 377778 208294 377874 208350
rect 377930 208294 377998 208350
rect 378054 208294 378122 208350
rect 378178 208294 378246 208350
rect 378302 208294 378398 208350
rect 377778 208226 378398 208294
rect 377778 208170 377874 208226
rect 377930 208170 377998 208226
rect 378054 208170 378122 208226
rect 378178 208170 378246 208226
rect 378302 208170 378398 208226
rect 377778 208102 378398 208170
rect 377778 208046 377874 208102
rect 377930 208046 377998 208102
rect 378054 208046 378122 208102
rect 378178 208046 378246 208102
rect 378302 208046 378398 208102
rect 377778 207978 378398 208046
rect 377778 207922 377874 207978
rect 377930 207922 377998 207978
rect 378054 207922 378122 207978
rect 378178 207922 378246 207978
rect 378302 207922 378398 207978
rect 377778 190350 378398 207922
rect 377778 190294 377874 190350
rect 377930 190294 377998 190350
rect 378054 190294 378122 190350
rect 378178 190294 378246 190350
rect 378302 190294 378398 190350
rect 377778 190226 378398 190294
rect 377778 190170 377874 190226
rect 377930 190170 377998 190226
rect 378054 190170 378122 190226
rect 378178 190170 378246 190226
rect 378302 190170 378398 190226
rect 377778 190102 378398 190170
rect 377778 190046 377874 190102
rect 377930 190046 377998 190102
rect 378054 190046 378122 190102
rect 378178 190046 378246 190102
rect 378302 190046 378398 190102
rect 377778 189978 378398 190046
rect 377778 189922 377874 189978
rect 377930 189922 377998 189978
rect 378054 189922 378122 189978
rect 378178 189922 378246 189978
rect 378302 189922 378398 189978
rect 377778 172350 378398 189922
rect 377778 172294 377874 172350
rect 377930 172294 377998 172350
rect 378054 172294 378122 172350
rect 378178 172294 378246 172350
rect 378302 172294 378398 172350
rect 377778 172226 378398 172294
rect 377778 172170 377874 172226
rect 377930 172170 377998 172226
rect 378054 172170 378122 172226
rect 378178 172170 378246 172226
rect 378302 172170 378398 172226
rect 377778 172102 378398 172170
rect 377778 172046 377874 172102
rect 377930 172046 377998 172102
rect 378054 172046 378122 172102
rect 378178 172046 378246 172102
rect 378302 172046 378398 172102
rect 377778 171978 378398 172046
rect 377778 171922 377874 171978
rect 377930 171922 377998 171978
rect 378054 171922 378122 171978
rect 378178 171922 378246 171978
rect 378302 171922 378398 171978
rect 375452 153906 375508 153916
rect 377778 154350 378398 171922
rect 377778 154294 377874 154350
rect 377930 154294 377998 154350
rect 378054 154294 378122 154350
rect 378178 154294 378246 154350
rect 378302 154294 378398 154350
rect 377778 154226 378398 154294
rect 377778 154170 377874 154226
rect 377930 154170 377998 154226
rect 378054 154170 378122 154226
rect 378178 154170 378246 154226
rect 378302 154170 378398 154226
rect 377778 154102 378398 154170
rect 377778 154046 377874 154102
rect 377930 154046 377998 154102
rect 378054 154046 378122 154102
rect 378178 154046 378246 154102
rect 378302 154046 378398 154102
rect 377778 153978 378398 154046
rect 377778 153922 377874 153978
rect 377930 153922 377998 153978
rect 378054 153922 378122 153978
rect 378178 153922 378246 153978
rect 378302 153922 378398 153978
rect 374058 148294 374154 148350
rect 374210 148294 374278 148350
rect 374334 148294 374402 148350
rect 374458 148294 374526 148350
rect 374582 148294 374678 148350
rect 374058 148226 374678 148294
rect 374058 148170 374154 148226
rect 374210 148170 374278 148226
rect 374334 148170 374402 148226
rect 374458 148170 374526 148226
rect 374582 148170 374678 148226
rect 374058 148102 374678 148170
rect 374058 148046 374154 148102
rect 374210 148046 374278 148102
rect 374334 148046 374402 148102
rect 374458 148046 374526 148102
rect 374582 148046 374678 148102
rect 374058 147978 374678 148046
rect 374058 147922 374154 147978
rect 374210 147922 374278 147978
rect 374334 147922 374402 147978
rect 374458 147922 374526 147978
rect 374582 147922 374678 147978
rect 374058 130350 374678 147922
rect 374058 130294 374154 130350
rect 374210 130294 374278 130350
rect 374334 130294 374402 130350
rect 374458 130294 374526 130350
rect 374582 130294 374678 130350
rect 374058 130226 374678 130294
rect 374058 130170 374154 130226
rect 374210 130170 374278 130226
rect 374334 130170 374402 130226
rect 374458 130170 374526 130226
rect 374582 130170 374678 130226
rect 374058 130102 374678 130170
rect 374058 130046 374154 130102
rect 374210 130046 374278 130102
rect 374334 130046 374402 130102
rect 374458 130046 374526 130102
rect 374582 130046 374678 130102
rect 374058 129978 374678 130046
rect 374058 129922 374154 129978
rect 374210 129922 374278 129978
rect 374334 129922 374402 129978
rect 374458 129922 374526 129978
rect 374582 129922 374678 129978
rect 374058 115262 374678 129922
rect 377778 136350 378398 153922
rect 380492 139300 380548 330876
rect 380492 139234 380548 139244
rect 382172 326452 382228 326462
rect 377778 136294 377874 136350
rect 377930 136294 377998 136350
rect 378054 136294 378122 136350
rect 378178 136294 378246 136350
rect 378302 136294 378398 136350
rect 377778 136226 378398 136294
rect 377778 136170 377874 136226
rect 377930 136170 377998 136226
rect 378054 136170 378122 136226
rect 378178 136170 378246 136226
rect 378302 136170 378398 136226
rect 377778 136102 378398 136170
rect 377778 136046 377874 136102
rect 377930 136046 377998 136102
rect 378054 136046 378122 136102
rect 378178 136046 378246 136102
rect 378302 136046 378398 136102
rect 377778 135978 378398 136046
rect 377778 135922 377874 135978
rect 377930 135922 377998 135978
rect 378054 135922 378122 135978
rect 378178 135922 378246 135978
rect 378302 135922 378398 135978
rect 377778 118350 378398 135922
rect 382172 127652 382228 326396
rect 383852 324212 383908 324222
rect 383068 309652 383124 309662
rect 383068 246820 383124 309596
rect 383068 246754 383124 246764
rect 382172 127586 382228 127596
rect 383852 121828 383908 324156
rect 383964 200116 384020 388682
rect 404778 382350 405398 399922
rect 404778 382294 404874 382350
rect 404930 382294 404998 382350
rect 405054 382294 405122 382350
rect 405178 382294 405246 382350
rect 405302 382294 405398 382350
rect 404778 382226 405398 382294
rect 404778 382170 404874 382226
rect 404930 382170 404998 382226
rect 405054 382170 405122 382226
rect 405178 382170 405246 382226
rect 405302 382170 405398 382226
rect 404778 382102 405398 382170
rect 404778 382046 404874 382102
rect 404930 382046 404998 382102
rect 405054 382046 405122 382102
rect 405178 382046 405246 382102
rect 405302 382046 405398 382102
rect 404778 381978 405398 382046
rect 404778 381922 404874 381978
rect 404930 381922 404998 381978
rect 405054 381922 405122 381978
rect 405178 381922 405246 381978
rect 405302 381922 405398 381978
rect 404778 364350 405398 381922
rect 404778 364294 404874 364350
rect 404930 364294 404998 364350
rect 405054 364294 405122 364350
rect 405178 364294 405246 364350
rect 405302 364294 405398 364350
rect 404778 364226 405398 364294
rect 404778 364170 404874 364226
rect 404930 364170 404998 364226
rect 405054 364170 405122 364226
rect 405178 364170 405246 364226
rect 405302 364170 405398 364226
rect 404778 364102 405398 364170
rect 404778 364046 404874 364102
rect 404930 364046 404998 364102
rect 405054 364046 405122 364102
rect 405178 364046 405246 364102
rect 405302 364046 405398 364102
rect 404778 363978 405398 364046
rect 404778 363922 404874 363978
rect 404930 363922 404998 363978
rect 405054 363922 405122 363978
rect 405178 363922 405246 363978
rect 405302 363922 405398 363978
rect 404778 346350 405398 363922
rect 404778 346294 404874 346350
rect 404930 346294 404998 346350
rect 405054 346294 405122 346350
rect 405178 346294 405246 346350
rect 405302 346294 405398 346350
rect 404778 346226 405398 346294
rect 404778 346170 404874 346226
rect 404930 346170 404998 346226
rect 405054 346170 405122 346226
rect 405178 346170 405246 346226
rect 405302 346170 405398 346226
rect 404778 346102 405398 346170
rect 404778 346046 404874 346102
rect 404930 346046 404998 346102
rect 405054 346046 405122 346102
rect 405178 346046 405246 346102
rect 405302 346046 405398 346102
rect 404778 345978 405398 346046
rect 404778 345922 404874 345978
rect 404930 345922 404998 345978
rect 405054 345922 405122 345978
rect 405178 345922 405246 345978
rect 405302 345922 405398 345978
rect 389116 344372 389172 344382
rect 388892 332052 388948 332062
rect 387212 329812 387268 329822
rect 385532 328692 385588 328702
rect 384748 308532 384804 308542
rect 384748 246708 384804 308476
rect 384748 246642 384804 246652
rect 383964 200050 384020 200060
rect 385532 133476 385588 328636
rect 387212 136388 387268 329756
rect 388892 142212 388948 331996
rect 389116 331828 389172 344316
rect 393932 334292 393988 334302
rect 389116 331762 389172 331772
rect 390572 333172 390628 333182
rect 390572 145124 390628 333116
rect 390572 145058 390628 145068
rect 392252 325332 392308 325342
rect 388892 142146 388948 142156
rect 387212 136322 387268 136332
rect 385532 133410 385588 133420
rect 392252 124740 392308 325276
rect 393932 152068 393988 334236
rect 404778 328350 405398 345922
rect 404778 328294 404874 328350
rect 404930 328294 404998 328350
rect 405054 328294 405122 328350
rect 405178 328294 405246 328350
rect 405302 328294 405398 328350
rect 404778 328226 405398 328294
rect 404778 328170 404874 328226
rect 404930 328170 404998 328226
rect 405054 328170 405122 328226
rect 405178 328170 405246 328226
rect 405302 328170 405398 328226
rect 404778 328102 405398 328170
rect 404778 328046 404874 328102
rect 404930 328046 404998 328102
rect 405054 328046 405122 328102
rect 405178 328046 405246 328102
rect 405302 328046 405398 328102
rect 404778 327978 405398 328046
rect 404778 327922 404874 327978
rect 404930 327922 404998 327978
rect 405054 327922 405122 327978
rect 405178 327922 405246 327978
rect 405302 327922 405398 327978
rect 404778 310350 405398 327922
rect 404778 310294 404874 310350
rect 404930 310294 404998 310350
rect 405054 310294 405122 310350
rect 405178 310294 405246 310350
rect 405302 310294 405398 310350
rect 404778 310226 405398 310294
rect 404778 310170 404874 310226
rect 404930 310170 404998 310226
rect 405054 310170 405122 310226
rect 405178 310170 405246 310226
rect 405302 310170 405398 310226
rect 404778 310102 405398 310170
rect 404778 310046 404874 310102
rect 404930 310046 404998 310102
rect 405054 310046 405122 310102
rect 405178 310046 405246 310102
rect 405302 310046 405398 310102
rect 404778 309978 405398 310046
rect 404778 309922 404874 309978
rect 404930 309922 404998 309978
rect 405054 309922 405122 309978
rect 405178 309922 405246 309978
rect 405302 309922 405398 309978
rect 404778 292350 405398 309922
rect 404778 292294 404874 292350
rect 404930 292294 404998 292350
rect 405054 292294 405122 292350
rect 405178 292294 405246 292350
rect 405302 292294 405398 292350
rect 404778 292226 405398 292294
rect 404778 292170 404874 292226
rect 404930 292170 404998 292226
rect 405054 292170 405122 292226
rect 405178 292170 405246 292226
rect 405302 292170 405398 292226
rect 404778 292102 405398 292170
rect 404778 292046 404874 292102
rect 404930 292046 404998 292102
rect 405054 292046 405122 292102
rect 405178 292046 405246 292102
rect 405302 292046 405398 292102
rect 404778 291978 405398 292046
rect 404778 291922 404874 291978
rect 404930 291922 404998 291978
rect 405054 291922 405122 291978
rect 405178 291922 405246 291978
rect 405302 291922 405398 291978
rect 404778 274350 405398 291922
rect 404778 274294 404874 274350
rect 404930 274294 404998 274350
rect 405054 274294 405122 274350
rect 405178 274294 405246 274350
rect 405302 274294 405398 274350
rect 404778 274226 405398 274294
rect 404778 274170 404874 274226
rect 404930 274170 404998 274226
rect 405054 274170 405122 274226
rect 405178 274170 405246 274226
rect 405302 274170 405398 274226
rect 404778 274102 405398 274170
rect 404778 274046 404874 274102
rect 404930 274046 404998 274102
rect 405054 274046 405122 274102
rect 405178 274046 405246 274102
rect 405302 274046 405398 274102
rect 404778 273978 405398 274046
rect 404778 273922 404874 273978
rect 404930 273922 404998 273978
rect 405054 273922 405122 273978
rect 405178 273922 405246 273978
rect 405302 273922 405398 273978
rect 404778 256350 405398 273922
rect 404778 256294 404874 256350
rect 404930 256294 404998 256350
rect 405054 256294 405122 256350
rect 405178 256294 405246 256350
rect 405302 256294 405398 256350
rect 404778 256226 405398 256294
rect 404778 256170 404874 256226
rect 404930 256170 404998 256226
rect 405054 256170 405122 256226
rect 405178 256170 405246 256226
rect 405302 256170 405398 256226
rect 404778 256102 405398 256170
rect 404778 256046 404874 256102
rect 404930 256046 404998 256102
rect 405054 256046 405122 256102
rect 405178 256046 405246 256102
rect 405302 256046 405398 256102
rect 404778 255978 405398 256046
rect 404778 255922 404874 255978
rect 404930 255922 404998 255978
rect 405054 255922 405122 255978
rect 405178 255922 405246 255978
rect 405302 255922 405398 255978
rect 393932 152002 393988 152012
rect 395612 246820 395668 246830
rect 395612 128548 395668 246764
rect 395612 128482 395668 128492
rect 404012 246372 404068 246382
rect 392252 124674 392308 124684
rect 383852 121762 383908 121772
rect 404012 120148 404068 246316
rect 404012 120082 404068 120092
rect 404778 238350 405398 255922
rect 404778 238294 404874 238350
rect 404930 238294 404998 238350
rect 405054 238294 405122 238350
rect 405178 238294 405246 238350
rect 405302 238294 405398 238350
rect 404778 238226 405398 238294
rect 404778 238170 404874 238226
rect 404930 238170 404998 238226
rect 405054 238170 405122 238226
rect 405178 238170 405246 238226
rect 405302 238170 405398 238226
rect 404778 238102 405398 238170
rect 404778 238046 404874 238102
rect 404930 238046 404998 238102
rect 405054 238046 405122 238102
rect 405178 238046 405246 238102
rect 405302 238046 405398 238102
rect 404778 237978 405398 238046
rect 404778 237922 404874 237978
rect 404930 237922 404998 237978
rect 405054 237922 405122 237978
rect 405178 237922 405246 237978
rect 405302 237922 405398 237978
rect 404778 220350 405398 237922
rect 404778 220294 404874 220350
rect 404930 220294 404998 220350
rect 405054 220294 405122 220350
rect 405178 220294 405246 220350
rect 405302 220294 405398 220350
rect 404778 220226 405398 220294
rect 404778 220170 404874 220226
rect 404930 220170 404998 220226
rect 405054 220170 405122 220226
rect 405178 220170 405246 220226
rect 405302 220170 405398 220226
rect 404778 220102 405398 220170
rect 404778 220046 404874 220102
rect 404930 220046 404998 220102
rect 405054 220046 405122 220102
rect 405178 220046 405246 220102
rect 405302 220046 405398 220102
rect 404778 219978 405398 220046
rect 404778 219922 404874 219978
rect 404930 219922 404998 219978
rect 405054 219922 405122 219978
rect 405178 219922 405246 219978
rect 405302 219922 405398 219978
rect 404778 202350 405398 219922
rect 404778 202294 404874 202350
rect 404930 202294 404998 202350
rect 405054 202294 405122 202350
rect 405178 202294 405246 202350
rect 405302 202294 405398 202350
rect 404778 202226 405398 202294
rect 404778 202170 404874 202226
rect 404930 202170 404998 202226
rect 405054 202170 405122 202226
rect 405178 202170 405246 202226
rect 405302 202170 405398 202226
rect 404778 202102 405398 202170
rect 404778 202046 404874 202102
rect 404930 202046 404998 202102
rect 405054 202046 405122 202102
rect 405178 202046 405246 202102
rect 405302 202046 405398 202102
rect 404778 201978 405398 202046
rect 404778 201922 404874 201978
rect 404930 201922 404998 201978
rect 405054 201922 405122 201978
rect 405178 201922 405246 201978
rect 405302 201922 405398 201978
rect 404778 184350 405398 201922
rect 404778 184294 404874 184350
rect 404930 184294 404998 184350
rect 405054 184294 405122 184350
rect 405178 184294 405246 184350
rect 405302 184294 405398 184350
rect 404778 184226 405398 184294
rect 404778 184170 404874 184226
rect 404930 184170 404998 184226
rect 405054 184170 405122 184226
rect 405178 184170 405246 184226
rect 405302 184170 405398 184226
rect 404778 184102 405398 184170
rect 404778 184046 404874 184102
rect 404930 184046 404998 184102
rect 405054 184046 405122 184102
rect 405178 184046 405246 184102
rect 405302 184046 405398 184102
rect 404778 183978 405398 184046
rect 404778 183922 404874 183978
rect 404930 183922 404998 183978
rect 405054 183922 405122 183978
rect 405178 183922 405246 183978
rect 405302 183922 405398 183978
rect 404778 166350 405398 183922
rect 404778 166294 404874 166350
rect 404930 166294 404998 166350
rect 405054 166294 405122 166350
rect 405178 166294 405246 166350
rect 405302 166294 405398 166350
rect 404778 166226 405398 166294
rect 404778 166170 404874 166226
rect 404930 166170 404998 166226
rect 405054 166170 405122 166226
rect 405178 166170 405246 166226
rect 405302 166170 405398 166226
rect 404778 166102 405398 166170
rect 404778 166046 404874 166102
rect 404930 166046 404998 166102
rect 405054 166046 405122 166102
rect 405178 166046 405246 166102
rect 405302 166046 405398 166102
rect 404778 165978 405398 166046
rect 404778 165922 404874 165978
rect 404930 165922 404998 165978
rect 405054 165922 405122 165978
rect 405178 165922 405246 165978
rect 405302 165922 405398 165978
rect 404778 148350 405398 165922
rect 404778 148294 404874 148350
rect 404930 148294 404998 148350
rect 405054 148294 405122 148350
rect 405178 148294 405246 148350
rect 405302 148294 405398 148350
rect 404778 148226 405398 148294
rect 404778 148170 404874 148226
rect 404930 148170 404998 148226
rect 405054 148170 405122 148226
rect 405178 148170 405246 148226
rect 405302 148170 405398 148226
rect 404778 148102 405398 148170
rect 404778 148046 404874 148102
rect 404930 148046 404998 148102
rect 405054 148046 405122 148102
rect 405178 148046 405246 148102
rect 405302 148046 405398 148102
rect 404778 147978 405398 148046
rect 404778 147922 404874 147978
rect 404930 147922 404998 147978
rect 405054 147922 405122 147978
rect 405178 147922 405246 147978
rect 405302 147922 405398 147978
rect 404778 130350 405398 147922
rect 404778 130294 404874 130350
rect 404930 130294 404998 130350
rect 405054 130294 405122 130350
rect 405178 130294 405246 130350
rect 405302 130294 405398 130350
rect 404778 130226 405398 130294
rect 404778 130170 404874 130226
rect 404930 130170 404998 130226
rect 405054 130170 405122 130226
rect 405178 130170 405246 130226
rect 405302 130170 405398 130226
rect 404778 130102 405398 130170
rect 404778 130046 404874 130102
rect 404930 130046 404998 130102
rect 405054 130046 405122 130102
rect 405178 130046 405246 130102
rect 405302 130046 405398 130102
rect 404778 129978 405398 130046
rect 404778 129922 404874 129978
rect 404930 129922 404998 129978
rect 405054 129922 405122 129978
rect 405178 129922 405246 129978
rect 405302 129922 405398 129978
rect 377778 118294 377874 118350
rect 377930 118294 377998 118350
rect 378054 118294 378122 118350
rect 378178 118294 378246 118350
rect 378302 118294 378398 118350
rect 377778 118226 378398 118294
rect 377778 118170 377874 118226
rect 377930 118170 377998 118226
rect 378054 118170 378122 118226
rect 378178 118170 378246 118226
rect 378302 118170 378398 118226
rect 377778 118102 378398 118170
rect 377778 118046 377874 118102
rect 377930 118046 377998 118102
rect 378054 118046 378122 118102
rect 378178 118046 378246 118102
rect 378302 118046 378398 118102
rect 377778 117978 378398 118046
rect 377778 117922 377874 117978
rect 377930 117922 377998 117978
rect 378054 117922 378122 117978
rect 378178 117922 378246 117978
rect 378302 117922 378398 117978
rect 377778 115262 378398 117922
rect 404778 115262 405398 129922
rect 408498 406350 409118 408578
rect 408498 406294 408594 406350
rect 408650 406294 408718 406350
rect 408774 406294 408842 406350
rect 408898 406294 408966 406350
rect 409022 406294 409118 406350
rect 408498 406226 409118 406294
rect 408498 406170 408594 406226
rect 408650 406170 408718 406226
rect 408774 406170 408842 406226
rect 408898 406170 408966 406226
rect 409022 406170 409118 406226
rect 408498 406102 409118 406170
rect 408498 406046 408594 406102
rect 408650 406046 408718 406102
rect 408774 406046 408842 406102
rect 408898 406046 408966 406102
rect 409022 406046 409118 406102
rect 408498 405978 409118 406046
rect 408498 405922 408594 405978
rect 408650 405922 408718 405978
rect 408774 405922 408842 405978
rect 408898 405922 408966 405978
rect 409022 405922 409118 405978
rect 408498 388350 409118 405922
rect 408498 388294 408594 388350
rect 408650 388294 408718 388350
rect 408774 388294 408842 388350
rect 408898 388294 408966 388350
rect 409022 388294 409118 388350
rect 408498 388226 409118 388294
rect 408498 388170 408594 388226
rect 408650 388170 408718 388226
rect 408774 388170 408842 388226
rect 408898 388170 408966 388226
rect 409022 388170 409118 388226
rect 408498 388102 409118 388170
rect 408498 388046 408594 388102
rect 408650 388046 408718 388102
rect 408774 388046 408842 388102
rect 408898 388046 408966 388102
rect 409022 388046 409118 388102
rect 408498 387978 409118 388046
rect 408498 387922 408594 387978
rect 408650 387922 408718 387978
rect 408774 387922 408842 387978
rect 408898 387922 408966 387978
rect 409022 387922 409118 387978
rect 408498 370350 409118 387922
rect 408498 370294 408594 370350
rect 408650 370294 408718 370350
rect 408774 370294 408842 370350
rect 408898 370294 408966 370350
rect 409022 370294 409118 370350
rect 408498 370226 409118 370294
rect 408498 370170 408594 370226
rect 408650 370170 408718 370226
rect 408774 370170 408842 370226
rect 408898 370170 408966 370226
rect 409022 370170 409118 370226
rect 408498 370102 409118 370170
rect 408498 370046 408594 370102
rect 408650 370046 408718 370102
rect 408774 370046 408842 370102
rect 408898 370046 408966 370102
rect 409022 370046 409118 370102
rect 408498 369978 409118 370046
rect 408498 369922 408594 369978
rect 408650 369922 408718 369978
rect 408774 369922 408842 369978
rect 408898 369922 408966 369978
rect 409022 369922 409118 369978
rect 408498 352350 409118 369922
rect 408498 352294 408594 352350
rect 408650 352294 408718 352350
rect 408774 352294 408842 352350
rect 408898 352294 408966 352350
rect 409022 352294 409118 352350
rect 408498 352226 409118 352294
rect 408498 352170 408594 352226
rect 408650 352170 408718 352226
rect 408774 352170 408842 352226
rect 408898 352170 408966 352226
rect 409022 352170 409118 352226
rect 408498 352102 409118 352170
rect 408498 352046 408594 352102
rect 408650 352046 408718 352102
rect 408774 352046 408842 352102
rect 408898 352046 408966 352102
rect 409022 352046 409118 352102
rect 408498 351978 409118 352046
rect 408498 351922 408594 351978
rect 408650 351922 408718 351978
rect 408774 351922 408842 351978
rect 408898 351922 408966 351978
rect 409022 351922 409118 351978
rect 408498 334350 409118 351922
rect 435498 400350 436118 408578
rect 435498 400294 435594 400350
rect 435650 400294 435718 400350
rect 435774 400294 435842 400350
rect 435898 400294 435966 400350
rect 436022 400294 436118 400350
rect 435498 400226 436118 400294
rect 435498 400170 435594 400226
rect 435650 400170 435718 400226
rect 435774 400170 435842 400226
rect 435898 400170 435966 400226
rect 436022 400170 436118 400226
rect 435498 400102 436118 400170
rect 435498 400046 435594 400102
rect 435650 400046 435718 400102
rect 435774 400046 435842 400102
rect 435898 400046 435966 400102
rect 436022 400046 436118 400102
rect 435498 399978 436118 400046
rect 435498 399922 435594 399978
rect 435650 399922 435718 399978
rect 435774 399922 435842 399978
rect 435898 399922 435966 399978
rect 436022 399922 436118 399978
rect 435498 382350 436118 399922
rect 435498 382294 435594 382350
rect 435650 382294 435718 382350
rect 435774 382294 435842 382350
rect 435898 382294 435966 382350
rect 436022 382294 436118 382350
rect 435498 382226 436118 382294
rect 435498 382170 435594 382226
rect 435650 382170 435718 382226
rect 435774 382170 435842 382226
rect 435898 382170 435966 382226
rect 436022 382170 436118 382226
rect 435498 382102 436118 382170
rect 435498 382046 435594 382102
rect 435650 382046 435718 382102
rect 435774 382046 435842 382102
rect 435898 382046 435966 382102
rect 436022 382046 436118 382102
rect 435498 381978 436118 382046
rect 435498 381922 435594 381978
rect 435650 381922 435718 381978
rect 435774 381922 435842 381978
rect 435898 381922 435966 381978
rect 436022 381922 436118 381978
rect 435498 364350 436118 381922
rect 435498 364294 435594 364350
rect 435650 364294 435718 364350
rect 435774 364294 435842 364350
rect 435898 364294 435966 364350
rect 436022 364294 436118 364350
rect 435498 364226 436118 364294
rect 435498 364170 435594 364226
rect 435650 364170 435718 364226
rect 435774 364170 435842 364226
rect 435898 364170 435966 364226
rect 436022 364170 436118 364226
rect 435498 364102 436118 364170
rect 435498 364046 435594 364102
rect 435650 364046 435718 364102
rect 435774 364046 435842 364102
rect 435898 364046 435966 364102
rect 436022 364046 436118 364102
rect 435498 363978 436118 364046
rect 435498 363922 435594 363978
rect 435650 363922 435718 363978
rect 435774 363922 435842 363978
rect 435898 363922 435966 363978
rect 436022 363922 436118 363978
rect 435498 346350 436118 363922
rect 435498 346294 435594 346350
rect 435650 346294 435718 346350
rect 435774 346294 435842 346350
rect 435898 346294 435966 346350
rect 436022 346294 436118 346350
rect 435498 346226 436118 346294
rect 435498 346170 435594 346226
rect 435650 346170 435718 346226
rect 435774 346170 435842 346226
rect 435898 346170 435966 346226
rect 436022 346170 436118 346226
rect 435498 346102 436118 346170
rect 435498 346046 435594 346102
rect 435650 346046 435718 346102
rect 435774 346046 435842 346102
rect 435898 346046 435966 346102
rect 436022 346046 436118 346102
rect 435498 345978 436118 346046
rect 435498 345922 435594 345978
rect 435650 345922 435718 345978
rect 435774 345922 435842 345978
rect 435898 345922 435966 345978
rect 436022 345922 436118 345978
rect 408498 334294 408594 334350
rect 408650 334294 408718 334350
rect 408774 334294 408842 334350
rect 408898 334294 408966 334350
rect 409022 334294 409118 334350
rect 408498 334226 409118 334294
rect 408498 334170 408594 334226
rect 408650 334170 408718 334226
rect 408774 334170 408842 334226
rect 408898 334170 408966 334226
rect 409022 334170 409118 334226
rect 408498 334102 409118 334170
rect 408498 334046 408594 334102
rect 408650 334046 408718 334102
rect 408774 334046 408842 334102
rect 408898 334046 408966 334102
rect 409022 334046 409118 334102
rect 408498 333978 409118 334046
rect 408498 333922 408594 333978
rect 408650 333922 408718 333978
rect 408774 333922 408842 333978
rect 408898 333922 408966 333978
rect 409022 333922 409118 333978
rect 408498 316350 409118 333922
rect 408498 316294 408594 316350
rect 408650 316294 408718 316350
rect 408774 316294 408842 316350
rect 408898 316294 408966 316350
rect 409022 316294 409118 316350
rect 408498 316226 409118 316294
rect 408498 316170 408594 316226
rect 408650 316170 408718 316226
rect 408774 316170 408842 316226
rect 408898 316170 408966 316226
rect 409022 316170 409118 316226
rect 408498 316102 409118 316170
rect 408498 316046 408594 316102
rect 408650 316046 408718 316102
rect 408774 316046 408842 316102
rect 408898 316046 408966 316102
rect 409022 316046 409118 316102
rect 408498 315978 409118 316046
rect 408498 315922 408594 315978
rect 408650 315922 408718 315978
rect 408774 315922 408842 315978
rect 408898 315922 408966 315978
rect 409022 315922 409118 315978
rect 408498 298350 409118 315922
rect 408498 298294 408594 298350
rect 408650 298294 408718 298350
rect 408774 298294 408842 298350
rect 408898 298294 408966 298350
rect 409022 298294 409118 298350
rect 408498 298226 409118 298294
rect 408498 298170 408594 298226
rect 408650 298170 408718 298226
rect 408774 298170 408842 298226
rect 408898 298170 408966 298226
rect 409022 298170 409118 298226
rect 408498 298102 409118 298170
rect 408498 298046 408594 298102
rect 408650 298046 408718 298102
rect 408774 298046 408842 298102
rect 408898 298046 408966 298102
rect 409022 298046 409118 298102
rect 408498 297978 409118 298046
rect 408498 297922 408594 297978
rect 408650 297922 408718 297978
rect 408774 297922 408842 297978
rect 408898 297922 408966 297978
rect 409022 297922 409118 297978
rect 408498 280350 409118 297922
rect 425852 337652 425908 337662
rect 408498 280294 408594 280350
rect 408650 280294 408718 280350
rect 408774 280294 408842 280350
rect 408898 280294 408966 280350
rect 409022 280294 409118 280350
rect 408498 280226 409118 280294
rect 408498 280170 408594 280226
rect 408650 280170 408718 280226
rect 408774 280170 408842 280226
rect 408898 280170 408966 280226
rect 409022 280170 409118 280226
rect 408498 280102 409118 280170
rect 408498 280046 408594 280102
rect 408650 280046 408718 280102
rect 408774 280046 408842 280102
rect 408898 280046 408966 280102
rect 409022 280046 409118 280102
rect 408498 279978 409118 280046
rect 408498 279922 408594 279978
rect 408650 279922 408718 279978
rect 408774 279922 408842 279978
rect 408898 279922 408966 279978
rect 409022 279922 409118 279978
rect 408498 262350 409118 279922
rect 411740 289492 411796 289502
rect 408498 262294 408594 262350
rect 408650 262294 408718 262350
rect 408774 262294 408842 262350
rect 408898 262294 408966 262350
rect 409022 262294 409118 262350
rect 408498 262226 409118 262294
rect 408498 262170 408594 262226
rect 408650 262170 408718 262226
rect 408774 262170 408842 262226
rect 408898 262170 408966 262226
rect 409022 262170 409118 262226
rect 408498 262102 409118 262170
rect 408498 262046 408594 262102
rect 408650 262046 408718 262102
rect 408774 262046 408842 262102
rect 408898 262046 408966 262102
rect 409022 262046 409118 262102
rect 408498 261978 409118 262046
rect 408498 261922 408594 261978
rect 408650 261922 408718 261978
rect 408774 261922 408842 261978
rect 408898 261922 408966 261978
rect 409022 261922 409118 261978
rect 408498 244350 409118 261922
rect 408498 244294 408594 244350
rect 408650 244294 408718 244350
rect 408774 244294 408842 244350
rect 408898 244294 408966 244350
rect 409022 244294 409118 244350
rect 408498 244226 409118 244294
rect 408498 244170 408594 244226
rect 408650 244170 408718 244226
rect 408774 244170 408842 244226
rect 408898 244170 408966 244226
rect 409022 244170 409118 244226
rect 408498 244102 409118 244170
rect 408498 244046 408594 244102
rect 408650 244046 408718 244102
rect 408774 244046 408842 244102
rect 408898 244046 408966 244102
rect 409022 244046 409118 244102
rect 408498 243978 409118 244046
rect 408498 243922 408594 243978
rect 408650 243922 408718 243978
rect 408774 243922 408842 243978
rect 408898 243922 408966 243978
rect 409022 243922 409118 243978
rect 408498 226350 409118 243922
rect 408498 226294 408594 226350
rect 408650 226294 408718 226350
rect 408774 226294 408842 226350
rect 408898 226294 408966 226350
rect 409022 226294 409118 226350
rect 408498 226226 409118 226294
rect 408498 226170 408594 226226
rect 408650 226170 408718 226226
rect 408774 226170 408842 226226
rect 408898 226170 408966 226226
rect 409022 226170 409118 226226
rect 408498 226102 409118 226170
rect 408498 226046 408594 226102
rect 408650 226046 408718 226102
rect 408774 226046 408842 226102
rect 408898 226046 408966 226102
rect 409022 226046 409118 226102
rect 408498 225978 409118 226046
rect 408498 225922 408594 225978
rect 408650 225922 408718 225978
rect 408774 225922 408842 225978
rect 408898 225922 408966 225978
rect 409022 225922 409118 225978
rect 408498 208350 409118 225922
rect 408498 208294 408594 208350
rect 408650 208294 408718 208350
rect 408774 208294 408842 208350
rect 408898 208294 408966 208350
rect 409022 208294 409118 208350
rect 408498 208226 409118 208294
rect 408498 208170 408594 208226
rect 408650 208170 408718 208226
rect 408774 208170 408842 208226
rect 408898 208170 408966 208226
rect 409022 208170 409118 208226
rect 408498 208102 409118 208170
rect 408498 208046 408594 208102
rect 408650 208046 408718 208102
rect 408774 208046 408842 208102
rect 408898 208046 408966 208102
rect 409022 208046 409118 208102
rect 408498 207978 409118 208046
rect 408498 207922 408594 207978
rect 408650 207922 408718 207978
rect 408774 207922 408842 207978
rect 408898 207922 408966 207978
rect 409022 207922 409118 207978
rect 408498 190350 409118 207922
rect 408498 190294 408594 190350
rect 408650 190294 408718 190350
rect 408774 190294 408842 190350
rect 408898 190294 408966 190350
rect 409022 190294 409118 190350
rect 408498 190226 409118 190294
rect 408498 190170 408594 190226
rect 408650 190170 408718 190226
rect 408774 190170 408842 190226
rect 408898 190170 408966 190226
rect 409022 190170 409118 190226
rect 408498 190102 409118 190170
rect 408498 190046 408594 190102
rect 408650 190046 408718 190102
rect 408774 190046 408842 190102
rect 408898 190046 408966 190102
rect 409022 190046 409118 190102
rect 408498 189978 409118 190046
rect 408498 189922 408594 189978
rect 408650 189922 408718 189978
rect 408774 189922 408842 189978
rect 408898 189922 408966 189978
rect 409022 189922 409118 189978
rect 408498 172350 409118 189922
rect 408498 172294 408594 172350
rect 408650 172294 408718 172350
rect 408774 172294 408842 172350
rect 408898 172294 408966 172350
rect 409022 172294 409118 172350
rect 408498 172226 409118 172294
rect 408498 172170 408594 172226
rect 408650 172170 408718 172226
rect 408774 172170 408842 172226
rect 408898 172170 408966 172226
rect 409022 172170 409118 172226
rect 408498 172102 409118 172170
rect 408498 172046 408594 172102
rect 408650 172046 408718 172102
rect 408774 172046 408842 172102
rect 408898 172046 408966 172102
rect 409022 172046 409118 172102
rect 408498 171978 409118 172046
rect 408498 171922 408594 171978
rect 408650 171922 408718 171978
rect 408774 171922 408842 171978
rect 408898 171922 408966 171978
rect 409022 171922 409118 171978
rect 408498 154350 409118 171922
rect 408498 154294 408594 154350
rect 408650 154294 408718 154350
rect 408774 154294 408842 154350
rect 408898 154294 408966 154350
rect 409022 154294 409118 154350
rect 408498 154226 409118 154294
rect 408498 154170 408594 154226
rect 408650 154170 408718 154226
rect 408774 154170 408842 154226
rect 408898 154170 408966 154226
rect 409022 154170 409118 154226
rect 408498 154102 409118 154170
rect 408498 154046 408594 154102
rect 408650 154046 408718 154102
rect 408774 154046 408842 154102
rect 408898 154046 408966 154102
rect 409022 154046 409118 154102
rect 408498 153978 409118 154046
rect 408498 153922 408594 153978
rect 408650 153922 408718 153978
rect 408774 153922 408842 153978
rect 408898 153922 408966 153978
rect 409022 153922 409118 153978
rect 408498 136350 409118 153922
rect 408498 136294 408594 136350
rect 408650 136294 408718 136350
rect 408774 136294 408842 136350
rect 408898 136294 408966 136350
rect 409022 136294 409118 136350
rect 408498 136226 409118 136294
rect 408498 136170 408594 136226
rect 408650 136170 408718 136226
rect 408774 136170 408842 136226
rect 408898 136170 408966 136226
rect 409022 136170 409118 136226
rect 408498 136102 409118 136170
rect 408498 136046 408594 136102
rect 408650 136046 408718 136102
rect 408774 136046 408842 136102
rect 408898 136046 408966 136102
rect 409022 136046 409118 136102
rect 408498 135978 409118 136046
rect 408498 135922 408594 135978
rect 408650 135922 408718 135978
rect 408774 135922 408842 135978
rect 408898 135922 408966 135978
rect 409022 135922 409118 135978
rect 408498 118350 409118 135922
rect 408498 118294 408594 118350
rect 408650 118294 408718 118350
rect 408774 118294 408842 118350
rect 408898 118294 408966 118350
rect 409022 118294 409118 118350
rect 408498 118226 409118 118294
rect 408498 118170 408594 118226
rect 408650 118170 408718 118226
rect 408774 118170 408842 118226
rect 408898 118170 408966 118226
rect 409022 118170 409118 118226
rect 408498 118102 409118 118170
rect 408498 118046 408594 118102
rect 408650 118046 408718 118102
rect 408774 118046 408842 118102
rect 408898 118046 408966 118102
rect 409022 118046 409118 118102
rect 408498 117978 409118 118046
rect 408498 117922 408594 117978
rect 408650 117922 408718 117978
rect 408774 117922 408842 117978
rect 408898 117922 408966 117978
rect 409022 117922 409118 117978
rect 408498 115262 409118 117922
rect 411628 278292 411684 278302
rect 364448 112350 364768 112384
rect 364448 112294 364518 112350
rect 364574 112294 364642 112350
rect 364698 112294 364768 112350
rect 364448 112226 364768 112294
rect 364448 112170 364518 112226
rect 364574 112170 364642 112226
rect 364698 112170 364768 112226
rect 364448 112102 364768 112170
rect 364448 112046 364518 112102
rect 364574 112046 364642 112102
rect 364698 112046 364768 112102
rect 364448 111978 364768 112046
rect 364448 111922 364518 111978
rect 364574 111922 364642 111978
rect 364698 111922 364768 111978
rect 364448 111888 364768 111922
rect 395168 112350 395488 112384
rect 395168 112294 395238 112350
rect 395294 112294 395362 112350
rect 395418 112294 395488 112350
rect 395168 112226 395488 112294
rect 395168 112170 395238 112226
rect 395294 112170 395362 112226
rect 395418 112170 395488 112226
rect 395168 112102 395488 112170
rect 395168 112046 395238 112102
rect 395294 112046 395362 112102
rect 395418 112046 395488 112102
rect 395168 111978 395488 112046
rect 395168 111922 395238 111978
rect 395294 111922 395362 111978
rect 395418 111922 395488 111978
rect 395168 111888 395488 111922
rect 379808 100350 380128 100384
rect 379808 100294 379878 100350
rect 379934 100294 380002 100350
rect 380058 100294 380128 100350
rect 379808 100226 380128 100294
rect 379808 100170 379878 100226
rect 379934 100170 380002 100226
rect 380058 100170 380128 100226
rect 379808 100102 380128 100170
rect 379808 100046 379878 100102
rect 379934 100046 380002 100102
rect 380058 100046 380128 100102
rect 379808 99978 380128 100046
rect 379808 99922 379878 99978
rect 379934 99922 380002 99978
rect 380058 99922 380128 99978
rect 379808 99888 380128 99922
rect 410528 100350 410848 100384
rect 410528 100294 410598 100350
rect 410654 100294 410722 100350
rect 410778 100294 410848 100350
rect 410528 100226 410848 100294
rect 410528 100170 410598 100226
rect 410654 100170 410722 100226
rect 410778 100170 410848 100226
rect 410528 100102 410848 100170
rect 410528 100046 410598 100102
rect 410654 100046 410722 100102
rect 410778 100046 410848 100102
rect 410528 99978 410848 100046
rect 410528 99922 410598 99978
rect 410654 99922 410722 99978
rect 410778 99922 410848 99978
rect 410528 99888 410848 99922
rect 364448 94350 364768 94384
rect 364448 94294 364518 94350
rect 364574 94294 364642 94350
rect 364698 94294 364768 94350
rect 364448 94226 364768 94294
rect 364448 94170 364518 94226
rect 364574 94170 364642 94226
rect 364698 94170 364768 94226
rect 364448 94102 364768 94170
rect 364448 94046 364518 94102
rect 364574 94046 364642 94102
rect 364698 94046 364768 94102
rect 364448 93978 364768 94046
rect 364448 93922 364518 93978
rect 364574 93922 364642 93978
rect 364698 93922 364768 93978
rect 364448 93888 364768 93922
rect 395168 94350 395488 94384
rect 395168 94294 395238 94350
rect 395294 94294 395362 94350
rect 395418 94294 395488 94350
rect 395168 94226 395488 94294
rect 395168 94170 395238 94226
rect 395294 94170 395362 94226
rect 395418 94170 395488 94226
rect 395168 94102 395488 94170
rect 395168 94046 395238 94102
rect 395294 94046 395362 94102
rect 395418 94046 395488 94102
rect 395168 93978 395488 94046
rect 395168 93922 395238 93978
rect 395294 93922 395362 93978
rect 395418 93922 395488 93978
rect 395168 93888 395488 93922
rect 379808 82350 380128 82384
rect 379808 82294 379878 82350
rect 379934 82294 380002 82350
rect 380058 82294 380128 82350
rect 379808 82226 380128 82294
rect 379808 82170 379878 82226
rect 379934 82170 380002 82226
rect 380058 82170 380128 82226
rect 379808 82102 380128 82170
rect 379808 82046 379878 82102
rect 379934 82046 380002 82102
rect 380058 82046 380128 82102
rect 379808 81978 380128 82046
rect 379808 81922 379878 81978
rect 379934 81922 380002 81978
rect 380058 81922 380128 81978
rect 379808 81888 380128 81922
rect 410528 82350 410848 82384
rect 410528 82294 410598 82350
rect 410654 82294 410722 82350
rect 410778 82294 410848 82350
rect 410528 82226 410848 82294
rect 410528 82170 410598 82226
rect 410654 82170 410722 82226
rect 410778 82170 410848 82226
rect 410528 82102 410848 82170
rect 410528 82046 410598 82102
rect 410654 82046 410722 82102
rect 410778 82046 410848 82102
rect 410528 81978 410848 82046
rect 410528 81922 410598 81978
rect 410654 81922 410722 81978
rect 410778 81922 410848 81978
rect 410528 81888 410848 81922
rect 364448 76350 364768 76384
rect 364448 76294 364518 76350
rect 364574 76294 364642 76350
rect 364698 76294 364768 76350
rect 364448 76226 364768 76294
rect 364448 76170 364518 76226
rect 364574 76170 364642 76226
rect 364698 76170 364768 76226
rect 364448 76102 364768 76170
rect 364448 76046 364518 76102
rect 364574 76046 364642 76102
rect 364698 76046 364768 76102
rect 364448 75978 364768 76046
rect 364448 75922 364518 75978
rect 364574 75922 364642 75978
rect 364698 75922 364768 75978
rect 364448 75888 364768 75922
rect 395168 76350 395488 76384
rect 395168 76294 395238 76350
rect 395294 76294 395362 76350
rect 395418 76294 395488 76350
rect 395168 76226 395488 76294
rect 395168 76170 395238 76226
rect 395294 76170 395362 76226
rect 395418 76170 395488 76226
rect 395168 76102 395488 76170
rect 395168 76046 395238 76102
rect 395294 76046 395362 76102
rect 395418 76046 395488 76102
rect 395168 75978 395488 76046
rect 395168 75922 395238 75978
rect 395294 75922 395362 75978
rect 395418 75922 395488 75978
rect 395168 75888 395488 75922
rect 379808 64350 380128 64384
rect 379808 64294 379878 64350
rect 379934 64294 380002 64350
rect 380058 64294 380128 64350
rect 379808 64226 380128 64294
rect 379808 64170 379878 64226
rect 379934 64170 380002 64226
rect 380058 64170 380128 64226
rect 379808 64102 380128 64170
rect 379808 64046 379878 64102
rect 379934 64046 380002 64102
rect 380058 64046 380128 64102
rect 379808 63978 380128 64046
rect 379808 63922 379878 63978
rect 379934 63922 380002 63978
rect 380058 63922 380128 63978
rect 379808 63888 380128 63922
rect 410528 64350 410848 64384
rect 410528 64294 410598 64350
rect 410654 64294 410722 64350
rect 410778 64294 410848 64350
rect 410528 64226 410848 64294
rect 410528 64170 410598 64226
rect 410654 64170 410722 64226
rect 410778 64170 410848 64226
rect 410528 64102 410848 64170
rect 410528 64046 410598 64102
rect 410654 64046 410722 64102
rect 410778 64046 410848 64102
rect 410528 63978 410848 64046
rect 410528 63922 410598 63978
rect 410654 63922 410722 63978
rect 410778 63922 410848 63978
rect 410528 63888 410848 63922
rect 364448 58350 364768 58384
rect 364448 58294 364518 58350
rect 364574 58294 364642 58350
rect 364698 58294 364768 58350
rect 364448 58226 364768 58294
rect 364448 58170 364518 58226
rect 364574 58170 364642 58226
rect 364698 58170 364768 58226
rect 364448 58102 364768 58170
rect 364448 58046 364518 58102
rect 364574 58046 364642 58102
rect 364698 58046 364768 58102
rect 364448 57978 364768 58046
rect 364448 57922 364518 57978
rect 364574 57922 364642 57978
rect 364698 57922 364768 57978
rect 364448 57888 364768 57922
rect 395168 58350 395488 58384
rect 395168 58294 395238 58350
rect 395294 58294 395362 58350
rect 395418 58294 395488 58350
rect 395168 58226 395488 58294
rect 395168 58170 395238 58226
rect 395294 58170 395362 58226
rect 395418 58170 395488 58226
rect 395168 58102 395488 58170
rect 395168 58046 395238 58102
rect 395294 58046 395362 58102
rect 395418 58046 395488 58102
rect 395168 57978 395488 58046
rect 395168 57922 395238 57978
rect 395294 57922 395362 57978
rect 395418 57922 395488 57978
rect 395168 57888 395488 57922
rect 362124 49522 362180 49532
rect 362012 41234 362068 41244
rect 358764 38098 358820 38108
rect 374058 40350 374678 53730
rect 374058 40294 374154 40350
rect 374210 40294 374278 40350
rect 374334 40294 374402 40350
rect 374458 40294 374526 40350
rect 374582 40294 374678 40350
rect 374058 40226 374678 40294
rect 374058 40170 374154 40226
rect 374210 40170 374278 40226
rect 374334 40170 374402 40226
rect 374458 40170 374526 40226
rect 374582 40170 374678 40226
rect 374058 40102 374678 40170
rect 374058 40046 374154 40102
rect 374210 40046 374278 40102
rect 374334 40046 374402 40102
rect 374458 40046 374526 40102
rect 374582 40046 374678 40102
rect 374058 39978 374678 40046
rect 374058 39922 374154 39978
rect 374210 39922 374278 39978
rect 374334 39922 374402 39978
rect 374458 39922 374526 39978
rect 374582 39922 374678 39978
rect 348572 4722 348628 4732
rect 374058 22350 374678 39922
rect 374058 22294 374154 22350
rect 374210 22294 374278 22350
rect 374334 22294 374402 22350
rect 374458 22294 374526 22350
rect 374582 22294 374678 22350
rect 374058 22226 374678 22294
rect 374058 22170 374154 22226
rect 374210 22170 374278 22226
rect 374334 22170 374402 22226
rect 374458 22170 374526 22226
rect 374582 22170 374678 22226
rect 374058 22102 374678 22170
rect 374058 22046 374154 22102
rect 374210 22046 374278 22102
rect 374334 22046 374402 22102
rect 374458 22046 374526 22102
rect 374582 22046 374678 22102
rect 374058 21978 374678 22046
rect 374058 21922 374154 21978
rect 374210 21922 374278 21978
rect 374334 21922 374402 21978
rect 374458 21922 374526 21978
rect 374582 21922 374678 21978
rect 347058 -1176 347154 -1120
rect 347210 -1176 347278 -1120
rect 347334 -1176 347402 -1120
rect 347458 -1176 347526 -1120
rect 347582 -1176 347678 -1120
rect 347058 -1244 347678 -1176
rect 347058 -1300 347154 -1244
rect 347210 -1300 347278 -1244
rect 347334 -1300 347402 -1244
rect 347458 -1300 347526 -1244
rect 347582 -1300 347678 -1244
rect 347058 -1368 347678 -1300
rect 347058 -1424 347154 -1368
rect 347210 -1424 347278 -1368
rect 347334 -1424 347402 -1368
rect 347458 -1424 347526 -1368
rect 347582 -1424 347678 -1368
rect 347058 -1492 347678 -1424
rect 347058 -1548 347154 -1492
rect 347210 -1548 347278 -1492
rect 347334 -1548 347402 -1492
rect 347458 -1548 347526 -1492
rect 347582 -1548 347678 -1492
rect 347058 -1644 347678 -1548
rect 374058 4350 374678 21922
rect 374058 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 374678 4350
rect 374058 4226 374678 4294
rect 374058 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 374678 4226
rect 374058 4102 374678 4170
rect 374058 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 374678 4102
rect 374058 3978 374678 4046
rect 374058 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 374678 3978
rect 374058 -160 374678 3922
rect 374058 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 374678 -160
rect 374058 -284 374678 -216
rect 374058 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 374678 -284
rect 374058 -408 374678 -340
rect 374058 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 374678 -408
rect 374058 -532 374678 -464
rect 374058 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 374678 -532
rect 374058 -1644 374678 -588
rect 377778 46350 378398 53730
rect 377778 46294 377874 46350
rect 377930 46294 377998 46350
rect 378054 46294 378122 46350
rect 378178 46294 378246 46350
rect 378302 46294 378398 46350
rect 377778 46226 378398 46294
rect 377778 46170 377874 46226
rect 377930 46170 377998 46226
rect 378054 46170 378122 46226
rect 378178 46170 378246 46226
rect 378302 46170 378398 46226
rect 377778 46102 378398 46170
rect 377778 46046 377874 46102
rect 377930 46046 377998 46102
rect 378054 46046 378122 46102
rect 378178 46046 378246 46102
rect 378302 46046 378398 46102
rect 377778 45978 378398 46046
rect 377778 45922 377874 45978
rect 377930 45922 377998 45978
rect 378054 45922 378122 45978
rect 378178 45922 378246 45978
rect 378302 45922 378398 45978
rect 377778 28350 378398 45922
rect 377778 28294 377874 28350
rect 377930 28294 377998 28350
rect 378054 28294 378122 28350
rect 378178 28294 378246 28350
rect 378302 28294 378398 28350
rect 377778 28226 378398 28294
rect 377778 28170 377874 28226
rect 377930 28170 377998 28226
rect 378054 28170 378122 28226
rect 378178 28170 378246 28226
rect 378302 28170 378398 28226
rect 377778 28102 378398 28170
rect 377778 28046 377874 28102
rect 377930 28046 377998 28102
rect 378054 28046 378122 28102
rect 378178 28046 378246 28102
rect 378302 28046 378398 28102
rect 377778 27978 378398 28046
rect 377778 27922 377874 27978
rect 377930 27922 377998 27978
rect 378054 27922 378122 27978
rect 378178 27922 378246 27978
rect 378302 27922 378398 27978
rect 377778 10350 378398 27922
rect 377778 10294 377874 10350
rect 377930 10294 377998 10350
rect 378054 10294 378122 10350
rect 378178 10294 378246 10350
rect 378302 10294 378398 10350
rect 377778 10226 378398 10294
rect 377778 10170 377874 10226
rect 377930 10170 377998 10226
rect 378054 10170 378122 10226
rect 378178 10170 378246 10226
rect 378302 10170 378398 10226
rect 377778 10102 378398 10170
rect 377778 10046 377874 10102
rect 377930 10046 377998 10102
rect 378054 10046 378122 10102
rect 378178 10046 378246 10102
rect 378302 10046 378398 10102
rect 377778 9978 378398 10046
rect 377778 9922 377874 9978
rect 377930 9922 377998 9978
rect 378054 9922 378122 9978
rect 378178 9922 378246 9978
rect 378302 9922 378398 9978
rect 377778 -1120 378398 9922
rect 377778 -1176 377874 -1120
rect 377930 -1176 377998 -1120
rect 378054 -1176 378122 -1120
rect 378178 -1176 378246 -1120
rect 378302 -1176 378398 -1120
rect 377778 -1244 378398 -1176
rect 377778 -1300 377874 -1244
rect 377930 -1300 377998 -1244
rect 378054 -1300 378122 -1244
rect 378178 -1300 378246 -1244
rect 378302 -1300 378398 -1244
rect 377778 -1368 378398 -1300
rect 377778 -1424 377874 -1368
rect 377930 -1424 377998 -1368
rect 378054 -1424 378122 -1368
rect 378178 -1424 378246 -1368
rect 378302 -1424 378398 -1368
rect 377778 -1492 378398 -1424
rect 377778 -1548 377874 -1492
rect 377930 -1548 377998 -1492
rect 378054 -1548 378122 -1492
rect 378178 -1548 378246 -1492
rect 378302 -1548 378398 -1492
rect 377778 -1644 378398 -1548
rect 404778 40350 405398 53730
rect 404778 40294 404874 40350
rect 404930 40294 404998 40350
rect 405054 40294 405122 40350
rect 405178 40294 405246 40350
rect 405302 40294 405398 40350
rect 404778 40226 405398 40294
rect 404778 40170 404874 40226
rect 404930 40170 404998 40226
rect 405054 40170 405122 40226
rect 405178 40170 405246 40226
rect 405302 40170 405398 40226
rect 404778 40102 405398 40170
rect 404778 40046 404874 40102
rect 404930 40046 404998 40102
rect 405054 40046 405122 40102
rect 405178 40046 405246 40102
rect 405302 40046 405398 40102
rect 404778 39978 405398 40046
rect 404778 39922 404874 39978
rect 404930 39922 404998 39978
rect 405054 39922 405122 39978
rect 405178 39922 405246 39978
rect 405302 39922 405398 39978
rect 404778 22350 405398 39922
rect 404778 22294 404874 22350
rect 404930 22294 404998 22350
rect 405054 22294 405122 22350
rect 405178 22294 405246 22350
rect 405302 22294 405398 22350
rect 404778 22226 405398 22294
rect 404778 22170 404874 22226
rect 404930 22170 404998 22226
rect 405054 22170 405122 22226
rect 405178 22170 405246 22226
rect 405302 22170 405398 22226
rect 404778 22102 405398 22170
rect 404778 22046 404874 22102
rect 404930 22046 404998 22102
rect 405054 22046 405122 22102
rect 405178 22046 405246 22102
rect 405302 22046 405398 22102
rect 404778 21978 405398 22046
rect 404778 21922 404874 21978
rect 404930 21922 404998 21978
rect 405054 21922 405122 21978
rect 405178 21922 405246 21978
rect 405302 21922 405398 21978
rect 404778 4350 405398 21922
rect 404778 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 405398 4350
rect 404778 4226 405398 4294
rect 404778 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 405398 4226
rect 404778 4102 405398 4170
rect 404778 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 405398 4102
rect 404778 3978 405398 4046
rect 404778 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 405398 3978
rect 404778 -160 405398 3922
rect 404778 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 405398 -160
rect 404778 -284 405398 -216
rect 404778 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 405398 -284
rect 404778 -408 405398 -340
rect 404778 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 405398 -408
rect 404778 -532 405398 -464
rect 404778 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 405398 -532
rect 404778 -1644 405398 -588
rect 408498 46350 409118 53730
rect 408498 46294 408594 46350
rect 408650 46294 408718 46350
rect 408774 46294 408842 46350
rect 408898 46294 408966 46350
rect 409022 46294 409118 46350
rect 408498 46226 409118 46294
rect 408498 46170 408594 46226
rect 408650 46170 408718 46226
rect 408774 46170 408842 46226
rect 408898 46170 408966 46226
rect 409022 46170 409118 46226
rect 408498 46102 409118 46170
rect 408498 46046 408594 46102
rect 408650 46046 408718 46102
rect 408774 46046 408842 46102
rect 408898 46046 408966 46102
rect 409022 46046 409118 46102
rect 408498 45978 409118 46046
rect 408498 45922 408594 45978
rect 408650 45922 408718 45978
rect 408774 45922 408842 45978
rect 408898 45922 408966 45978
rect 409022 45922 409118 45978
rect 408498 28350 409118 45922
rect 408498 28294 408594 28350
rect 408650 28294 408718 28350
rect 408774 28294 408842 28350
rect 408898 28294 408966 28350
rect 409022 28294 409118 28350
rect 408498 28226 409118 28294
rect 408498 28170 408594 28226
rect 408650 28170 408718 28226
rect 408774 28170 408842 28226
rect 408898 28170 408966 28226
rect 409022 28170 409118 28226
rect 408498 28102 409118 28170
rect 408498 28046 408594 28102
rect 408650 28046 408718 28102
rect 408774 28046 408842 28102
rect 408898 28046 408966 28102
rect 409022 28046 409118 28102
rect 408498 27978 409118 28046
rect 408498 27922 408594 27978
rect 408650 27922 408718 27978
rect 408774 27922 408842 27978
rect 408898 27922 408966 27978
rect 409022 27922 409118 27978
rect 408498 10350 409118 27922
rect 408498 10294 408594 10350
rect 408650 10294 408718 10350
rect 408774 10294 408842 10350
rect 408898 10294 408966 10350
rect 409022 10294 409118 10350
rect 408498 10226 409118 10294
rect 408498 10170 408594 10226
rect 408650 10170 408718 10226
rect 408774 10170 408842 10226
rect 408898 10170 408966 10226
rect 409022 10170 409118 10226
rect 408498 10102 409118 10170
rect 408498 10046 408594 10102
rect 408650 10046 408718 10102
rect 408774 10046 408842 10102
rect 408898 10046 408966 10102
rect 409022 10046 409118 10102
rect 408498 9978 409118 10046
rect 408498 9922 408594 9978
rect 408650 9922 408718 9978
rect 408774 9922 408842 9978
rect 408898 9922 408966 9978
rect 409022 9922 409118 9978
rect 408498 -1120 409118 9922
rect 411628 9268 411684 278236
rect 411740 42868 411796 289436
rect 424172 284004 424228 284014
rect 420812 280644 420868 280654
rect 411740 42802 411796 42812
rect 411852 272692 411908 272702
rect 411852 32788 411908 272636
rect 419356 263844 419412 263854
rect 419356 116116 419412 263788
rect 419356 116050 419412 116060
rect 420812 86884 420868 280588
rect 422492 260484 422548 260494
rect 422492 235172 422548 260428
rect 422492 235106 422548 235116
rect 423276 235172 423332 235182
rect 423276 234612 423332 235116
rect 423276 109172 423332 234556
rect 423276 109106 423332 109116
rect 424172 89796 424228 283948
rect 424172 89730 424228 89740
rect 420812 86818 420868 86828
rect 419244 52948 419300 52958
rect 419244 52052 419300 52892
rect 419244 51986 419300 51996
rect 425852 50372 425908 337596
rect 435498 328350 436118 345922
rect 435498 328294 435594 328350
rect 435650 328294 435718 328350
rect 435774 328294 435842 328350
rect 435898 328294 435966 328350
rect 436022 328294 436118 328350
rect 435498 328226 436118 328294
rect 435498 328170 435594 328226
rect 435650 328170 435718 328226
rect 435774 328170 435842 328226
rect 435898 328170 435966 328226
rect 436022 328170 436118 328226
rect 435498 328102 436118 328170
rect 435498 328046 435594 328102
rect 435650 328046 435718 328102
rect 435774 328046 435842 328102
rect 435898 328046 435966 328102
rect 436022 328046 436118 328102
rect 435498 327978 436118 328046
rect 435498 327922 435594 327978
rect 435650 327922 435718 327978
rect 435774 327922 435842 327978
rect 435898 327922 435966 327978
rect 436022 327922 436118 327978
rect 434252 319732 434308 319742
rect 432572 318388 432628 318398
rect 427532 316708 427588 316718
rect 425964 313460 426020 313470
rect 425964 92708 426020 313404
rect 427532 101444 427588 316652
rect 430892 315140 430948 315150
rect 429212 315028 429268 315038
rect 427532 101378 427588 101388
rect 427644 109172 427700 109182
rect 425964 92642 426020 92652
rect 427644 59668 427700 109116
rect 429212 98532 429268 314972
rect 430892 104356 430948 315084
rect 432572 107268 432628 318332
rect 434252 110180 434308 319676
rect 434252 110114 434308 110124
rect 435498 310350 436118 327922
rect 439218 406350 439838 408578
rect 439218 406294 439314 406350
rect 439370 406294 439438 406350
rect 439494 406294 439562 406350
rect 439618 406294 439686 406350
rect 439742 406294 439838 406350
rect 439218 406226 439838 406294
rect 439218 406170 439314 406226
rect 439370 406170 439438 406226
rect 439494 406170 439562 406226
rect 439618 406170 439686 406226
rect 439742 406170 439838 406226
rect 439218 406102 439838 406170
rect 439218 406046 439314 406102
rect 439370 406046 439438 406102
rect 439494 406046 439562 406102
rect 439618 406046 439686 406102
rect 439742 406046 439838 406102
rect 439218 405978 439838 406046
rect 439218 405922 439314 405978
rect 439370 405922 439438 405978
rect 439494 405922 439562 405978
rect 439618 405922 439686 405978
rect 439742 405922 439838 405978
rect 439218 388350 439838 405922
rect 439218 388294 439314 388350
rect 439370 388294 439438 388350
rect 439494 388294 439562 388350
rect 439618 388294 439686 388350
rect 439742 388294 439838 388350
rect 439218 388226 439838 388294
rect 439218 388170 439314 388226
rect 439370 388170 439438 388226
rect 439494 388170 439562 388226
rect 439618 388170 439686 388226
rect 439742 388170 439838 388226
rect 439218 388102 439838 388170
rect 439218 388046 439314 388102
rect 439370 388046 439438 388102
rect 439494 388046 439562 388102
rect 439618 388046 439686 388102
rect 439742 388046 439838 388102
rect 439218 387978 439838 388046
rect 439218 387922 439314 387978
rect 439370 387922 439438 387978
rect 439494 387922 439562 387978
rect 439618 387922 439686 387978
rect 439742 387922 439838 387978
rect 439218 370350 439838 387922
rect 466218 400350 466838 408578
rect 466218 400294 466314 400350
rect 466370 400294 466438 400350
rect 466494 400294 466562 400350
rect 466618 400294 466686 400350
rect 466742 400294 466838 400350
rect 466218 400226 466838 400294
rect 466218 400170 466314 400226
rect 466370 400170 466438 400226
rect 466494 400170 466562 400226
rect 466618 400170 466686 400226
rect 466742 400170 466838 400226
rect 466218 400102 466838 400170
rect 466218 400046 466314 400102
rect 466370 400046 466438 400102
rect 466494 400046 466562 400102
rect 466618 400046 466686 400102
rect 466742 400046 466838 400102
rect 466218 399978 466838 400046
rect 466218 399922 466314 399978
rect 466370 399922 466438 399978
rect 466494 399922 466562 399978
rect 466618 399922 466686 399978
rect 466742 399922 466838 399978
rect 439218 370294 439314 370350
rect 439370 370294 439438 370350
rect 439494 370294 439562 370350
rect 439618 370294 439686 370350
rect 439742 370294 439838 370350
rect 439218 370226 439838 370294
rect 439218 370170 439314 370226
rect 439370 370170 439438 370226
rect 439494 370170 439562 370226
rect 439618 370170 439686 370226
rect 439742 370170 439838 370226
rect 439218 370102 439838 370170
rect 439218 370046 439314 370102
rect 439370 370046 439438 370102
rect 439494 370046 439562 370102
rect 439618 370046 439686 370102
rect 439742 370046 439838 370102
rect 439218 369978 439838 370046
rect 439218 369922 439314 369978
rect 439370 369922 439438 369978
rect 439494 369922 439562 369978
rect 439618 369922 439686 369978
rect 439742 369922 439838 369978
rect 439218 352350 439838 369922
rect 439218 352294 439314 352350
rect 439370 352294 439438 352350
rect 439494 352294 439562 352350
rect 439618 352294 439686 352350
rect 439742 352294 439838 352350
rect 439218 352226 439838 352294
rect 439218 352170 439314 352226
rect 439370 352170 439438 352226
rect 439494 352170 439562 352226
rect 439618 352170 439686 352226
rect 439742 352170 439838 352226
rect 439218 352102 439838 352170
rect 439218 352046 439314 352102
rect 439370 352046 439438 352102
rect 439494 352046 439562 352102
rect 439618 352046 439686 352102
rect 439742 352046 439838 352102
rect 439218 351978 439838 352046
rect 439218 351922 439314 351978
rect 439370 351922 439438 351978
rect 439494 351922 439562 351978
rect 439618 351922 439686 351978
rect 439742 351922 439838 351978
rect 439218 334350 439838 351922
rect 439218 334294 439314 334350
rect 439370 334294 439438 334350
rect 439494 334294 439562 334350
rect 439618 334294 439686 334350
rect 439742 334294 439838 334350
rect 439218 334226 439838 334294
rect 439218 334170 439314 334226
rect 439370 334170 439438 334226
rect 439494 334170 439562 334226
rect 439618 334170 439686 334226
rect 439742 334170 439838 334226
rect 439218 334102 439838 334170
rect 439218 334046 439314 334102
rect 439370 334046 439438 334102
rect 439494 334046 439562 334102
rect 439618 334046 439686 334102
rect 439742 334046 439838 334102
rect 439218 333978 439838 334046
rect 439218 333922 439314 333978
rect 439370 333922 439438 333978
rect 439494 333922 439562 333978
rect 439618 333922 439686 333978
rect 439742 333922 439838 333978
rect 435498 310294 435594 310350
rect 435650 310294 435718 310350
rect 435774 310294 435842 310350
rect 435898 310294 435966 310350
rect 436022 310294 436118 310350
rect 435498 310226 436118 310294
rect 435498 310170 435594 310226
rect 435650 310170 435718 310226
rect 435774 310170 435842 310226
rect 435898 310170 435966 310226
rect 436022 310170 436118 310226
rect 435498 310102 436118 310170
rect 435498 310046 435594 310102
rect 435650 310046 435718 310102
rect 435774 310046 435842 310102
rect 435898 310046 435966 310102
rect 436022 310046 436118 310102
rect 435498 309978 436118 310046
rect 435498 309922 435594 309978
rect 435650 309922 435718 309978
rect 435774 309922 435842 309978
rect 435898 309922 435966 309978
rect 436022 309922 436118 309978
rect 435498 292350 436118 309922
rect 435498 292294 435594 292350
rect 435650 292294 435718 292350
rect 435774 292294 435842 292350
rect 435898 292294 435966 292350
rect 436022 292294 436118 292350
rect 435498 292226 436118 292294
rect 435498 292170 435594 292226
rect 435650 292170 435718 292226
rect 435774 292170 435842 292226
rect 435898 292170 435966 292226
rect 436022 292170 436118 292226
rect 435498 292102 436118 292170
rect 435498 292046 435594 292102
rect 435650 292046 435718 292102
rect 435774 292046 435842 292102
rect 435898 292046 435966 292102
rect 436022 292046 436118 292102
rect 435498 291978 436118 292046
rect 435498 291922 435594 291978
rect 435650 291922 435718 291978
rect 435774 291922 435842 291978
rect 435898 291922 435966 291978
rect 436022 291922 436118 291978
rect 435498 274350 436118 291922
rect 435498 274294 435594 274350
rect 435650 274294 435718 274350
rect 435774 274294 435842 274350
rect 435898 274294 435966 274350
rect 436022 274294 436118 274350
rect 435498 274226 436118 274294
rect 435498 274170 435594 274226
rect 435650 274170 435718 274226
rect 435774 274170 435842 274226
rect 435898 274170 435966 274226
rect 436022 274170 436118 274226
rect 435498 274102 436118 274170
rect 435498 274046 435594 274102
rect 435650 274046 435718 274102
rect 435774 274046 435842 274102
rect 435898 274046 435966 274102
rect 436022 274046 436118 274102
rect 435498 273978 436118 274046
rect 435498 273922 435594 273978
rect 435650 273922 435718 273978
rect 435774 273922 435842 273978
rect 435898 273922 435966 273978
rect 436022 273922 436118 273978
rect 435498 256350 436118 273922
rect 435498 256294 435594 256350
rect 435650 256294 435718 256350
rect 435774 256294 435842 256350
rect 435898 256294 435966 256350
rect 436022 256294 436118 256350
rect 435498 256226 436118 256294
rect 435498 256170 435594 256226
rect 435650 256170 435718 256226
rect 435774 256170 435842 256226
rect 435898 256170 435966 256226
rect 436022 256170 436118 256226
rect 435498 256102 436118 256170
rect 435498 256046 435594 256102
rect 435650 256046 435718 256102
rect 435774 256046 435842 256102
rect 435898 256046 435966 256102
rect 436022 256046 436118 256102
rect 435498 255978 436118 256046
rect 435498 255922 435594 255978
rect 435650 255922 435718 255978
rect 435774 255922 435842 255978
rect 435898 255922 435966 255978
rect 436022 255922 436118 255978
rect 435498 238350 436118 255922
rect 435498 238294 435594 238350
rect 435650 238294 435718 238350
rect 435774 238294 435842 238350
rect 435898 238294 435966 238350
rect 436022 238294 436118 238350
rect 435498 238226 436118 238294
rect 435498 238170 435594 238226
rect 435650 238170 435718 238226
rect 435774 238170 435842 238226
rect 435898 238170 435966 238226
rect 436022 238170 436118 238226
rect 435498 238102 436118 238170
rect 435498 238046 435594 238102
rect 435650 238046 435718 238102
rect 435774 238046 435842 238102
rect 435898 238046 435966 238102
rect 436022 238046 436118 238102
rect 435498 237978 436118 238046
rect 435498 237922 435594 237978
rect 435650 237922 435718 237978
rect 435774 237922 435842 237978
rect 435898 237922 435966 237978
rect 436022 237922 436118 237978
rect 435498 220350 436118 237922
rect 435498 220294 435594 220350
rect 435650 220294 435718 220350
rect 435774 220294 435842 220350
rect 435898 220294 435966 220350
rect 436022 220294 436118 220350
rect 435498 220226 436118 220294
rect 435498 220170 435594 220226
rect 435650 220170 435718 220226
rect 435774 220170 435842 220226
rect 435898 220170 435966 220226
rect 436022 220170 436118 220226
rect 435498 220102 436118 220170
rect 435498 220046 435594 220102
rect 435650 220046 435718 220102
rect 435774 220046 435842 220102
rect 435898 220046 435966 220102
rect 436022 220046 436118 220102
rect 435498 219978 436118 220046
rect 435498 219922 435594 219978
rect 435650 219922 435718 219978
rect 435774 219922 435842 219978
rect 435898 219922 435966 219978
rect 436022 219922 436118 219978
rect 435498 202350 436118 219922
rect 435498 202294 435594 202350
rect 435650 202294 435718 202350
rect 435774 202294 435842 202350
rect 435898 202294 435966 202350
rect 436022 202294 436118 202350
rect 435498 202226 436118 202294
rect 435498 202170 435594 202226
rect 435650 202170 435718 202226
rect 435774 202170 435842 202226
rect 435898 202170 435966 202226
rect 436022 202170 436118 202226
rect 435498 202102 436118 202170
rect 435498 202046 435594 202102
rect 435650 202046 435718 202102
rect 435774 202046 435842 202102
rect 435898 202046 435966 202102
rect 436022 202046 436118 202102
rect 435498 201978 436118 202046
rect 435498 201922 435594 201978
rect 435650 201922 435718 201978
rect 435774 201922 435842 201978
rect 435898 201922 435966 201978
rect 436022 201922 436118 201978
rect 435498 184350 436118 201922
rect 435498 184294 435594 184350
rect 435650 184294 435718 184350
rect 435774 184294 435842 184350
rect 435898 184294 435966 184350
rect 436022 184294 436118 184350
rect 435498 184226 436118 184294
rect 435498 184170 435594 184226
rect 435650 184170 435718 184226
rect 435774 184170 435842 184226
rect 435898 184170 435966 184226
rect 436022 184170 436118 184226
rect 435498 184102 436118 184170
rect 435498 184046 435594 184102
rect 435650 184046 435718 184102
rect 435774 184046 435842 184102
rect 435898 184046 435966 184102
rect 436022 184046 436118 184102
rect 435498 183978 436118 184046
rect 435498 183922 435594 183978
rect 435650 183922 435718 183978
rect 435774 183922 435842 183978
rect 435898 183922 435966 183978
rect 436022 183922 436118 183978
rect 435498 166350 436118 183922
rect 435498 166294 435594 166350
rect 435650 166294 435718 166350
rect 435774 166294 435842 166350
rect 435898 166294 435966 166350
rect 436022 166294 436118 166350
rect 435498 166226 436118 166294
rect 435498 166170 435594 166226
rect 435650 166170 435718 166226
rect 435774 166170 435842 166226
rect 435898 166170 435966 166226
rect 436022 166170 436118 166226
rect 435498 166102 436118 166170
rect 435498 166046 435594 166102
rect 435650 166046 435718 166102
rect 435774 166046 435842 166102
rect 435898 166046 435966 166102
rect 436022 166046 436118 166102
rect 435498 165978 436118 166046
rect 435498 165922 435594 165978
rect 435650 165922 435718 165978
rect 435774 165922 435842 165978
rect 435898 165922 435966 165978
rect 436022 165922 436118 165978
rect 435498 148350 436118 165922
rect 435498 148294 435594 148350
rect 435650 148294 435718 148350
rect 435774 148294 435842 148350
rect 435898 148294 435966 148350
rect 436022 148294 436118 148350
rect 435498 148226 436118 148294
rect 435498 148170 435594 148226
rect 435650 148170 435718 148226
rect 435774 148170 435842 148226
rect 435898 148170 435966 148226
rect 436022 148170 436118 148226
rect 435498 148102 436118 148170
rect 435498 148046 435594 148102
rect 435650 148046 435718 148102
rect 435774 148046 435842 148102
rect 435898 148046 435966 148102
rect 436022 148046 436118 148102
rect 435498 147978 436118 148046
rect 435498 147922 435594 147978
rect 435650 147922 435718 147978
rect 435774 147922 435842 147978
rect 435898 147922 435966 147978
rect 436022 147922 436118 147978
rect 435498 130350 436118 147922
rect 435498 130294 435594 130350
rect 435650 130294 435718 130350
rect 435774 130294 435842 130350
rect 435898 130294 435966 130350
rect 436022 130294 436118 130350
rect 435498 130226 436118 130294
rect 435498 130170 435594 130226
rect 435650 130170 435718 130226
rect 435774 130170 435842 130226
rect 435898 130170 435966 130226
rect 436022 130170 436118 130226
rect 435498 130102 436118 130170
rect 435498 130046 435594 130102
rect 435650 130046 435718 130102
rect 435774 130046 435842 130102
rect 435898 130046 435966 130102
rect 436022 130046 436118 130102
rect 435498 129978 436118 130046
rect 435498 129922 435594 129978
rect 435650 129922 435718 129978
rect 435774 129922 435842 129978
rect 435898 129922 435966 129978
rect 436022 129922 436118 129978
rect 435498 112350 436118 129922
rect 437612 320068 437668 320078
rect 437612 113092 437668 320012
rect 437612 113026 437668 113036
rect 439218 316350 439838 333922
rect 464492 384418 464548 384428
rect 451052 327572 451108 327582
rect 439218 316294 439314 316350
rect 439370 316294 439438 316350
rect 439494 316294 439562 316350
rect 439618 316294 439686 316350
rect 439742 316294 439838 316350
rect 439218 316226 439838 316294
rect 439218 316170 439314 316226
rect 439370 316170 439438 316226
rect 439494 316170 439562 316226
rect 439618 316170 439686 316226
rect 439742 316170 439838 316226
rect 439218 316102 439838 316170
rect 439218 316046 439314 316102
rect 439370 316046 439438 316102
rect 439494 316046 439562 316102
rect 439618 316046 439686 316102
rect 439742 316046 439838 316102
rect 439218 315978 439838 316046
rect 439218 315922 439314 315978
rect 439370 315922 439438 315978
rect 439494 315922 439562 315978
rect 439618 315922 439686 315978
rect 439742 315922 439838 315978
rect 439218 298350 439838 315922
rect 439218 298294 439314 298350
rect 439370 298294 439438 298350
rect 439494 298294 439562 298350
rect 439618 298294 439686 298350
rect 439742 298294 439838 298350
rect 439218 298226 439838 298294
rect 439218 298170 439314 298226
rect 439370 298170 439438 298226
rect 439494 298170 439562 298226
rect 439618 298170 439686 298226
rect 439742 298170 439838 298226
rect 439218 298102 439838 298170
rect 439218 298046 439314 298102
rect 439370 298046 439438 298102
rect 439494 298046 439562 298102
rect 439618 298046 439686 298102
rect 439742 298046 439838 298102
rect 439218 297978 439838 298046
rect 439218 297922 439314 297978
rect 439370 297922 439438 297978
rect 439494 297922 439562 297978
rect 439618 297922 439686 297978
rect 439742 297922 439838 297978
rect 439218 280350 439838 297922
rect 439218 280294 439314 280350
rect 439370 280294 439438 280350
rect 439494 280294 439562 280350
rect 439618 280294 439686 280350
rect 439742 280294 439838 280350
rect 439218 280226 439838 280294
rect 439218 280170 439314 280226
rect 439370 280170 439438 280226
rect 439494 280170 439562 280226
rect 439618 280170 439686 280226
rect 439742 280170 439838 280226
rect 439218 280102 439838 280170
rect 439218 280046 439314 280102
rect 439370 280046 439438 280102
rect 439494 280046 439562 280102
rect 439618 280046 439686 280102
rect 439742 280046 439838 280102
rect 439218 279978 439838 280046
rect 439218 279922 439314 279978
rect 439370 279922 439438 279978
rect 439494 279922 439562 279978
rect 439618 279922 439686 279978
rect 439742 279922 439838 279978
rect 439218 262350 439838 279922
rect 442652 321972 442708 321982
rect 439218 262294 439314 262350
rect 439370 262294 439438 262350
rect 439494 262294 439562 262350
rect 439618 262294 439686 262350
rect 439742 262294 439838 262350
rect 439218 262226 439838 262294
rect 439218 262170 439314 262226
rect 439370 262170 439438 262226
rect 439494 262170 439562 262226
rect 439618 262170 439686 262226
rect 439742 262170 439838 262226
rect 439218 262102 439838 262170
rect 439218 262046 439314 262102
rect 439370 262046 439438 262102
rect 439494 262046 439562 262102
rect 439618 262046 439686 262102
rect 439742 262046 439838 262102
rect 439218 261978 439838 262046
rect 439218 261922 439314 261978
rect 439370 261922 439438 261978
rect 439494 261922 439562 261978
rect 439618 261922 439686 261978
rect 439742 261922 439838 261978
rect 439218 244350 439838 261922
rect 439218 244294 439314 244350
rect 439370 244294 439438 244350
rect 439494 244294 439562 244350
rect 439618 244294 439686 244350
rect 439742 244294 439838 244350
rect 439218 244226 439838 244294
rect 439218 244170 439314 244226
rect 439370 244170 439438 244226
rect 439494 244170 439562 244226
rect 439618 244170 439686 244226
rect 439742 244170 439838 244226
rect 439218 244102 439838 244170
rect 439218 244046 439314 244102
rect 439370 244046 439438 244102
rect 439494 244046 439562 244102
rect 439618 244046 439686 244102
rect 439742 244046 439838 244102
rect 439218 243978 439838 244046
rect 439218 243922 439314 243978
rect 439370 243922 439438 243978
rect 439494 243922 439562 243978
rect 439618 243922 439686 243978
rect 439742 243922 439838 243978
rect 439218 226350 439838 243922
rect 439218 226294 439314 226350
rect 439370 226294 439438 226350
rect 439494 226294 439562 226350
rect 439618 226294 439686 226350
rect 439742 226294 439838 226350
rect 439218 226226 439838 226294
rect 439218 226170 439314 226226
rect 439370 226170 439438 226226
rect 439494 226170 439562 226226
rect 439618 226170 439686 226226
rect 439742 226170 439838 226226
rect 439218 226102 439838 226170
rect 439218 226046 439314 226102
rect 439370 226046 439438 226102
rect 439494 226046 439562 226102
rect 439618 226046 439686 226102
rect 439742 226046 439838 226102
rect 439218 225978 439838 226046
rect 439218 225922 439314 225978
rect 439370 225922 439438 225978
rect 439494 225922 439562 225978
rect 439618 225922 439686 225978
rect 439742 225922 439838 225978
rect 439218 208350 439838 225922
rect 439218 208294 439314 208350
rect 439370 208294 439438 208350
rect 439494 208294 439562 208350
rect 439618 208294 439686 208350
rect 439742 208294 439838 208350
rect 439218 208226 439838 208294
rect 439218 208170 439314 208226
rect 439370 208170 439438 208226
rect 439494 208170 439562 208226
rect 439618 208170 439686 208226
rect 439742 208170 439838 208226
rect 439218 208102 439838 208170
rect 439218 208046 439314 208102
rect 439370 208046 439438 208102
rect 439494 208046 439562 208102
rect 439618 208046 439686 208102
rect 439742 208046 439838 208102
rect 439218 207978 439838 208046
rect 439218 207922 439314 207978
rect 439370 207922 439438 207978
rect 439494 207922 439562 207978
rect 439618 207922 439686 207978
rect 439742 207922 439838 207978
rect 439218 190350 439838 207922
rect 439218 190294 439314 190350
rect 439370 190294 439438 190350
rect 439494 190294 439562 190350
rect 439618 190294 439686 190350
rect 439742 190294 439838 190350
rect 439218 190226 439838 190294
rect 439218 190170 439314 190226
rect 439370 190170 439438 190226
rect 439494 190170 439562 190226
rect 439618 190170 439686 190226
rect 439742 190170 439838 190226
rect 439218 190102 439838 190170
rect 439218 190046 439314 190102
rect 439370 190046 439438 190102
rect 439494 190046 439562 190102
rect 439618 190046 439686 190102
rect 439742 190046 439838 190102
rect 439218 189978 439838 190046
rect 439218 189922 439314 189978
rect 439370 189922 439438 189978
rect 439494 189922 439562 189978
rect 439618 189922 439686 189978
rect 439742 189922 439838 189978
rect 439218 172350 439838 189922
rect 439218 172294 439314 172350
rect 439370 172294 439438 172350
rect 439494 172294 439562 172350
rect 439618 172294 439686 172350
rect 439742 172294 439838 172350
rect 439218 172226 439838 172294
rect 439218 172170 439314 172226
rect 439370 172170 439438 172226
rect 439494 172170 439562 172226
rect 439618 172170 439686 172226
rect 439742 172170 439838 172226
rect 439218 172102 439838 172170
rect 439218 172046 439314 172102
rect 439370 172046 439438 172102
rect 439494 172046 439562 172102
rect 439618 172046 439686 172102
rect 439742 172046 439838 172102
rect 439218 171978 439838 172046
rect 439218 171922 439314 171978
rect 439370 171922 439438 171978
rect 439494 171922 439562 171978
rect 439618 171922 439686 171978
rect 439742 171922 439838 171978
rect 439218 154350 439838 171922
rect 439218 154294 439314 154350
rect 439370 154294 439438 154350
rect 439494 154294 439562 154350
rect 439618 154294 439686 154350
rect 439742 154294 439838 154350
rect 439218 154226 439838 154294
rect 439218 154170 439314 154226
rect 439370 154170 439438 154226
rect 439494 154170 439562 154226
rect 439618 154170 439686 154226
rect 439742 154170 439838 154226
rect 439218 154102 439838 154170
rect 439218 154046 439314 154102
rect 439370 154046 439438 154102
rect 439494 154046 439562 154102
rect 439618 154046 439686 154102
rect 439742 154046 439838 154102
rect 439218 153978 439838 154046
rect 439218 153922 439314 153978
rect 439370 153922 439438 153978
rect 439494 153922 439562 153978
rect 439618 153922 439686 153978
rect 439742 153922 439838 153978
rect 439218 136350 439838 153922
rect 439218 136294 439314 136350
rect 439370 136294 439438 136350
rect 439494 136294 439562 136350
rect 439618 136294 439686 136350
rect 439742 136294 439838 136350
rect 439218 136226 439838 136294
rect 439218 136170 439314 136226
rect 439370 136170 439438 136226
rect 439494 136170 439562 136226
rect 439618 136170 439686 136226
rect 439742 136170 439838 136226
rect 439218 136102 439838 136170
rect 439218 136046 439314 136102
rect 439370 136046 439438 136102
rect 439494 136046 439562 136102
rect 439618 136046 439686 136102
rect 439742 136046 439838 136102
rect 439218 135978 439838 136046
rect 439218 135922 439314 135978
rect 439370 135922 439438 135978
rect 439494 135922 439562 135978
rect 439618 135922 439686 135978
rect 439742 135922 439838 135978
rect 439218 118350 439838 135922
rect 439218 118294 439314 118350
rect 439370 118294 439438 118350
rect 439494 118294 439562 118350
rect 439618 118294 439686 118350
rect 439742 118294 439838 118350
rect 439218 118226 439838 118294
rect 439218 118170 439314 118226
rect 439370 118170 439438 118226
rect 439494 118170 439562 118226
rect 439618 118170 439686 118226
rect 439742 118170 439838 118226
rect 439218 118102 439838 118170
rect 439218 118046 439314 118102
rect 439370 118046 439438 118102
rect 439494 118046 439562 118102
rect 439618 118046 439686 118102
rect 439742 118046 439838 118102
rect 439218 117978 439838 118046
rect 439218 117922 439314 117978
rect 439370 117922 439438 117978
rect 439494 117922 439562 117978
rect 439618 117922 439686 117978
rect 439742 117922 439838 117978
rect 435498 112294 435594 112350
rect 435650 112294 435718 112350
rect 435774 112294 435842 112350
rect 435898 112294 435966 112350
rect 436022 112294 436118 112350
rect 435498 112226 436118 112294
rect 435498 112170 435594 112226
rect 435650 112170 435718 112226
rect 435774 112170 435842 112226
rect 435898 112170 435966 112226
rect 436022 112170 436118 112226
rect 435498 112102 436118 112170
rect 435498 112046 435594 112102
rect 435650 112046 435718 112102
rect 435774 112046 435842 112102
rect 435898 112046 435966 112102
rect 436022 112046 436118 112102
rect 435498 111978 436118 112046
rect 435498 111922 435594 111978
rect 435650 111922 435718 111978
rect 435774 111922 435842 111978
rect 435898 111922 435966 111978
rect 436022 111922 436118 111978
rect 432572 107202 432628 107212
rect 430892 104290 430948 104300
rect 429212 98466 429268 98476
rect 427644 59602 427700 59612
rect 435498 94350 436118 111922
rect 435498 94294 435594 94350
rect 435650 94294 435718 94350
rect 435774 94294 435842 94350
rect 435898 94294 435966 94350
rect 436022 94294 436118 94350
rect 435498 94226 436118 94294
rect 435498 94170 435594 94226
rect 435650 94170 435718 94226
rect 435774 94170 435842 94226
rect 435898 94170 435966 94226
rect 436022 94170 436118 94226
rect 435498 94102 436118 94170
rect 435498 94046 435594 94102
rect 435650 94046 435718 94102
rect 435774 94046 435842 94102
rect 435898 94046 435966 94102
rect 436022 94046 436118 94102
rect 435498 93978 436118 94046
rect 435498 93922 435594 93978
rect 435650 93922 435718 93978
rect 435774 93922 435842 93978
rect 435898 93922 435966 93978
rect 436022 93922 436118 93978
rect 435498 76350 436118 93922
rect 435498 76294 435594 76350
rect 435650 76294 435718 76350
rect 435774 76294 435842 76350
rect 435898 76294 435966 76350
rect 436022 76294 436118 76350
rect 435498 76226 436118 76294
rect 435498 76170 435594 76226
rect 435650 76170 435718 76226
rect 435774 76170 435842 76226
rect 435898 76170 435966 76226
rect 436022 76170 436118 76226
rect 435498 76102 436118 76170
rect 435498 76046 435594 76102
rect 435650 76046 435718 76102
rect 435774 76046 435842 76102
rect 435898 76046 435966 76102
rect 436022 76046 436118 76102
rect 435498 75978 436118 76046
rect 435498 75922 435594 75978
rect 435650 75922 435718 75978
rect 435774 75922 435842 75978
rect 435898 75922 435966 75978
rect 436022 75922 436118 75978
rect 425852 50306 425908 50316
rect 435498 58350 436118 75922
rect 435498 58294 435594 58350
rect 435650 58294 435718 58350
rect 435774 58294 435842 58350
rect 435898 58294 435966 58350
rect 436022 58294 436118 58350
rect 435498 58226 436118 58294
rect 435498 58170 435594 58226
rect 435650 58170 435718 58226
rect 435774 58170 435842 58226
rect 435898 58170 435966 58226
rect 436022 58170 436118 58226
rect 435498 58102 436118 58170
rect 435498 58046 435594 58102
rect 435650 58046 435718 58102
rect 435774 58046 435842 58102
rect 435898 58046 435966 58102
rect 436022 58046 436118 58102
rect 435498 57978 436118 58046
rect 435498 57922 435594 57978
rect 435650 57922 435718 57978
rect 435774 57922 435842 57978
rect 435898 57922 435966 57978
rect 436022 57922 436118 57978
rect 411852 32722 411908 32732
rect 435498 40350 436118 57922
rect 435498 40294 435594 40350
rect 435650 40294 435718 40350
rect 435774 40294 435842 40350
rect 435898 40294 435966 40350
rect 436022 40294 436118 40350
rect 435498 40226 436118 40294
rect 435498 40170 435594 40226
rect 435650 40170 435718 40226
rect 435774 40170 435842 40226
rect 435898 40170 435966 40226
rect 436022 40170 436118 40226
rect 435498 40102 436118 40170
rect 435498 40046 435594 40102
rect 435650 40046 435718 40102
rect 435774 40046 435842 40102
rect 435898 40046 435966 40102
rect 436022 40046 436118 40102
rect 435498 39978 436118 40046
rect 435498 39922 435594 39978
rect 435650 39922 435718 39978
rect 435774 39922 435842 39978
rect 435898 39922 435966 39978
rect 436022 39922 436118 39978
rect 411628 9202 411684 9212
rect 435498 22350 436118 39922
rect 435498 22294 435594 22350
rect 435650 22294 435718 22350
rect 435774 22294 435842 22350
rect 435898 22294 435966 22350
rect 436022 22294 436118 22350
rect 435498 22226 436118 22294
rect 435498 22170 435594 22226
rect 435650 22170 435718 22226
rect 435774 22170 435842 22226
rect 435898 22170 435966 22226
rect 436022 22170 436118 22226
rect 435498 22102 436118 22170
rect 435498 22046 435594 22102
rect 435650 22046 435718 22102
rect 435774 22046 435842 22102
rect 435898 22046 435966 22102
rect 436022 22046 436118 22102
rect 435498 21978 436118 22046
rect 435498 21922 435594 21978
rect 435650 21922 435718 21978
rect 435774 21922 435842 21978
rect 435898 21922 435966 21978
rect 436022 21922 436118 21978
rect 408498 -1176 408594 -1120
rect 408650 -1176 408718 -1120
rect 408774 -1176 408842 -1120
rect 408898 -1176 408966 -1120
rect 409022 -1176 409118 -1120
rect 408498 -1244 409118 -1176
rect 408498 -1300 408594 -1244
rect 408650 -1300 408718 -1244
rect 408774 -1300 408842 -1244
rect 408898 -1300 408966 -1244
rect 409022 -1300 409118 -1244
rect 408498 -1368 409118 -1300
rect 408498 -1424 408594 -1368
rect 408650 -1424 408718 -1368
rect 408774 -1424 408842 -1368
rect 408898 -1424 408966 -1368
rect 409022 -1424 409118 -1368
rect 408498 -1492 409118 -1424
rect 408498 -1548 408594 -1492
rect 408650 -1548 408718 -1492
rect 408774 -1548 408842 -1492
rect 408898 -1548 408966 -1492
rect 409022 -1548 409118 -1492
rect 408498 -1644 409118 -1548
rect 435498 4350 436118 21922
rect 435498 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 436118 4350
rect 435498 4226 436118 4294
rect 435498 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 436118 4226
rect 435498 4102 436118 4170
rect 435498 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 436118 4102
rect 435498 3978 436118 4046
rect 435498 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 436118 3978
rect 435498 -160 436118 3922
rect 435498 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 436118 -160
rect 435498 -284 436118 -216
rect 435498 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 436118 -284
rect 435498 -408 436118 -340
rect 435498 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 436118 -408
rect 435498 -532 436118 -464
rect 435498 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 436118 -532
rect 435498 -1644 436118 -588
rect 439218 100350 439838 117922
rect 439218 100294 439314 100350
rect 439370 100294 439438 100350
rect 439494 100294 439562 100350
rect 439618 100294 439686 100350
rect 439742 100294 439838 100350
rect 439218 100226 439838 100294
rect 439218 100170 439314 100226
rect 439370 100170 439438 100226
rect 439494 100170 439562 100226
rect 439618 100170 439686 100226
rect 439742 100170 439838 100226
rect 439218 100102 439838 100170
rect 439218 100046 439314 100102
rect 439370 100046 439438 100102
rect 439494 100046 439562 100102
rect 439618 100046 439686 100102
rect 439742 100046 439838 100102
rect 439218 99978 439838 100046
rect 439218 99922 439314 99978
rect 439370 99922 439438 99978
rect 439494 99922 439562 99978
rect 439618 99922 439686 99978
rect 439742 99922 439838 99978
rect 439218 82350 439838 99922
rect 439218 82294 439314 82350
rect 439370 82294 439438 82350
rect 439494 82294 439562 82350
rect 439618 82294 439686 82350
rect 439742 82294 439838 82350
rect 439218 82226 439838 82294
rect 439218 82170 439314 82226
rect 439370 82170 439438 82226
rect 439494 82170 439562 82226
rect 439618 82170 439686 82226
rect 439742 82170 439838 82226
rect 439218 82102 439838 82170
rect 439218 82046 439314 82102
rect 439370 82046 439438 82102
rect 439494 82046 439562 82102
rect 439618 82046 439686 82102
rect 439742 82046 439838 82102
rect 439218 81978 439838 82046
rect 439218 81922 439314 81978
rect 439370 81922 439438 81978
rect 439494 81922 439562 81978
rect 439618 81922 439686 81978
rect 439742 81922 439838 81978
rect 439218 64350 439838 81922
rect 440972 273924 441028 273934
rect 440972 75236 441028 273868
rect 440972 75170 441028 75180
rect 441084 116116 441140 116126
rect 439218 64294 439314 64350
rect 439370 64294 439438 64350
rect 439494 64294 439562 64350
rect 439618 64294 439686 64350
rect 439742 64294 439838 64350
rect 439218 64226 439838 64294
rect 439218 64170 439314 64226
rect 439370 64170 439438 64226
rect 439494 64170 439562 64226
rect 439618 64170 439686 64226
rect 439742 64170 439838 64226
rect 439218 64102 439838 64170
rect 439218 64046 439314 64102
rect 439370 64046 439438 64102
rect 439494 64046 439562 64102
rect 439618 64046 439686 64102
rect 439742 64046 439838 64102
rect 439218 63978 439838 64046
rect 439218 63922 439314 63978
rect 439370 63922 439438 63978
rect 439494 63922 439562 63978
rect 439618 63922 439686 63978
rect 439742 63922 439838 63978
rect 439218 46350 439838 63922
rect 441084 60676 441140 116060
rect 442652 115892 442708 321916
rect 447692 270564 447748 270574
rect 446012 268884 446068 268894
rect 442652 115826 442708 115836
rect 444332 267204 444388 267214
rect 444332 66500 444388 267148
rect 446012 69412 446068 268828
rect 447692 72212 447748 270508
rect 447692 72146 447748 72156
rect 449372 265524 449428 265534
rect 446012 69346 446068 69356
rect 444332 66434 444388 66444
rect 449372 63588 449428 265468
rect 451052 130564 451108 327516
rect 456092 323092 456148 323102
rect 454412 313348 454468 313358
rect 451052 130498 451108 130508
rect 452732 275604 452788 275614
rect 452732 78148 452788 275548
rect 454412 95620 454468 313292
rect 456092 118916 456148 323036
rect 457772 214228 457828 214238
rect 456988 152068 457044 152078
rect 456988 148596 457044 152012
rect 456988 148530 457044 148540
rect 456092 118850 456148 118860
rect 454412 95554 454468 95564
rect 452732 78082 452788 78092
rect 449372 63522 449428 63532
rect 441084 60610 441140 60620
rect 457660 59668 457716 59678
rect 457660 57764 457716 59612
rect 457660 57698 457716 57708
rect 457772 54852 457828 214172
rect 464492 198118 464548 384362
rect 464492 198052 464548 198062
rect 466218 382350 466838 399922
rect 466218 382294 466314 382350
rect 466370 382294 466438 382350
rect 466494 382294 466562 382350
rect 466618 382294 466686 382350
rect 466742 382294 466838 382350
rect 466218 382226 466838 382294
rect 466218 382170 466314 382226
rect 466370 382170 466438 382226
rect 466494 382170 466562 382226
rect 466618 382170 466686 382226
rect 466742 382170 466838 382226
rect 466218 382102 466838 382170
rect 466218 382046 466314 382102
rect 466370 382046 466438 382102
rect 466494 382046 466562 382102
rect 466618 382046 466686 382102
rect 466742 382046 466838 382102
rect 466218 381978 466838 382046
rect 466218 381922 466314 381978
rect 466370 381922 466438 381978
rect 466494 381922 466562 381978
rect 466618 381922 466686 381978
rect 466742 381922 466838 381978
rect 466218 364350 466838 381922
rect 466218 364294 466314 364350
rect 466370 364294 466438 364350
rect 466494 364294 466562 364350
rect 466618 364294 466686 364350
rect 466742 364294 466838 364350
rect 466218 364226 466838 364294
rect 466218 364170 466314 364226
rect 466370 364170 466438 364226
rect 466494 364170 466562 364226
rect 466618 364170 466686 364226
rect 466742 364170 466838 364226
rect 466218 364102 466838 364170
rect 466218 364046 466314 364102
rect 466370 364046 466438 364102
rect 466494 364046 466562 364102
rect 466618 364046 466686 364102
rect 466742 364046 466838 364102
rect 466218 363978 466838 364046
rect 466218 363922 466314 363978
rect 466370 363922 466438 363978
rect 466494 363922 466562 363978
rect 466618 363922 466686 363978
rect 466742 363922 466838 363978
rect 466218 346350 466838 363922
rect 466218 346294 466314 346350
rect 466370 346294 466438 346350
rect 466494 346294 466562 346350
rect 466618 346294 466686 346350
rect 466742 346294 466838 346350
rect 466218 346226 466838 346294
rect 466218 346170 466314 346226
rect 466370 346170 466438 346226
rect 466494 346170 466562 346226
rect 466618 346170 466686 346226
rect 466742 346170 466838 346226
rect 466218 346102 466838 346170
rect 466218 346046 466314 346102
rect 466370 346046 466438 346102
rect 466494 346046 466562 346102
rect 466618 346046 466686 346102
rect 466742 346046 466838 346102
rect 466218 345978 466838 346046
rect 466218 345922 466314 345978
rect 466370 345922 466438 345978
rect 466494 345922 466562 345978
rect 466618 345922 466686 345978
rect 466742 345922 466838 345978
rect 466218 328350 466838 345922
rect 466218 328294 466314 328350
rect 466370 328294 466438 328350
rect 466494 328294 466562 328350
rect 466618 328294 466686 328350
rect 466742 328294 466838 328350
rect 466218 328226 466838 328294
rect 466218 328170 466314 328226
rect 466370 328170 466438 328226
rect 466494 328170 466562 328226
rect 466618 328170 466686 328226
rect 466742 328170 466838 328226
rect 466218 328102 466838 328170
rect 466218 328046 466314 328102
rect 466370 328046 466438 328102
rect 466494 328046 466562 328102
rect 466618 328046 466686 328102
rect 466742 328046 466838 328102
rect 466218 327978 466838 328046
rect 466218 327922 466314 327978
rect 466370 327922 466438 327978
rect 466494 327922 466562 327978
rect 466618 327922 466686 327978
rect 466742 327922 466838 327978
rect 466218 310350 466838 327922
rect 466218 310294 466314 310350
rect 466370 310294 466438 310350
rect 466494 310294 466562 310350
rect 466618 310294 466686 310350
rect 466742 310294 466838 310350
rect 466218 310226 466838 310294
rect 466218 310170 466314 310226
rect 466370 310170 466438 310226
rect 466494 310170 466562 310226
rect 466618 310170 466686 310226
rect 466742 310170 466838 310226
rect 466218 310102 466838 310170
rect 466218 310046 466314 310102
rect 466370 310046 466438 310102
rect 466494 310046 466562 310102
rect 466618 310046 466686 310102
rect 466742 310046 466838 310102
rect 466218 309978 466838 310046
rect 466218 309922 466314 309978
rect 466370 309922 466438 309978
rect 466494 309922 466562 309978
rect 466618 309922 466686 309978
rect 466742 309922 466838 309978
rect 466218 292350 466838 309922
rect 466218 292294 466314 292350
rect 466370 292294 466438 292350
rect 466494 292294 466562 292350
rect 466618 292294 466686 292350
rect 466742 292294 466838 292350
rect 466218 292226 466838 292294
rect 466218 292170 466314 292226
rect 466370 292170 466438 292226
rect 466494 292170 466562 292226
rect 466618 292170 466686 292226
rect 466742 292170 466838 292226
rect 466218 292102 466838 292170
rect 466218 292046 466314 292102
rect 466370 292046 466438 292102
rect 466494 292046 466562 292102
rect 466618 292046 466686 292102
rect 466742 292046 466838 292102
rect 466218 291978 466838 292046
rect 466218 291922 466314 291978
rect 466370 291922 466438 291978
rect 466494 291922 466562 291978
rect 466618 291922 466686 291978
rect 466742 291922 466838 291978
rect 466218 274350 466838 291922
rect 466218 274294 466314 274350
rect 466370 274294 466438 274350
rect 466494 274294 466562 274350
rect 466618 274294 466686 274350
rect 466742 274294 466838 274350
rect 466218 274226 466838 274294
rect 466218 274170 466314 274226
rect 466370 274170 466438 274226
rect 466494 274170 466562 274226
rect 466618 274170 466686 274226
rect 466742 274170 466838 274226
rect 466218 274102 466838 274170
rect 466218 274046 466314 274102
rect 466370 274046 466438 274102
rect 466494 274046 466562 274102
rect 466618 274046 466686 274102
rect 466742 274046 466838 274102
rect 466218 273978 466838 274046
rect 466218 273922 466314 273978
rect 466370 273922 466438 273978
rect 466494 273922 466562 273978
rect 466618 273922 466686 273978
rect 466742 273922 466838 273978
rect 466218 256350 466838 273922
rect 466218 256294 466314 256350
rect 466370 256294 466438 256350
rect 466494 256294 466562 256350
rect 466618 256294 466686 256350
rect 466742 256294 466838 256350
rect 466218 256226 466838 256294
rect 466218 256170 466314 256226
rect 466370 256170 466438 256226
rect 466494 256170 466562 256226
rect 466618 256170 466686 256226
rect 466742 256170 466838 256226
rect 466218 256102 466838 256170
rect 466218 256046 466314 256102
rect 466370 256046 466438 256102
rect 466494 256046 466562 256102
rect 466618 256046 466686 256102
rect 466742 256046 466838 256102
rect 466218 255978 466838 256046
rect 466218 255922 466314 255978
rect 466370 255922 466438 255978
rect 466494 255922 466562 255978
rect 466618 255922 466686 255978
rect 466742 255922 466838 255978
rect 466218 238350 466838 255922
rect 466218 238294 466314 238350
rect 466370 238294 466438 238350
rect 466494 238294 466562 238350
rect 466618 238294 466686 238350
rect 466742 238294 466838 238350
rect 466218 238226 466838 238294
rect 466218 238170 466314 238226
rect 466370 238170 466438 238226
rect 466494 238170 466562 238226
rect 466618 238170 466686 238226
rect 466742 238170 466838 238226
rect 466218 238102 466838 238170
rect 466218 238046 466314 238102
rect 466370 238046 466438 238102
rect 466494 238046 466562 238102
rect 466618 238046 466686 238102
rect 466742 238046 466838 238102
rect 466218 237978 466838 238046
rect 466218 237922 466314 237978
rect 466370 237922 466438 237978
rect 466494 237922 466562 237978
rect 466618 237922 466686 237978
rect 466742 237922 466838 237978
rect 466218 220350 466838 237922
rect 466218 220294 466314 220350
rect 466370 220294 466438 220350
rect 466494 220294 466562 220350
rect 466618 220294 466686 220350
rect 466742 220294 466838 220350
rect 466218 220226 466838 220294
rect 466218 220170 466314 220226
rect 466370 220170 466438 220226
rect 466494 220170 466562 220226
rect 466618 220170 466686 220226
rect 466742 220170 466838 220226
rect 466218 220102 466838 220170
rect 466218 220046 466314 220102
rect 466370 220046 466438 220102
rect 466494 220046 466562 220102
rect 466618 220046 466686 220102
rect 466742 220046 466838 220102
rect 466218 219978 466838 220046
rect 466218 219922 466314 219978
rect 466370 219922 466438 219978
rect 466494 219922 466562 219978
rect 466618 219922 466686 219978
rect 466742 219922 466838 219978
rect 466218 202350 466838 219922
rect 466218 202294 466314 202350
rect 466370 202294 466438 202350
rect 466494 202294 466562 202350
rect 466618 202294 466686 202350
rect 466742 202294 466838 202350
rect 466218 202226 466838 202294
rect 466218 202170 466314 202226
rect 466370 202170 466438 202226
rect 466494 202170 466562 202226
rect 466618 202170 466686 202226
rect 466742 202170 466838 202226
rect 466218 202102 466838 202170
rect 466218 202046 466314 202102
rect 466370 202046 466438 202102
rect 466494 202046 466562 202102
rect 466618 202046 466686 202102
rect 466742 202046 466838 202102
rect 466218 201978 466838 202046
rect 466218 201922 466314 201978
rect 466370 201922 466438 201978
rect 466494 201922 466562 201978
rect 466618 201922 466686 201978
rect 466742 201922 466838 201978
rect 466218 184350 466838 201922
rect 466218 184294 466314 184350
rect 466370 184294 466438 184350
rect 466494 184294 466562 184350
rect 466618 184294 466686 184350
rect 466742 184294 466838 184350
rect 466218 184226 466838 184294
rect 466218 184170 466314 184226
rect 466370 184170 466438 184226
rect 466494 184170 466562 184226
rect 466618 184170 466686 184226
rect 466742 184170 466838 184226
rect 466218 184102 466838 184170
rect 466218 184046 466314 184102
rect 466370 184046 466438 184102
rect 466494 184046 466562 184102
rect 466618 184046 466686 184102
rect 466742 184046 466838 184102
rect 466218 183978 466838 184046
rect 466218 183922 466314 183978
rect 466370 183922 466438 183978
rect 466494 183922 466562 183978
rect 466618 183922 466686 183978
rect 466742 183922 466838 183978
rect 466218 166350 466838 183922
rect 466218 166294 466314 166350
rect 466370 166294 466438 166350
rect 466494 166294 466562 166350
rect 466618 166294 466686 166350
rect 466742 166294 466838 166350
rect 466218 166226 466838 166294
rect 466218 166170 466314 166226
rect 466370 166170 466438 166226
rect 466494 166170 466562 166226
rect 466618 166170 466686 166226
rect 466742 166170 466838 166226
rect 466218 166102 466838 166170
rect 466218 166046 466314 166102
rect 466370 166046 466438 166102
rect 466494 166046 466562 166102
rect 466618 166046 466686 166102
rect 466742 166046 466838 166102
rect 466218 165978 466838 166046
rect 466218 165922 466314 165978
rect 466370 165922 466438 165978
rect 466494 165922 466562 165978
rect 466618 165922 466686 165978
rect 466742 165922 466838 165978
rect 466218 149870 466838 165922
rect 469938 406350 470558 408578
rect 477148 407764 477204 407774
rect 475468 407652 475524 407662
rect 475468 407458 475524 407596
rect 477148 407638 477204 407708
rect 477148 407572 477204 407582
rect 475468 407392 475524 407402
rect 469938 406294 470034 406350
rect 470090 406294 470158 406350
rect 470214 406294 470282 406350
rect 470338 406294 470406 406350
rect 470462 406294 470558 406350
rect 469938 406226 470558 406294
rect 469938 406170 470034 406226
rect 470090 406170 470158 406226
rect 470214 406170 470282 406226
rect 470338 406170 470406 406226
rect 470462 406170 470558 406226
rect 469938 406102 470558 406170
rect 469938 406046 470034 406102
rect 470090 406046 470158 406102
rect 470214 406046 470282 406102
rect 470338 406046 470406 406102
rect 470462 406046 470558 406102
rect 469938 405978 470558 406046
rect 469938 405922 470034 405978
rect 470090 405922 470158 405978
rect 470214 405922 470282 405978
rect 470338 405922 470406 405978
rect 470462 405922 470558 405978
rect 469938 388350 470558 405922
rect 469938 388294 470034 388350
rect 470090 388294 470158 388350
rect 470214 388294 470282 388350
rect 470338 388294 470406 388350
rect 470462 388294 470558 388350
rect 469938 388226 470558 388294
rect 469938 388170 470034 388226
rect 470090 388170 470158 388226
rect 470214 388170 470282 388226
rect 470338 388170 470406 388226
rect 470462 388170 470558 388226
rect 469938 388102 470558 388170
rect 469938 388046 470034 388102
rect 470090 388046 470158 388102
rect 470214 388046 470282 388102
rect 470338 388046 470406 388102
rect 470462 388046 470558 388102
rect 469938 387978 470558 388046
rect 469938 387922 470034 387978
rect 470090 387922 470158 387978
rect 470214 387922 470282 387978
rect 470338 387922 470406 387978
rect 470462 387922 470558 387978
rect 469938 370350 470558 387922
rect 496938 400350 497558 408578
rect 496938 400294 497034 400350
rect 497090 400294 497158 400350
rect 497214 400294 497282 400350
rect 497338 400294 497406 400350
rect 497462 400294 497558 400350
rect 496938 400226 497558 400294
rect 496938 400170 497034 400226
rect 497090 400170 497158 400226
rect 497214 400170 497282 400226
rect 497338 400170 497406 400226
rect 497462 400170 497558 400226
rect 496938 400102 497558 400170
rect 496938 400046 497034 400102
rect 497090 400046 497158 400102
rect 497214 400046 497282 400102
rect 497338 400046 497406 400102
rect 497462 400046 497558 400102
rect 496938 399978 497558 400046
rect 496938 399922 497034 399978
rect 497090 399922 497158 399978
rect 497214 399922 497282 399978
rect 497338 399922 497406 399978
rect 497462 399922 497558 399978
rect 469938 370294 470034 370350
rect 470090 370294 470158 370350
rect 470214 370294 470282 370350
rect 470338 370294 470406 370350
rect 470462 370294 470558 370350
rect 469938 370226 470558 370294
rect 469938 370170 470034 370226
rect 470090 370170 470158 370226
rect 470214 370170 470282 370226
rect 470338 370170 470406 370226
rect 470462 370170 470558 370226
rect 469938 370102 470558 370170
rect 469938 370046 470034 370102
rect 470090 370046 470158 370102
rect 470214 370046 470282 370102
rect 470338 370046 470406 370102
rect 470462 370046 470558 370102
rect 469938 369978 470558 370046
rect 469938 369922 470034 369978
rect 470090 369922 470158 369978
rect 470214 369922 470282 369978
rect 470338 369922 470406 369978
rect 470462 369922 470558 369978
rect 469938 352350 470558 369922
rect 469938 352294 470034 352350
rect 470090 352294 470158 352350
rect 470214 352294 470282 352350
rect 470338 352294 470406 352350
rect 470462 352294 470558 352350
rect 469938 352226 470558 352294
rect 469938 352170 470034 352226
rect 470090 352170 470158 352226
rect 470214 352170 470282 352226
rect 470338 352170 470406 352226
rect 470462 352170 470558 352226
rect 469938 352102 470558 352170
rect 469938 352046 470034 352102
rect 470090 352046 470158 352102
rect 470214 352046 470282 352102
rect 470338 352046 470406 352102
rect 470462 352046 470558 352102
rect 469938 351978 470558 352046
rect 469938 351922 470034 351978
rect 470090 351922 470158 351978
rect 470214 351922 470282 351978
rect 470338 351922 470406 351978
rect 470462 351922 470558 351978
rect 469938 334350 470558 351922
rect 469938 334294 470034 334350
rect 470090 334294 470158 334350
rect 470214 334294 470282 334350
rect 470338 334294 470406 334350
rect 470462 334294 470558 334350
rect 469938 334226 470558 334294
rect 469938 334170 470034 334226
rect 470090 334170 470158 334226
rect 470214 334170 470282 334226
rect 470338 334170 470406 334226
rect 470462 334170 470558 334226
rect 469938 334102 470558 334170
rect 469938 334046 470034 334102
rect 470090 334046 470158 334102
rect 470214 334046 470282 334102
rect 470338 334046 470406 334102
rect 470462 334046 470558 334102
rect 469938 333978 470558 334046
rect 469938 333922 470034 333978
rect 470090 333922 470158 333978
rect 470214 333922 470282 333978
rect 470338 333922 470406 333978
rect 470462 333922 470558 333978
rect 469938 316350 470558 333922
rect 469938 316294 470034 316350
rect 470090 316294 470158 316350
rect 470214 316294 470282 316350
rect 470338 316294 470406 316350
rect 470462 316294 470558 316350
rect 469938 316226 470558 316294
rect 469938 316170 470034 316226
rect 470090 316170 470158 316226
rect 470214 316170 470282 316226
rect 470338 316170 470406 316226
rect 470462 316170 470558 316226
rect 469938 316102 470558 316170
rect 469938 316046 470034 316102
rect 470090 316046 470158 316102
rect 470214 316046 470282 316102
rect 470338 316046 470406 316102
rect 470462 316046 470558 316102
rect 469938 315978 470558 316046
rect 469938 315922 470034 315978
rect 470090 315922 470158 315978
rect 470214 315922 470282 315978
rect 470338 315922 470406 315978
rect 470462 315922 470558 315978
rect 469938 298350 470558 315922
rect 469938 298294 470034 298350
rect 470090 298294 470158 298350
rect 470214 298294 470282 298350
rect 470338 298294 470406 298350
rect 470462 298294 470558 298350
rect 469938 298226 470558 298294
rect 469938 298170 470034 298226
rect 470090 298170 470158 298226
rect 470214 298170 470282 298226
rect 470338 298170 470406 298226
rect 470462 298170 470558 298226
rect 469938 298102 470558 298170
rect 469938 298046 470034 298102
rect 470090 298046 470158 298102
rect 470214 298046 470282 298102
rect 470338 298046 470406 298102
rect 470462 298046 470558 298102
rect 469938 297978 470558 298046
rect 469938 297922 470034 297978
rect 470090 297922 470158 297978
rect 470214 297922 470282 297978
rect 470338 297922 470406 297978
rect 470462 297922 470558 297978
rect 469938 280350 470558 297922
rect 469938 280294 470034 280350
rect 470090 280294 470158 280350
rect 470214 280294 470282 280350
rect 470338 280294 470406 280350
rect 470462 280294 470558 280350
rect 469938 280226 470558 280294
rect 469938 280170 470034 280226
rect 470090 280170 470158 280226
rect 470214 280170 470282 280226
rect 470338 280170 470406 280226
rect 470462 280170 470558 280226
rect 469938 280102 470558 280170
rect 469938 280046 470034 280102
rect 470090 280046 470158 280102
rect 470214 280046 470282 280102
rect 470338 280046 470406 280102
rect 470462 280046 470558 280102
rect 469938 279978 470558 280046
rect 469938 279922 470034 279978
rect 470090 279922 470158 279978
rect 470214 279922 470282 279978
rect 470338 279922 470406 279978
rect 470462 279922 470558 279978
rect 469938 262350 470558 279922
rect 469938 262294 470034 262350
rect 470090 262294 470158 262350
rect 470214 262294 470282 262350
rect 470338 262294 470406 262350
rect 470462 262294 470558 262350
rect 469938 262226 470558 262294
rect 469938 262170 470034 262226
rect 470090 262170 470158 262226
rect 470214 262170 470282 262226
rect 470338 262170 470406 262226
rect 470462 262170 470558 262226
rect 469938 262102 470558 262170
rect 469938 262046 470034 262102
rect 470090 262046 470158 262102
rect 470214 262046 470282 262102
rect 470338 262046 470406 262102
rect 470462 262046 470558 262102
rect 469938 261978 470558 262046
rect 469938 261922 470034 261978
rect 470090 261922 470158 261978
rect 470214 261922 470282 261978
rect 470338 261922 470406 261978
rect 470462 261922 470558 261978
rect 469938 244350 470558 261922
rect 469938 244294 470034 244350
rect 470090 244294 470158 244350
rect 470214 244294 470282 244350
rect 470338 244294 470406 244350
rect 470462 244294 470558 244350
rect 469938 244226 470558 244294
rect 469938 244170 470034 244226
rect 470090 244170 470158 244226
rect 470214 244170 470282 244226
rect 470338 244170 470406 244226
rect 470462 244170 470558 244226
rect 469938 244102 470558 244170
rect 469938 244046 470034 244102
rect 470090 244046 470158 244102
rect 470214 244046 470282 244102
rect 470338 244046 470406 244102
rect 470462 244046 470558 244102
rect 469938 243978 470558 244046
rect 469938 243922 470034 243978
rect 470090 243922 470158 243978
rect 470214 243922 470282 243978
rect 470338 243922 470406 243978
rect 470462 243922 470558 243978
rect 469938 226350 470558 243922
rect 469938 226294 470034 226350
rect 470090 226294 470158 226350
rect 470214 226294 470282 226350
rect 470338 226294 470406 226350
rect 470462 226294 470558 226350
rect 469938 226226 470558 226294
rect 469938 226170 470034 226226
rect 470090 226170 470158 226226
rect 470214 226170 470282 226226
rect 470338 226170 470406 226226
rect 470462 226170 470558 226226
rect 469938 226102 470558 226170
rect 469938 226046 470034 226102
rect 470090 226046 470158 226102
rect 470214 226046 470282 226102
rect 470338 226046 470406 226102
rect 470462 226046 470558 226102
rect 469938 225978 470558 226046
rect 469938 225922 470034 225978
rect 470090 225922 470158 225978
rect 470214 225922 470282 225978
rect 470338 225922 470406 225978
rect 470462 225922 470558 225978
rect 469938 208350 470558 225922
rect 469938 208294 470034 208350
rect 470090 208294 470158 208350
rect 470214 208294 470282 208350
rect 470338 208294 470406 208350
rect 470462 208294 470558 208350
rect 469938 208226 470558 208294
rect 469938 208170 470034 208226
rect 470090 208170 470158 208226
rect 470214 208170 470282 208226
rect 470338 208170 470406 208226
rect 470462 208170 470558 208226
rect 469938 208102 470558 208170
rect 469938 208046 470034 208102
rect 470090 208046 470158 208102
rect 470214 208046 470282 208102
rect 470338 208046 470406 208102
rect 470462 208046 470558 208102
rect 469938 207978 470558 208046
rect 469938 207922 470034 207978
rect 470090 207922 470158 207978
rect 470214 207922 470282 207978
rect 470338 207922 470406 207978
rect 470462 207922 470558 207978
rect 469938 190350 470558 207922
rect 476252 384238 476308 384248
rect 476252 197938 476308 384182
rect 476252 197872 476308 197882
rect 479612 384058 479668 384068
rect 479612 197758 479668 384002
rect 481292 383878 481348 383888
rect 481292 198100 481348 383822
rect 496938 382350 497558 399922
rect 496938 382294 497034 382350
rect 497090 382294 497158 382350
rect 497214 382294 497282 382350
rect 497338 382294 497406 382350
rect 497462 382294 497558 382350
rect 496938 382226 497558 382294
rect 496938 382170 497034 382226
rect 497090 382170 497158 382226
rect 497214 382170 497282 382226
rect 497338 382170 497406 382226
rect 497462 382170 497558 382226
rect 496938 382102 497558 382170
rect 496938 382046 497034 382102
rect 497090 382046 497158 382102
rect 497214 382046 497282 382102
rect 497338 382046 497406 382102
rect 497462 382046 497558 382102
rect 496938 381978 497558 382046
rect 496938 381922 497034 381978
rect 497090 381922 497158 381978
rect 497214 381922 497282 381978
rect 497338 381922 497406 381978
rect 497462 381922 497558 381978
rect 496938 364350 497558 381922
rect 496938 364294 497034 364350
rect 497090 364294 497158 364350
rect 497214 364294 497282 364350
rect 497338 364294 497406 364350
rect 497462 364294 497558 364350
rect 496938 364226 497558 364294
rect 496938 364170 497034 364226
rect 497090 364170 497158 364226
rect 497214 364170 497282 364226
rect 497338 364170 497406 364226
rect 497462 364170 497558 364226
rect 496938 364102 497558 364170
rect 496938 364046 497034 364102
rect 497090 364046 497158 364102
rect 497214 364046 497282 364102
rect 497338 364046 497406 364102
rect 497462 364046 497558 364102
rect 496938 363978 497558 364046
rect 496938 363922 497034 363978
rect 497090 363922 497158 363978
rect 497214 363922 497282 363978
rect 497338 363922 497406 363978
rect 497462 363922 497558 363978
rect 496938 346350 497558 363922
rect 496938 346294 497034 346350
rect 497090 346294 497158 346350
rect 497214 346294 497282 346350
rect 497338 346294 497406 346350
rect 497462 346294 497558 346350
rect 496938 346226 497558 346294
rect 496938 346170 497034 346226
rect 497090 346170 497158 346226
rect 497214 346170 497282 346226
rect 497338 346170 497406 346226
rect 497462 346170 497558 346226
rect 496938 346102 497558 346170
rect 496938 346046 497034 346102
rect 497090 346046 497158 346102
rect 497214 346046 497282 346102
rect 497338 346046 497406 346102
rect 497462 346046 497558 346102
rect 496938 345978 497558 346046
rect 496938 345922 497034 345978
rect 497090 345922 497158 345978
rect 497214 345922 497282 345978
rect 497338 345922 497406 345978
rect 497462 345922 497558 345978
rect 496938 328350 497558 345922
rect 496938 328294 497034 328350
rect 497090 328294 497158 328350
rect 497214 328294 497282 328350
rect 497338 328294 497406 328350
rect 497462 328294 497558 328350
rect 496938 328226 497558 328294
rect 496938 328170 497034 328226
rect 497090 328170 497158 328226
rect 497214 328170 497282 328226
rect 497338 328170 497406 328226
rect 497462 328170 497558 328226
rect 496938 328102 497558 328170
rect 496938 328046 497034 328102
rect 497090 328046 497158 328102
rect 497214 328046 497282 328102
rect 497338 328046 497406 328102
rect 497462 328046 497558 328102
rect 496938 327978 497558 328046
rect 496938 327922 497034 327978
rect 497090 327922 497158 327978
rect 497214 327922 497282 327978
rect 497338 327922 497406 327978
rect 497462 327922 497558 327978
rect 496938 310350 497558 327922
rect 496938 310294 497034 310350
rect 497090 310294 497158 310350
rect 497214 310294 497282 310350
rect 497338 310294 497406 310350
rect 497462 310294 497558 310350
rect 496938 310226 497558 310294
rect 496938 310170 497034 310226
rect 497090 310170 497158 310226
rect 497214 310170 497282 310226
rect 497338 310170 497406 310226
rect 497462 310170 497558 310226
rect 496938 310102 497558 310170
rect 496938 310046 497034 310102
rect 497090 310046 497158 310102
rect 497214 310046 497282 310102
rect 497338 310046 497406 310102
rect 497462 310046 497558 310102
rect 496938 309978 497558 310046
rect 496938 309922 497034 309978
rect 497090 309922 497158 309978
rect 497214 309922 497282 309978
rect 497338 309922 497406 309978
rect 497462 309922 497558 309978
rect 496938 292350 497558 309922
rect 496938 292294 497034 292350
rect 497090 292294 497158 292350
rect 497214 292294 497282 292350
rect 497338 292294 497406 292350
rect 497462 292294 497558 292350
rect 496938 292226 497558 292294
rect 496938 292170 497034 292226
rect 497090 292170 497158 292226
rect 497214 292170 497282 292226
rect 497338 292170 497406 292226
rect 497462 292170 497558 292226
rect 496938 292102 497558 292170
rect 496938 292046 497034 292102
rect 497090 292046 497158 292102
rect 497214 292046 497282 292102
rect 497338 292046 497406 292102
rect 497462 292046 497558 292102
rect 496938 291978 497558 292046
rect 496938 291922 497034 291978
rect 497090 291922 497158 291978
rect 497214 291922 497282 291978
rect 497338 291922 497406 291978
rect 497462 291922 497558 291978
rect 496938 274350 497558 291922
rect 496938 274294 497034 274350
rect 497090 274294 497158 274350
rect 497214 274294 497282 274350
rect 497338 274294 497406 274350
rect 497462 274294 497558 274350
rect 496938 274226 497558 274294
rect 496938 274170 497034 274226
rect 497090 274170 497158 274226
rect 497214 274170 497282 274226
rect 497338 274170 497406 274226
rect 497462 274170 497558 274226
rect 496938 274102 497558 274170
rect 496938 274046 497034 274102
rect 497090 274046 497158 274102
rect 497214 274046 497282 274102
rect 497338 274046 497406 274102
rect 497462 274046 497558 274102
rect 496938 273978 497558 274046
rect 496938 273922 497034 273978
rect 497090 273922 497158 273978
rect 497214 273922 497282 273978
rect 497338 273922 497406 273978
rect 497462 273922 497558 273978
rect 496938 256350 497558 273922
rect 496938 256294 497034 256350
rect 497090 256294 497158 256350
rect 497214 256294 497282 256350
rect 497338 256294 497406 256350
rect 497462 256294 497558 256350
rect 496938 256226 497558 256294
rect 496938 256170 497034 256226
rect 497090 256170 497158 256226
rect 497214 256170 497282 256226
rect 497338 256170 497406 256226
rect 497462 256170 497558 256226
rect 496938 256102 497558 256170
rect 496938 256046 497034 256102
rect 497090 256046 497158 256102
rect 497214 256046 497282 256102
rect 497338 256046 497406 256102
rect 497462 256046 497558 256102
rect 496938 255978 497558 256046
rect 496938 255922 497034 255978
rect 497090 255922 497158 255978
rect 497214 255922 497282 255978
rect 497338 255922 497406 255978
rect 497462 255922 497558 255978
rect 496938 238350 497558 255922
rect 496938 238294 497034 238350
rect 497090 238294 497158 238350
rect 497214 238294 497282 238350
rect 497338 238294 497406 238350
rect 497462 238294 497558 238350
rect 496938 238226 497558 238294
rect 496938 238170 497034 238226
rect 497090 238170 497158 238226
rect 497214 238170 497282 238226
rect 497338 238170 497406 238226
rect 497462 238170 497558 238226
rect 496938 238102 497558 238170
rect 496938 238046 497034 238102
rect 497090 238046 497158 238102
rect 497214 238046 497282 238102
rect 497338 238046 497406 238102
rect 497462 238046 497558 238102
rect 496938 237978 497558 238046
rect 496938 237922 497034 237978
rect 497090 237922 497158 237978
rect 497214 237922 497282 237978
rect 497338 237922 497406 237978
rect 497462 237922 497558 237978
rect 496938 233230 497558 237922
rect 500658 406350 501278 408578
rect 500658 406294 500754 406350
rect 500810 406294 500878 406350
rect 500934 406294 501002 406350
rect 501058 406294 501126 406350
rect 501182 406294 501278 406350
rect 500658 406226 501278 406294
rect 500658 406170 500754 406226
rect 500810 406170 500878 406226
rect 500934 406170 501002 406226
rect 501058 406170 501126 406226
rect 501182 406170 501278 406226
rect 500658 406102 501278 406170
rect 500658 406046 500754 406102
rect 500810 406046 500878 406102
rect 500934 406046 501002 406102
rect 501058 406046 501126 406102
rect 501182 406046 501278 406102
rect 500658 405978 501278 406046
rect 500658 405922 500754 405978
rect 500810 405922 500878 405978
rect 500934 405922 501002 405978
rect 501058 405922 501126 405978
rect 501182 405922 501278 405978
rect 500658 388350 501278 405922
rect 500658 388294 500754 388350
rect 500810 388294 500878 388350
rect 500934 388294 501002 388350
rect 501058 388294 501126 388350
rect 501182 388294 501278 388350
rect 500658 388226 501278 388294
rect 500658 388170 500754 388226
rect 500810 388170 500878 388226
rect 500934 388170 501002 388226
rect 501058 388170 501126 388226
rect 501182 388170 501278 388226
rect 500658 388102 501278 388170
rect 500658 388046 500754 388102
rect 500810 388046 500878 388102
rect 500934 388046 501002 388102
rect 501058 388046 501126 388102
rect 501182 388046 501278 388102
rect 500658 387978 501278 388046
rect 500658 387922 500754 387978
rect 500810 387922 500878 387978
rect 500934 387922 501002 387978
rect 501058 387922 501126 387978
rect 501182 387922 501278 387978
rect 500658 370350 501278 387922
rect 527658 400350 528278 408578
rect 527658 400294 527754 400350
rect 527810 400294 527878 400350
rect 527934 400294 528002 400350
rect 528058 400294 528126 400350
rect 528182 400294 528278 400350
rect 527658 400226 528278 400294
rect 527658 400170 527754 400226
rect 527810 400170 527878 400226
rect 527934 400170 528002 400226
rect 528058 400170 528126 400226
rect 528182 400170 528278 400226
rect 527658 400102 528278 400170
rect 527658 400046 527754 400102
rect 527810 400046 527878 400102
rect 527934 400046 528002 400102
rect 528058 400046 528126 400102
rect 528182 400046 528278 400102
rect 527658 399978 528278 400046
rect 527658 399922 527754 399978
rect 527810 399922 527878 399978
rect 527934 399922 528002 399978
rect 528058 399922 528126 399978
rect 528182 399922 528278 399978
rect 500658 370294 500754 370350
rect 500810 370294 500878 370350
rect 500934 370294 501002 370350
rect 501058 370294 501126 370350
rect 501182 370294 501278 370350
rect 500658 370226 501278 370294
rect 500658 370170 500754 370226
rect 500810 370170 500878 370226
rect 500934 370170 501002 370226
rect 501058 370170 501126 370226
rect 501182 370170 501278 370226
rect 500658 370102 501278 370170
rect 500658 370046 500754 370102
rect 500810 370046 500878 370102
rect 500934 370046 501002 370102
rect 501058 370046 501126 370102
rect 501182 370046 501278 370102
rect 500658 369978 501278 370046
rect 500658 369922 500754 369978
rect 500810 369922 500878 369978
rect 500934 369922 501002 369978
rect 501058 369922 501126 369978
rect 501182 369922 501278 369978
rect 500658 352350 501278 369922
rect 500658 352294 500754 352350
rect 500810 352294 500878 352350
rect 500934 352294 501002 352350
rect 501058 352294 501126 352350
rect 501182 352294 501278 352350
rect 500658 352226 501278 352294
rect 500658 352170 500754 352226
rect 500810 352170 500878 352226
rect 500934 352170 501002 352226
rect 501058 352170 501126 352226
rect 501182 352170 501278 352226
rect 500658 352102 501278 352170
rect 500658 352046 500754 352102
rect 500810 352046 500878 352102
rect 500934 352046 501002 352102
rect 501058 352046 501126 352102
rect 501182 352046 501278 352102
rect 500658 351978 501278 352046
rect 500658 351922 500754 351978
rect 500810 351922 500878 351978
rect 500934 351922 501002 351978
rect 501058 351922 501126 351978
rect 501182 351922 501278 351978
rect 500658 334350 501278 351922
rect 519932 382618 519988 382628
rect 519932 349468 519988 382562
rect 527658 382350 528278 399922
rect 527658 382294 527754 382350
rect 527810 382294 527878 382350
rect 527934 382294 528002 382350
rect 528058 382294 528126 382350
rect 528182 382294 528278 382350
rect 527658 382226 528278 382294
rect 527658 382170 527754 382226
rect 527810 382170 527878 382226
rect 527934 382170 528002 382226
rect 528058 382170 528126 382226
rect 528182 382170 528278 382226
rect 527658 382102 528278 382170
rect 527658 382046 527754 382102
rect 527810 382046 527878 382102
rect 527934 382046 528002 382102
rect 528058 382046 528126 382102
rect 528182 382046 528278 382102
rect 527658 381978 528278 382046
rect 527658 381922 527754 381978
rect 527810 381922 527878 381978
rect 527934 381922 528002 381978
rect 528058 381922 528126 381978
rect 528182 381922 528278 381978
rect 527658 364350 528278 381922
rect 527658 364294 527754 364350
rect 527810 364294 527878 364350
rect 527934 364294 528002 364350
rect 528058 364294 528126 364350
rect 528182 364294 528278 364350
rect 527658 364226 528278 364294
rect 527658 364170 527754 364226
rect 527810 364170 527878 364226
rect 527934 364170 528002 364226
rect 528058 364170 528126 364226
rect 528182 364170 528278 364226
rect 527658 364102 528278 364170
rect 527658 364046 527754 364102
rect 527810 364046 527878 364102
rect 527934 364046 528002 364102
rect 528058 364046 528126 364102
rect 528182 364046 528278 364102
rect 527658 363978 528278 364046
rect 527658 363922 527754 363978
rect 527810 363922 527878 363978
rect 527934 363922 528002 363978
rect 528058 363922 528126 363978
rect 528182 363922 528278 363978
rect 519932 349412 520100 349468
rect 500658 334294 500754 334350
rect 500810 334294 500878 334350
rect 500934 334294 501002 334350
rect 501058 334294 501126 334350
rect 501182 334294 501278 334350
rect 500658 334226 501278 334294
rect 500658 334170 500754 334226
rect 500810 334170 500878 334226
rect 500934 334170 501002 334226
rect 501058 334170 501126 334226
rect 501182 334170 501278 334226
rect 500658 334102 501278 334170
rect 500658 334046 500754 334102
rect 500810 334046 500878 334102
rect 500934 334046 501002 334102
rect 501058 334046 501126 334102
rect 501182 334046 501278 334102
rect 500658 333978 501278 334046
rect 500658 333922 500754 333978
rect 500810 333922 500878 333978
rect 500934 333922 501002 333978
rect 501058 333922 501126 333978
rect 501182 333922 501278 333978
rect 500658 316350 501278 333922
rect 520044 324324 520100 349412
rect 520044 324258 520100 324268
rect 527658 346350 528278 363922
rect 527658 346294 527754 346350
rect 527810 346294 527878 346350
rect 527934 346294 528002 346350
rect 528058 346294 528126 346350
rect 528182 346294 528278 346350
rect 527658 346226 528278 346294
rect 527658 346170 527754 346226
rect 527810 346170 527878 346226
rect 527934 346170 528002 346226
rect 528058 346170 528126 346226
rect 528182 346170 528278 346226
rect 527658 346102 528278 346170
rect 527658 346046 527754 346102
rect 527810 346046 527878 346102
rect 527934 346046 528002 346102
rect 528058 346046 528126 346102
rect 528182 346046 528278 346102
rect 527658 345978 528278 346046
rect 527658 345922 527754 345978
rect 527810 345922 527878 345978
rect 527934 345922 528002 345978
rect 528058 345922 528126 345978
rect 528182 345922 528278 345978
rect 527658 328350 528278 345922
rect 527658 328294 527754 328350
rect 527810 328294 527878 328350
rect 527934 328294 528002 328350
rect 528058 328294 528126 328350
rect 528182 328294 528278 328350
rect 527658 328226 528278 328294
rect 527658 328170 527754 328226
rect 527810 328170 527878 328226
rect 527934 328170 528002 328226
rect 528058 328170 528126 328226
rect 528182 328170 528278 328226
rect 527658 328102 528278 328170
rect 527658 328046 527754 328102
rect 527810 328046 527878 328102
rect 527934 328046 528002 328102
rect 528058 328046 528126 328102
rect 528182 328046 528278 328102
rect 527658 327978 528278 328046
rect 527658 327922 527754 327978
rect 527810 327922 527878 327978
rect 527934 327922 528002 327978
rect 528058 327922 528126 327978
rect 528182 327922 528278 327978
rect 500658 316294 500754 316350
rect 500810 316294 500878 316350
rect 500934 316294 501002 316350
rect 501058 316294 501126 316350
rect 501182 316294 501278 316350
rect 500658 316226 501278 316294
rect 500658 316170 500754 316226
rect 500810 316170 500878 316226
rect 500934 316170 501002 316226
rect 501058 316170 501126 316226
rect 501182 316170 501278 316226
rect 500658 316102 501278 316170
rect 500658 316046 500754 316102
rect 500810 316046 500878 316102
rect 500934 316046 501002 316102
rect 501058 316046 501126 316102
rect 501182 316046 501278 316102
rect 500658 315978 501278 316046
rect 500658 315922 500754 315978
rect 500810 315922 500878 315978
rect 500934 315922 501002 315978
rect 501058 315922 501126 315978
rect 501182 315922 501278 315978
rect 500658 298350 501278 315922
rect 500658 298294 500754 298350
rect 500810 298294 500878 298350
rect 500934 298294 501002 298350
rect 501058 298294 501126 298350
rect 501182 298294 501278 298350
rect 500658 298226 501278 298294
rect 500658 298170 500754 298226
rect 500810 298170 500878 298226
rect 500934 298170 501002 298226
rect 501058 298170 501126 298226
rect 501182 298170 501278 298226
rect 500658 298102 501278 298170
rect 500658 298046 500754 298102
rect 500810 298046 500878 298102
rect 500934 298046 501002 298102
rect 501058 298046 501126 298102
rect 501182 298046 501278 298102
rect 500658 297978 501278 298046
rect 500658 297922 500754 297978
rect 500810 297922 500878 297978
rect 500934 297922 501002 297978
rect 501058 297922 501126 297978
rect 501182 297922 501278 297978
rect 500658 280350 501278 297922
rect 500658 280294 500754 280350
rect 500810 280294 500878 280350
rect 500934 280294 501002 280350
rect 501058 280294 501126 280350
rect 501182 280294 501278 280350
rect 500658 280226 501278 280294
rect 500658 280170 500754 280226
rect 500810 280170 500878 280226
rect 500934 280170 501002 280226
rect 501058 280170 501126 280226
rect 501182 280170 501278 280226
rect 500658 280102 501278 280170
rect 500658 280046 500754 280102
rect 500810 280046 500878 280102
rect 500934 280046 501002 280102
rect 501058 280046 501126 280102
rect 501182 280046 501278 280102
rect 500658 279978 501278 280046
rect 500658 279922 500754 279978
rect 500810 279922 500878 279978
rect 500934 279922 501002 279978
rect 501058 279922 501126 279978
rect 501182 279922 501278 279978
rect 500658 262350 501278 279922
rect 500658 262294 500754 262350
rect 500810 262294 500878 262350
rect 500934 262294 501002 262350
rect 501058 262294 501126 262350
rect 501182 262294 501278 262350
rect 500658 262226 501278 262294
rect 500658 262170 500754 262226
rect 500810 262170 500878 262226
rect 500934 262170 501002 262226
rect 501058 262170 501126 262226
rect 501182 262170 501278 262226
rect 500658 262102 501278 262170
rect 500658 262046 500754 262102
rect 500810 262046 500878 262102
rect 500934 262046 501002 262102
rect 501058 262046 501126 262102
rect 501182 262046 501278 262102
rect 500658 261978 501278 262046
rect 500658 261922 500754 261978
rect 500810 261922 500878 261978
rect 500934 261922 501002 261978
rect 501058 261922 501126 261978
rect 501182 261922 501278 261978
rect 500658 244350 501278 261922
rect 500658 244294 500754 244350
rect 500810 244294 500878 244350
rect 500934 244294 501002 244350
rect 501058 244294 501126 244350
rect 501182 244294 501278 244350
rect 500658 244226 501278 244294
rect 500658 244170 500754 244226
rect 500810 244170 500878 244226
rect 500934 244170 501002 244226
rect 501058 244170 501126 244226
rect 501182 244170 501278 244226
rect 500658 244102 501278 244170
rect 500658 244046 500754 244102
rect 500810 244046 500878 244102
rect 500934 244046 501002 244102
rect 501058 244046 501126 244102
rect 501182 244046 501278 244102
rect 500658 243978 501278 244046
rect 500658 243922 500754 243978
rect 500810 243922 500878 243978
rect 500934 243922 501002 243978
rect 501058 243922 501126 243978
rect 501182 243922 501278 243978
rect 500658 233230 501278 243922
rect 527658 310350 528278 327922
rect 527658 310294 527754 310350
rect 527810 310294 527878 310350
rect 527934 310294 528002 310350
rect 528058 310294 528126 310350
rect 528182 310294 528278 310350
rect 527658 310226 528278 310294
rect 527658 310170 527754 310226
rect 527810 310170 527878 310226
rect 527934 310170 528002 310226
rect 528058 310170 528126 310226
rect 528182 310170 528278 310226
rect 527658 310102 528278 310170
rect 527658 310046 527754 310102
rect 527810 310046 527878 310102
rect 527934 310046 528002 310102
rect 528058 310046 528126 310102
rect 528182 310046 528278 310102
rect 527658 309978 528278 310046
rect 527658 309922 527754 309978
rect 527810 309922 527878 309978
rect 527934 309922 528002 309978
rect 528058 309922 528126 309978
rect 528182 309922 528278 309978
rect 527658 292350 528278 309922
rect 527658 292294 527754 292350
rect 527810 292294 527878 292350
rect 527934 292294 528002 292350
rect 528058 292294 528126 292350
rect 528182 292294 528278 292350
rect 527658 292226 528278 292294
rect 527658 292170 527754 292226
rect 527810 292170 527878 292226
rect 527934 292170 528002 292226
rect 528058 292170 528126 292226
rect 528182 292170 528278 292226
rect 527658 292102 528278 292170
rect 527658 292046 527754 292102
rect 527810 292046 527878 292102
rect 527934 292046 528002 292102
rect 528058 292046 528126 292102
rect 528182 292046 528278 292102
rect 527658 291978 528278 292046
rect 527658 291922 527754 291978
rect 527810 291922 527878 291978
rect 527934 291922 528002 291978
rect 528058 291922 528126 291978
rect 528182 291922 528278 291978
rect 527658 274350 528278 291922
rect 527658 274294 527754 274350
rect 527810 274294 527878 274350
rect 527934 274294 528002 274350
rect 528058 274294 528126 274350
rect 528182 274294 528278 274350
rect 527658 274226 528278 274294
rect 527658 274170 527754 274226
rect 527810 274170 527878 274226
rect 527934 274170 528002 274226
rect 528058 274170 528126 274226
rect 528182 274170 528278 274226
rect 527658 274102 528278 274170
rect 527658 274046 527754 274102
rect 527810 274046 527878 274102
rect 527934 274046 528002 274102
rect 528058 274046 528126 274102
rect 528182 274046 528278 274102
rect 527658 273978 528278 274046
rect 527658 273922 527754 273978
rect 527810 273922 527878 273978
rect 527934 273922 528002 273978
rect 528058 273922 528126 273978
rect 528182 273922 528278 273978
rect 527658 256350 528278 273922
rect 527658 256294 527754 256350
rect 527810 256294 527878 256350
rect 527934 256294 528002 256350
rect 528058 256294 528126 256350
rect 528182 256294 528278 256350
rect 527658 256226 528278 256294
rect 527658 256170 527754 256226
rect 527810 256170 527878 256226
rect 527934 256170 528002 256226
rect 528058 256170 528126 256226
rect 528182 256170 528278 256226
rect 527658 256102 528278 256170
rect 527658 256046 527754 256102
rect 527810 256046 527878 256102
rect 527934 256046 528002 256102
rect 528058 256046 528126 256102
rect 528182 256046 528278 256102
rect 527658 255978 528278 256046
rect 527658 255922 527754 255978
rect 527810 255922 527878 255978
rect 527934 255922 528002 255978
rect 528058 255922 528126 255978
rect 528182 255922 528278 255978
rect 527658 238350 528278 255922
rect 527658 238294 527754 238350
rect 527810 238294 527878 238350
rect 527934 238294 528002 238350
rect 528058 238294 528126 238350
rect 528182 238294 528278 238350
rect 527658 238226 528278 238294
rect 527658 238170 527754 238226
rect 527810 238170 527878 238226
rect 527934 238170 528002 238226
rect 528058 238170 528126 238226
rect 528182 238170 528278 238226
rect 527658 238102 528278 238170
rect 527658 238046 527754 238102
rect 527810 238046 527878 238102
rect 527934 238046 528002 238102
rect 528058 238046 528126 238102
rect 528182 238046 528278 238102
rect 527658 237978 528278 238046
rect 527658 237922 527754 237978
rect 527810 237922 527878 237978
rect 527934 237922 528002 237978
rect 528058 237922 528126 237978
rect 528182 237922 528278 237978
rect 519148 236740 519204 236750
rect 489752 226350 490072 226384
rect 489752 226294 489822 226350
rect 489878 226294 489946 226350
rect 490002 226294 490072 226350
rect 489752 226226 490072 226294
rect 489752 226170 489822 226226
rect 489878 226170 489946 226226
rect 490002 226170 490072 226226
rect 489752 226102 490072 226170
rect 489752 226046 489822 226102
rect 489878 226046 489946 226102
rect 490002 226046 490072 226102
rect 489752 225978 490072 226046
rect 489752 225922 489822 225978
rect 489878 225922 489946 225978
rect 490002 225922 490072 225978
rect 489752 225888 490072 225922
rect 498320 226350 498640 226384
rect 498320 226294 498390 226350
rect 498446 226294 498514 226350
rect 498570 226294 498640 226350
rect 498320 226226 498640 226294
rect 498320 226170 498390 226226
rect 498446 226170 498514 226226
rect 498570 226170 498640 226226
rect 498320 226102 498640 226170
rect 498320 226046 498390 226102
rect 498446 226046 498514 226102
rect 498570 226046 498640 226102
rect 498320 225978 498640 226046
rect 498320 225922 498390 225978
rect 498446 225922 498514 225978
rect 498570 225922 498640 225978
rect 498320 225888 498640 225922
rect 506888 226350 507208 226384
rect 506888 226294 506958 226350
rect 507014 226294 507082 226350
rect 507138 226294 507208 226350
rect 506888 226226 507208 226294
rect 506888 226170 506958 226226
rect 507014 226170 507082 226226
rect 507138 226170 507208 226226
rect 506888 226102 507208 226170
rect 506888 226046 506958 226102
rect 507014 226046 507082 226102
rect 507138 226046 507208 226102
rect 506888 225978 507208 226046
rect 506888 225922 506958 225978
rect 507014 225922 507082 225978
rect 507138 225922 507208 225978
rect 506888 225888 507208 225922
rect 515456 226350 515776 226384
rect 515456 226294 515526 226350
rect 515582 226294 515650 226350
rect 515706 226294 515776 226350
rect 515456 226226 515776 226294
rect 515456 226170 515526 226226
rect 515582 226170 515650 226226
rect 515706 226170 515776 226226
rect 515456 226102 515776 226170
rect 515456 226046 515526 226102
rect 515582 226046 515650 226102
rect 515706 226046 515776 226102
rect 515456 225978 515776 226046
rect 515456 225922 515526 225978
rect 515582 225922 515650 225978
rect 515706 225922 515776 225978
rect 515456 225888 515776 225922
rect 485468 220350 485788 220384
rect 485468 220294 485538 220350
rect 485594 220294 485662 220350
rect 485718 220294 485788 220350
rect 485468 220226 485788 220294
rect 485468 220170 485538 220226
rect 485594 220170 485662 220226
rect 485718 220170 485788 220226
rect 485468 220102 485788 220170
rect 485468 220046 485538 220102
rect 485594 220046 485662 220102
rect 485718 220046 485788 220102
rect 485468 219978 485788 220046
rect 485468 219922 485538 219978
rect 485594 219922 485662 219978
rect 485718 219922 485788 219978
rect 485468 219888 485788 219922
rect 494036 220350 494356 220384
rect 494036 220294 494106 220350
rect 494162 220294 494230 220350
rect 494286 220294 494356 220350
rect 494036 220226 494356 220294
rect 494036 220170 494106 220226
rect 494162 220170 494230 220226
rect 494286 220170 494356 220226
rect 494036 220102 494356 220170
rect 494036 220046 494106 220102
rect 494162 220046 494230 220102
rect 494286 220046 494356 220102
rect 494036 219978 494356 220046
rect 494036 219922 494106 219978
rect 494162 219922 494230 219978
rect 494286 219922 494356 219978
rect 494036 219888 494356 219922
rect 502604 220350 502924 220384
rect 502604 220294 502674 220350
rect 502730 220294 502798 220350
rect 502854 220294 502924 220350
rect 502604 220226 502924 220294
rect 502604 220170 502674 220226
rect 502730 220170 502798 220226
rect 502854 220170 502924 220226
rect 502604 220102 502924 220170
rect 502604 220046 502674 220102
rect 502730 220046 502798 220102
rect 502854 220046 502924 220102
rect 502604 219978 502924 220046
rect 502604 219922 502674 219978
rect 502730 219922 502798 219978
rect 502854 219922 502924 219978
rect 502604 219888 502924 219922
rect 511172 220350 511492 220384
rect 511172 220294 511242 220350
rect 511298 220294 511366 220350
rect 511422 220294 511492 220350
rect 511172 220226 511492 220294
rect 511172 220170 511242 220226
rect 511298 220170 511366 220226
rect 511422 220170 511492 220226
rect 511172 220102 511492 220170
rect 511172 220046 511242 220102
rect 511298 220046 511366 220102
rect 511422 220046 511492 220102
rect 511172 219978 511492 220046
rect 511172 219922 511242 219978
rect 511298 219922 511366 219978
rect 511422 219922 511492 219978
rect 511172 219888 511492 219922
rect 489752 208350 490072 208384
rect 489752 208294 489822 208350
rect 489878 208294 489946 208350
rect 490002 208294 490072 208350
rect 489752 208226 490072 208294
rect 489752 208170 489822 208226
rect 489878 208170 489946 208226
rect 490002 208170 490072 208226
rect 489752 208102 490072 208170
rect 489752 208046 489822 208102
rect 489878 208046 489946 208102
rect 490002 208046 490072 208102
rect 489752 207978 490072 208046
rect 489752 207922 489822 207978
rect 489878 207922 489946 207978
rect 490002 207922 490072 207978
rect 489752 207888 490072 207922
rect 498320 208350 498640 208384
rect 498320 208294 498390 208350
rect 498446 208294 498514 208350
rect 498570 208294 498640 208350
rect 498320 208226 498640 208294
rect 498320 208170 498390 208226
rect 498446 208170 498514 208226
rect 498570 208170 498640 208226
rect 498320 208102 498640 208170
rect 498320 208046 498390 208102
rect 498446 208046 498514 208102
rect 498570 208046 498640 208102
rect 498320 207978 498640 208046
rect 498320 207922 498390 207978
rect 498446 207922 498514 207978
rect 498570 207922 498640 207978
rect 498320 207888 498640 207922
rect 506888 208350 507208 208384
rect 506888 208294 506958 208350
rect 507014 208294 507082 208350
rect 507138 208294 507208 208350
rect 506888 208226 507208 208294
rect 506888 208170 506958 208226
rect 507014 208170 507082 208226
rect 507138 208170 507208 208226
rect 506888 208102 507208 208170
rect 506888 208046 506958 208102
rect 507014 208046 507082 208102
rect 507138 208046 507208 208102
rect 506888 207978 507208 208046
rect 506888 207922 506958 207978
rect 507014 207922 507082 207978
rect 507138 207922 507208 207978
rect 506888 207888 507208 207922
rect 515456 208350 515776 208384
rect 515456 208294 515526 208350
rect 515582 208294 515650 208350
rect 515706 208294 515776 208350
rect 515456 208226 515776 208294
rect 515456 208170 515526 208226
rect 515582 208170 515650 208226
rect 515706 208170 515776 208226
rect 515456 208102 515776 208170
rect 515456 208046 515526 208102
rect 515582 208046 515650 208102
rect 515706 208046 515776 208102
rect 515456 207978 515776 208046
rect 515456 207922 515526 207978
rect 515582 207922 515650 207978
rect 515706 207922 515776 207978
rect 515456 207888 515776 207922
rect 519148 205044 519204 236684
rect 519148 204978 519204 204988
rect 527658 220350 528278 237922
rect 527658 220294 527754 220350
rect 527810 220294 527878 220350
rect 527934 220294 528002 220350
rect 528058 220294 528126 220350
rect 528182 220294 528278 220350
rect 527658 220226 528278 220294
rect 527658 220170 527754 220226
rect 527810 220170 527878 220226
rect 527934 220170 528002 220226
rect 528058 220170 528126 220226
rect 528182 220170 528278 220226
rect 527658 220102 528278 220170
rect 527658 220046 527754 220102
rect 527810 220046 527878 220102
rect 527934 220046 528002 220102
rect 528058 220046 528126 220102
rect 528182 220046 528278 220102
rect 527658 219978 528278 220046
rect 527658 219922 527754 219978
rect 527810 219922 527878 219978
rect 527934 219922 528002 219978
rect 528058 219922 528126 219978
rect 528182 219922 528278 219978
rect 481292 198034 481348 198044
rect 496938 202350 497558 203170
rect 496938 202294 497034 202350
rect 497090 202294 497158 202350
rect 497214 202294 497282 202350
rect 497338 202294 497406 202350
rect 497462 202294 497558 202350
rect 496938 202226 497558 202294
rect 496938 202170 497034 202226
rect 497090 202170 497158 202226
rect 497214 202170 497282 202226
rect 497338 202170 497406 202226
rect 497462 202170 497558 202226
rect 496938 202102 497558 202170
rect 496938 202046 497034 202102
rect 497090 202046 497158 202102
rect 497214 202046 497282 202102
rect 497338 202046 497406 202102
rect 497462 202046 497558 202102
rect 496938 201978 497558 202046
rect 496938 201922 497034 201978
rect 497090 201922 497158 201978
rect 497214 201922 497282 201978
rect 497338 201922 497406 201978
rect 497462 201922 497558 201978
rect 479612 197692 479668 197702
rect 469938 190294 470034 190350
rect 470090 190294 470158 190350
rect 470214 190294 470282 190350
rect 470338 190294 470406 190350
rect 470462 190294 470558 190350
rect 469938 190226 470558 190294
rect 469938 190170 470034 190226
rect 470090 190170 470158 190226
rect 470214 190170 470282 190226
rect 470338 190170 470406 190226
rect 470462 190170 470558 190226
rect 469938 190102 470558 190170
rect 469938 190046 470034 190102
rect 470090 190046 470158 190102
rect 470214 190046 470282 190102
rect 470338 190046 470406 190102
rect 470462 190046 470558 190102
rect 469938 189978 470558 190046
rect 469938 189922 470034 189978
rect 470090 189922 470158 189978
rect 470214 189922 470282 189978
rect 470338 189922 470406 189978
rect 470462 189922 470558 189978
rect 469938 172350 470558 189922
rect 469938 172294 470034 172350
rect 470090 172294 470158 172350
rect 470214 172294 470282 172350
rect 470338 172294 470406 172350
rect 470462 172294 470558 172350
rect 469938 172226 470558 172294
rect 469938 172170 470034 172226
rect 470090 172170 470158 172226
rect 470214 172170 470282 172226
rect 470338 172170 470406 172226
rect 470462 172170 470558 172226
rect 469938 172102 470558 172170
rect 469938 172046 470034 172102
rect 470090 172046 470158 172102
rect 470214 172046 470282 172102
rect 470338 172046 470406 172102
rect 470462 172046 470558 172102
rect 469938 171978 470558 172046
rect 469938 171922 470034 171978
rect 470090 171922 470158 171978
rect 470214 171922 470282 171978
rect 470338 171922 470406 171978
rect 470462 171922 470558 171978
rect 469938 154350 470558 171922
rect 469938 154294 470034 154350
rect 470090 154294 470158 154350
rect 470214 154294 470282 154350
rect 470338 154294 470406 154350
rect 470462 154294 470558 154350
rect 469938 154226 470558 154294
rect 469938 154170 470034 154226
rect 470090 154170 470158 154226
rect 470214 154170 470282 154226
rect 470338 154170 470406 154226
rect 470462 154170 470558 154226
rect 469938 154102 470558 154170
rect 469938 154046 470034 154102
rect 470090 154046 470158 154102
rect 470214 154046 470282 154102
rect 470338 154046 470406 154102
rect 470462 154046 470558 154102
rect 469938 153978 470558 154046
rect 469938 153922 470034 153978
rect 470090 153922 470158 153978
rect 470214 153922 470282 153978
rect 470338 153922 470406 153978
rect 470462 153922 470558 153978
rect 469938 149870 470558 153922
rect 496938 184350 497558 201922
rect 497644 198212 497700 198222
rect 497644 198118 497700 198156
rect 497644 198052 497700 198062
rect 499100 198212 499156 198222
rect 499100 197938 499156 198156
rect 499100 197872 499156 197882
rect 496938 184294 497034 184350
rect 497090 184294 497158 184350
rect 497214 184294 497282 184350
rect 497338 184294 497406 184350
rect 497462 184294 497558 184350
rect 496938 184226 497558 184294
rect 496938 184170 497034 184226
rect 497090 184170 497158 184226
rect 497214 184170 497282 184226
rect 497338 184170 497406 184226
rect 497462 184170 497558 184226
rect 496938 184102 497558 184170
rect 496938 184046 497034 184102
rect 497090 184046 497158 184102
rect 497214 184046 497282 184102
rect 497338 184046 497406 184102
rect 497462 184046 497558 184102
rect 496938 183978 497558 184046
rect 496938 183922 497034 183978
rect 497090 183922 497158 183978
rect 497214 183922 497282 183978
rect 497338 183922 497406 183978
rect 497462 183922 497558 183978
rect 496938 166350 497558 183922
rect 496938 166294 497034 166350
rect 497090 166294 497158 166350
rect 497214 166294 497282 166350
rect 497338 166294 497406 166350
rect 497462 166294 497558 166350
rect 496938 166226 497558 166294
rect 496938 166170 497034 166226
rect 497090 166170 497158 166226
rect 497214 166170 497282 166226
rect 497338 166170 497406 166226
rect 497462 166170 497558 166226
rect 496938 166102 497558 166170
rect 496938 166046 497034 166102
rect 497090 166046 497158 166102
rect 497214 166046 497282 166102
rect 497338 166046 497406 166102
rect 497462 166046 497558 166102
rect 496938 165978 497558 166046
rect 496938 165922 497034 165978
rect 497090 165922 497158 165978
rect 497214 165922 497282 165978
rect 497338 165922 497406 165978
rect 497462 165922 497558 165978
rect 495852 153658 495908 153668
rect 495852 152964 495908 153602
rect 495852 152898 495908 152908
rect 496938 149870 497558 165922
rect 500658 190350 501278 203170
rect 527658 202350 528278 219922
rect 527658 202294 527754 202350
rect 527810 202294 527878 202350
rect 527934 202294 528002 202350
rect 528058 202294 528126 202350
rect 528182 202294 528278 202350
rect 527658 202226 528278 202294
rect 527658 202170 527754 202226
rect 527810 202170 527878 202226
rect 527934 202170 528002 202226
rect 528058 202170 528126 202226
rect 528182 202170 528278 202226
rect 527658 202102 528278 202170
rect 527658 202046 527754 202102
rect 527810 202046 527878 202102
rect 527934 202046 528002 202102
rect 528058 202046 528126 202102
rect 528182 202046 528278 202102
rect 527658 201978 528278 202046
rect 527658 201922 527754 201978
rect 527810 201922 527878 201978
rect 527934 201922 528002 201978
rect 528058 201922 528126 201978
rect 528182 201922 528278 201978
rect 516236 201684 516292 201694
rect 516236 199444 516292 201628
rect 516236 199378 516292 199388
rect 502236 198212 502292 198222
rect 502236 197758 502292 198156
rect 502236 197692 502292 197702
rect 500658 190294 500754 190350
rect 500810 190294 500878 190350
rect 500934 190294 501002 190350
rect 501058 190294 501126 190350
rect 501182 190294 501278 190350
rect 500658 190226 501278 190294
rect 500658 190170 500754 190226
rect 500810 190170 500878 190226
rect 500934 190170 501002 190226
rect 501058 190170 501126 190226
rect 501182 190170 501278 190226
rect 500658 190102 501278 190170
rect 500658 190046 500754 190102
rect 500810 190046 500878 190102
rect 500934 190046 501002 190102
rect 501058 190046 501126 190102
rect 501182 190046 501278 190102
rect 500658 189978 501278 190046
rect 500658 189922 500754 189978
rect 500810 189922 500878 189978
rect 500934 189922 501002 189978
rect 501058 189922 501126 189978
rect 501182 189922 501278 189978
rect 500658 172350 501278 189922
rect 500658 172294 500754 172350
rect 500810 172294 500878 172350
rect 500934 172294 501002 172350
rect 501058 172294 501126 172350
rect 501182 172294 501278 172350
rect 500658 172226 501278 172294
rect 500658 172170 500754 172226
rect 500810 172170 500878 172226
rect 500934 172170 501002 172226
rect 501058 172170 501126 172226
rect 501182 172170 501278 172226
rect 500658 172102 501278 172170
rect 500658 172046 500754 172102
rect 500810 172046 500878 172102
rect 500934 172046 501002 172102
rect 501058 172046 501126 172102
rect 501182 172046 501278 172102
rect 500658 171978 501278 172046
rect 500658 171922 500754 171978
rect 500810 171922 500878 171978
rect 500934 171922 501002 171978
rect 501058 171922 501126 171978
rect 501182 171922 501278 171978
rect 500658 154350 501278 171922
rect 500658 154294 500754 154350
rect 500810 154294 500878 154350
rect 500934 154294 501002 154350
rect 501058 154294 501126 154350
rect 501182 154294 501278 154350
rect 500658 154226 501278 154294
rect 500658 154170 500754 154226
rect 500810 154170 500878 154226
rect 500934 154170 501002 154226
rect 501058 154170 501126 154226
rect 501182 154170 501278 154226
rect 500658 154102 501278 154170
rect 500658 154046 500754 154102
rect 500810 154046 500878 154102
rect 500934 154046 501002 154102
rect 501058 154046 501126 154102
rect 501182 154046 501278 154102
rect 500658 153978 501278 154046
rect 500658 153922 500754 153978
rect 500810 153922 500878 153978
rect 500934 153922 501002 153978
rect 501058 153922 501126 153978
rect 501182 153922 501278 153978
rect 500658 149870 501278 153922
rect 527658 184350 528278 201922
rect 527658 184294 527754 184350
rect 527810 184294 527878 184350
rect 527934 184294 528002 184350
rect 528058 184294 528126 184350
rect 528182 184294 528278 184350
rect 527658 184226 528278 184294
rect 527658 184170 527754 184226
rect 527810 184170 527878 184226
rect 527934 184170 528002 184226
rect 528058 184170 528126 184226
rect 528182 184170 528278 184226
rect 527658 184102 528278 184170
rect 527658 184046 527754 184102
rect 527810 184046 527878 184102
rect 527934 184046 528002 184102
rect 528058 184046 528126 184102
rect 528182 184046 528278 184102
rect 527658 183978 528278 184046
rect 527658 183922 527754 183978
rect 527810 183922 527878 183978
rect 527934 183922 528002 183978
rect 528058 183922 528126 183978
rect 528182 183922 528278 183978
rect 527658 166350 528278 183922
rect 527658 166294 527754 166350
rect 527810 166294 527878 166350
rect 527934 166294 528002 166350
rect 528058 166294 528126 166350
rect 528182 166294 528278 166350
rect 527658 166226 528278 166294
rect 527658 166170 527754 166226
rect 527810 166170 527878 166226
rect 527934 166170 528002 166226
rect 528058 166170 528126 166226
rect 528182 166170 528278 166226
rect 527658 166102 528278 166170
rect 527658 166046 527754 166102
rect 527810 166046 527878 166102
rect 527934 166046 528002 166102
rect 528058 166046 528126 166102
rect 528182 166046 528278 166102
rect 527658 165978 528278 166046
rect 527658 165922 527754 165978
rect 527810 165922 527878 165978
rect 527934 165922 528002 165978
rect 528058 165922 528126 165978
rect 528182 165922 528278 165978
rect 501340 152964 501396 152976
rect 501340 152872 501396 152882
rect 527658 149870 528278 165922
rect 531378 406350 531998 408578
rect 545580 407540 545636 590492
rect 546028 409220 546084 590604
rect 558378 580350 558998 596784
rect 558378 580294 558474 580350
rect 558530 580294 558598 580350
rect 558654 580294 558722 580350
rect 558778 580294 558846 580350
rect 558902 580294 558998 580350
rect 558378 580226 558998 580294
rect 558378 580170 558474 580226
rect 558530 580170 558598 580226
rect 558654 580170 558722 580226
rect 558778 580170 558846 580226
rect 558902 580170 558998 580226
rect 558378 580102 558998 580170
rect 558378 580046 558474 580102
rect 558530 580046 558598 580102
rect 558654 580046 558722 580102
rect 558778 580046 558846 580102
rect 558902 580046 558998 580102
rect 558378 579978 558998 580046
rect 558378 579922 558474 579978
rect 558530 579922 558598 579978
rect 558654 579922 558722 579978
rect 558778 579922 558846 579978
rect 558902 579922 558998 579978
rect 558378 562350 558998 579922
rect 558378 562294 558474 562350
rect 558530 562294 558598 562350
rect 558654 562294 558722 562350
rect 558778 562294 558846 562350
rect 558902 562294 558998 562350
rect 558378 562226 558998 562294
rect 558378 562170 558474 562226
rect 558530 562170 558598 562226
rect 558654 562170 558722 562226
rect 558778 562170 558846 562226
rect 558902 562170 558998 562226
rect 558378 562102 558998 562170
rect 558378 562046 558474 562102
rect 558530 562046 558598 562102
rect 558654 562046 558722 562102
rect 558778 562046 558846 562102
rect 558902 562046 558998 562102
rect 558378 561978 558998 562046
rect 558378 561922 558474 561978
rect 558530 561922 558598 561978
rect 558654 561922 558722 561978
rect 558778 561922 558846 561978
rect 558902 561922 558998 561978
rect 547728 550350 548048 550384
rect 547728 550294 547798 550350
rect 547854 550294 547922 550350
rect 547978 550294 548048 550350
rect 547728 550226 548048 550294
rect 547728 550170 547798 550226
rect 547854 550170 547922 550226
rect 547978 550170 548048 550226
rect 547728 550102 548048 550170
rect 547728 550046 547798 550102
rect 547854 550046 547922 550102
rect 547978 550046 548048 550102
rect 547728 549978 548048 550046
rect 547728 549922 547798 549978
rect 547854 549922 547922 549978
rect 547978 549922 548048 549978
rect 547728 549888 548048 549922
rect 558378 544350 558998 561922
rect 558378 544294 558474 544350
rect 558530 544294 558598 544350
rect 558654 544294 558722 544350
rect 558778 544294 558846 544350
rect 558902 544294 558998 544350
rect 558378 544226 558998 544294
rect 558378 544170 558474 544226
rect 558530 544170 558598 544226
rect 558654 544170 558722 544226
rect 558778 544170 558846 544226
rect 558902 544170 558998 544226
rect 558378 544102 558998 544170
rect 558378 544046 558474 544102
rect 558530 544046 558598 544102
rect 558654 544046 558722 544102
rect 558778 544046 558846 544102
rect 558902 544046 558998 544102
rect 558378 543978 558998 544046
rect 558378 543922 558474 543978
rect 558530 543922 558598 543978
rect 558654 543922 558722 543978
rect 558778 543922 558846 543978
rect 558902 543922 558998 543978
rect 547728 532350 548048 532384
rect 547728 532294 547798 532350
rect 547854 532294 547922 532350
rect 547978 532294 548048 532350
rect 547728 532226 548048 532294
rect 547728 532170 547798 532226
rect 547854 532170 547922 532226
rect 547978 532170 548048 532226
rect 547728 532102 548048 532170
rect 547728 532046 547798 532102
rect 547854 532046 547922 532102
rect 547978 532046 548048 532102
rect 547728 531978 548048 532046
rect 547728 531922 547798 531978
rect 547854 531922 547922 531978
rect 547978 531922 548048 531978
rect 547728 531888 548048 531922
rect 558378 526350 558998 543922
rect 558378 526294 558474 526350
rect 558530 526294 558598 526350
rect 558654 526294 558722 526350
rect 558778 526294 558846 526350
rect 558902 526294 558998 526350
rect 558378 526226 558998 526294
rect 558378 526170 558474 526226
rect 558530 526170 558598 526226
rect 558654 526170 558722 526226
rect 558778 526170 558846 526226
rect 558902 526170 558998 526226
rect 558378 526102 558998 526170
rect 558378 526046 558474 526102
rect 558530 526046 558598 526102
rect 558654 526046 558722 526102
rect 558778 526046 558846 526102
rect 558902 526046 558998 526102
rect 558378 525978 558998 526046
rect 558378 525922 558474 525978
rect 558530 525922 558598 525978
rect 558654 525922 558722 525978
rect 558778 525922 558846 525978
rect 558902 525922 558998 525978
rect 547728 514350 548048 514384
rect 547728 514294 547798 514350
rect 547854 514294 547922 514350
rect 547978 514294 548048 514350
rect 547728 514226 548048 514294
rect 547728 514170 547798 514226
rect 547854 514170 547922 514226
rect 547978 514170 548048 514226
rect 547728 514102 548048 514170
rect 547728 514046 547798 514102
rect 547854 514046 547922 514102
rect 547978 514046 548048 514102
rect 547728 513978 548048 514046
rect 547728 513922 547798 513978
rect 547854 513922 547922 513978
rect 547978 513922 548048 513978
rect 547728 513888 548048 513922
rect 558378 508350 558998 525922
rect 558378 508294 558474 508350
rect 558530 508294 558598 508350
rect 558654 508294 558722 508350
rect 558778 508294 558846 508350
rect 558902 508294 558998 508350
rect 558378 508226 558998 508294
rect 558378 508170 558474 508226
rect 558530 508170 558598 508226
rect 558654 508170 558722 508226
rect 558778 508170 558846 508226
rect 558902 508170 558998 508226
rect 558378 508102 558998 508170
rect 558378 508046 558474 508102
rect 558530 508046 558598 508102
rect 558654 508046 558722 508102
rect 558778 508046 558846 508102
rect 558902 508046 558998 508102
rect 558378 507978 558998 508046
rect 558378 507922 558474 507978
rect 558530 507922 558598 507978
rect 558654 507922 558722 507978
rect 558778 507922 558846 507978
rect 558902 507922 558998 507978
rect 547728 496350 548048 496384
rect 547728 496294 547798 496350
rect 547854 496294 547922 496350
rect 547978 496294 548048 496350
rect 547728 496226 548048 496294
rect 547728 496170 547798 496226
rect 547854 496170 547922 496226
rect 547978 496170 548048 496226
rect 547728 496102 548048 496170
rect 547728 496046 547798 496102
rect 547854 496046 547922 496102
rect 547978 496046 548048 496102
rect 547728 495978 548048 496046
rect 547728 495922 547798 495978
rect 547854 495922 547922 495978
rect 547978 495922 548048 495978
rect 547728 495888 548048 495922
rect 558378 490350 558998 507922
rect 558378 490294 558474 490350
rect 558530 490294 558598 490350
rect 558654 490294 558722 490350
rect 558778 490294 558846 490350
rect 558902 490294 558998 490350
rect 558378 490226 558998 490294
rect 558378 490170 558474 490226
rect 558530 490170 558598 490226
rect 558654 490170 558722 490226
rect 558778 490170 558846 490226
rect 558902 490170 558998 490226
rect 558378 490102 558998 490170
rect 558378 490046 558474 490102
rect 558530 490046 558598 490102
rect 558654 490046 558722 490102
rect 558778 490046 558846 490102
rect 558902 490046 558998 490102
rect 558378 489978 558998 490046
rect 558378 489922 558474 489978
rect 558530 489922 558598 489978
rect 558654 489922 558722 489978
rect 558778 489922 558846 489978
rect 558902 489922 558998 489978
rect 547728 478350 548048 478384
rect 547728 478294 547798 478350
rect 547854 478294 547922 478350
rect 547978 478294 548048 478350
rect 547728 478226 548048 478294
rect 547728 478170 547798 478226
rect 547854 478170 547922 478226
rect 547978 478170 548048 478226
rect 547728 478102 548048 478170
rect 547728 478046 547798 478102
rect 547854 478046 547922 478102
rect 547978 478046 548048 478102
rect 547728 477978 548048 478046
rect 547728 477922 547798 477978
rect 547854 477922 547922 477978
rect 547978 477922 548048 477978
rect 547728 477888 548048 477922
rect 558378 472350 558998 489922
rect 558378 472294 558474 472350
rect 558530 472294 558598 472350
rect 558654 472294 558722 472350
rect 558778 472294 558846 472350
rect 558902 472294 558998 472350
rect 558378 472226 558998 472294
rect 558378 472170 558474 472226
rect 558530 472170 558598 472226
rect 558654 472170 558722 472226
rect 558778 472170 558846 472226
rect 558902 472170 558998 472226
rect 558378 472102 558998 472170
rect 558378 472046 558474 472102
rect 558530 472046 558598 472102
rect 558654 472046 558722 472102
rect 558778 472046 558846 472102
rect 558902 472046 558998 472102
rect 558378 471978 558998 472046
rect 558378 471922 558474 471978
rect 558530 471922 558598 471978
rect 558654 471922 558722 471978
rect 558778 471922 558846 471978
rect 558902 471922 558998 471978
rect 547728 460350 548048 460384
rect 547728 460294 547798 460350
rect 547854 460294 547922 460350
rect 547978 460294 548048 460350
rect 547728 460226 548048 460294
rect 547728 460170 547798 460226
rect 547854 460170 547922 460226
rect 547978 460170 548048 460226
rect 547728 460102 548048 460170
rect 547728 460046 547798 460102
rect 547854 460046 547922 460102
rect 547978 460046 548048 460102
rect 547728 459978 548048 460046
rect 547728 459922 547798 459978
rect 547854 459922 547922 459978
rect 547978 459922 548048 459978
rect 547728 459888 548048 459922
rect 558378 454350 558998 471922
rect 558378 454294 558474 454350
rect 558530 454294 558598 454350
rect 558654 454294 558722 454350
rect 558778 454294 558846 454350
rect 558902 454294 558998 454350
rect 558378 454226 558998 454294
rect 558378 454170 558474 454226
rect 558530 454170 558598 454226
rect 558654 454170 558722 454226
rect 558778 454170 558846 454226
rect 558902 454170 558998 454226
rect 558378 454102 558998 454170
rect 558378 454046 558474 454102
rect 558530 454046 558598 454102
rect 558654 454046 558722 454102
rect 558778 454046 558846 454102
rect 558902 454046 558998 454102
rect 558378 453978 558998 454046
rect 558378 453922 558474 453978
rect 558530 453922 558598 453978
rect 558654 453922 558722 453978
rect 558778 453922 558846 453978
rect 558902 453922 558998 453978
rect 547728 442350 548048 442384
rect 547728 442294 547798 442350
rect 547854 442294 547922 442350
rect 547978 442294 548048 442350
rect 547728 442226 548048 442294
rect 547728 442170 547798 442226
rect 547854 442170 547922 442226
rect 547978 442170 548048 442226
rect 547728 442102 548048 442170
rect 547728 442046 547798 442102
rect 547854 442046 547922 442102
rect 547978 442046 548048 442102
rect 547728 441978 548048 442046
rect 547728 441922 547798 441978
rect 547854 441922 547922 441978
rect 547978 441922 548048 441978
rect 547728 441888 548048 441922
rect 558378 436350 558998 453922
rect 558378 436294 558474 436350
rect 558530 436294 558598 436350
rect 558654 436294 558722 436350
rect 558778 436294 558846 436350
rect 558902 436294 558998 436350
rect 558378 436226 558998 436294
rect 558378 436170 558474 436226
rect 558530 436170 558598 436226
rect 558654 436170 558722 436226
rect 558778 436170 558846 436226
rect 558902 436170 558998 436226
rect 558378 436102 558998 436170
rect 558378 436046 558474 436102
rect 558530 436046 558598 436102
rect 558654 436046 558722 436102
rect 558778 436046 558846 436102
rect 558902 436046 558998 436102
rect 558378 435978 558998 436046
rect 558378 435922 558474 435978
rect 558530 435922 558598 435978
rect 558654 435922 558722 435978
rect 558778 435922 558846 435978
rect 558902 435922 558998 435978
rect 547728 424350 548048 424384
rect 547728 424294 547798 424350
rect 547854 424294 547922 424350
rect 547978 424294 548048 424350
rect 547728 424226 548048 424294
rect 547728 424170 547798 424226
rect 547854 424170 547922 424226
rect 547978 424170 548048 424226
rect 547728 424102 548048 424170
rect 547728 424046 547798 424102
rect 547854 424046 547922 424102
rect 547978 424046 548048 424102
rect 547728 423978 548048 424046
rect 547728 423922 547798 423978
rect 547854 423922 547922 423978
rect 547978 423922 548048 423978
rect 547728 423888 548048 423922
rect 546028 409154 546084 409164
rect 558378 418350 558998 435922
rect 558378 418294 558474 418350
rect 558530 418294 558598 418350
rect 558654 418294 558722 418350
rect 558778 418294 558846 418350
rect 558902 418294 558998 418350
rect 558378 418226 558998 418294
rect 558378 418170 558474 418226
rect 558530 418170 558598 418226
rect 558654 418170 558722 418226
rect 558778 418170 558846 418226
rect 558902 418170 558998 418226
rect 558378 418102 558998 418170
rect 558378 418046 558474 418102
rect 558530 418046 558598 418102
rect 558654 418046 558722 418102
rect 558778 418046 558846 418102
rect 558902 418046 558998 418102
rect 558378 417978 558998 418046
rect 558378 417922 558474 417978
rect 558530 417922 558598 417978
rect 558654 417922 558722 417978
rect 558778 417922 558846 417978
rect 558902 417922 558998 417978
rect 545580 407474 545636 407484
rect 531378 406294 531474 406350
rect 531530 406294 531598 406350
rect 531654 406294 531722 406350
rect 531778 406294 531846 406350
rect 531902 406294 531998 406350
rect 531378 406226 531998 406294
rect 531378 406170 531474 406226
rect 531530 406170 531598 406226
rect 531654 406170 531722 406226
rect 531778 406170 531846 406226
rect 531902 406170 531998 406226
rect 531378 406102 531998 406170
rect 531378 406046 531474 406102
rect 531530 406046 531598 406102
rect 531654 406046 531722 406102
rect 531778 406046 531846 406102
rect 531902 406046 531998 406102
rect 531378 405978 531998 406046
rect 531378 405922 531474 405978
rect 531530 405922 531598 405978
rect 531654 405922 531722 405978
rect 531778 405922 531846 405978
rect 531902 405922 531998 405978
rect 531378 388350 531998 405922
rect 531378 388294 531474 388350
rect 531530 388294 531598 388350
rect 531654 388294 531722 388350
rect 531778 388294 531846 388350
rect 531902 388294 531998 388350
rect 531378 388226 531998 388294
rect 531378 388170 531474 388226
rect 531530 388170 531598 388226
rect 531654 388170 531722 388226
rect 531778 388170 531846 388226
rect 531902 388170 531998 388226
rect 531378 388102 531998 388170
rect 531378 388046 531474 388102
rect 531530 388046 531598 388102
rect 531654 388046 531722 388102
rect 531778 388046 531846 388102
rect 531902 388046 531998 388102
rect 531378 387978 531998 388046
rect 531378 387922 531474 387978
rect 531530 387922 531598 387978
rect 531654 387922 531722 387978
rect 531778 387922 531846 387978
rect 531902 387922 531998 387978
rect 531378 370350 531998 387922
rect 531378 370294 531474 370350
rect 531530 370294 531598 370350
rect 531654 370294 531722 370350
rect 531778 370294 531846 370350
rect 531902 370294 531998 370350
rect 531378 370226 531998 370294
rect 531378 370170 531474 370226
rect 531530 370170 531598 370226
rect 531654 370170 531722 370226
rect 531778 370170 531846 370226
rect 531902 370170 531998 370226
rect 531378 370102 531998 370170
rect 531378 370046 531474 370102
rect 531530 370046 531598 370102
rect 531654 370046 531722 370102
rect 531778 370046 531846 370102
rect 531902 370046 531998 370102
rect 531378 369978 531998 370046
rect 531378 369922 531474 369978
rect 531530 369922 531598 369978
rect 531654 369922 531722 369978
rect 531778 369922 531846 369978
rect 531902 369922 531998 369978
rect 531378 352350 531998 369922
rect 531378 352294 531474 352350
rect 531530 352294 531598 352350
rect 531654 352294 531722 352350
rect 531778 352294 531846 352350
rect 531902 352294 531998 352350
rect 531378 352226 531998 352294
rect 531378 352170 531474 352226
rect 531530 352170 531598 352226
rect 531654 352170 531722 352226
rect 531778 352170 531846 352226
rect 531902 352170 531998 352226
rect 531378 352102 531998 352170
rect 531378 352046 531474 352102
rect 531530 352046 531598 352102
rect 531654 352046 531722 352102
rect 531778 352046 531846 352102
rect 531902 352046 531998 352102
rect 531378 351978 531998 352046
rect 531378 351922 531474 351978
rect 531530 351922 531598 351978
rect 531654 351922 531722 351978
rect 531778 351922 531846 351978
rect 531902 351922 531998 351978
rect 531378 334350 531998 351922
rect 558378 400350 558998 417922
rect 558378 400294 558474 400350
rect 558530 400294 558598 400350
rect 558654 400294 558722 400350
rect 558778 400294 558846 400350
rect 558902 400294 558998 400350
rect 558378 400226 558998 400294
rect 558378 400170 558474 400226
rect 558530 400170 558598 400226
rect 558654 400170 558722 400226
rect 558778 400170 558846 400226
rect 558902 400170 558998 400226
rect 558378 400102 558998 400170
rect 558378 400046 558474 400102
rect 558530 400046 558598 400102
rect 558654 400046 558722 400102
rect 558778 400046 558846 400102
rect 558902 400046 558998 400102
rect 558378 399978 558998 400046
rect 558378 399922 558474 399978
rect 558530 399922 558598 399978
rect 558654 399922 558722 399978
rect 558778 399922 558846 399978
rect 558902 399922 558998 399978
rect 558378 382350 558998 399922
rect 558378 382294 558474 382350
rect 558530 382294 558598 382350
rect 558654 382294 558722 382350
rect 558778 382294 558846 382350
rect 558902 382294 558998 382350
rect 558378 382226 558998 382294
rect 558378 382170 558474 382226
rect 558530 382170 558598 382226
rect 558654 382170 558722 382226
rect 558778 382170 558846 382226
rect 558902 382170 558998 382226
rect 558378 382102 558998 382170
rect 558378 382046 558474 382102
rect 558530 382046 558598 382102
rect 558654 382046 558722 382102
rect 558778 382046 558846 382102
rect 558902 382046 558998 382102
rect 558378 381978 558998 382046
rect 558378 381922 558474 381978
rect 558530 381922 558598 381978
rect 558654 381922 558722 381978
rect 558778 381922 558846 381978
rect 558902 381922 558998 381978
rect 558378 364350 558998 381922
rect 562098 598172 562718 598268
rect 562098 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 562718 598172
rect 562098 598048 562718 598116
rect 562098 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 562718 598048
rect 562098 597924 562718 597992
rect 562098 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 562718 597924
rect 562098 597800 562718 597868
rect 562098 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 562718 597800
rect 562098 586350 562718 597744
rect 562098 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 562718 586350
rect 562098 586226 562718 586294
rect 562098 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 562718 586226
rect 562098 586102 562718 586170
rect 562098 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 562718 586102
rect 562098 585978 562718 586046
rect 562098 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 562718 585978
rect 562098 568350 562718 585922
rect 562098 568294 562194 568350
rect 562250 568294 562318 568350
rect 562374 568294 562442 568350
rect 562498 568294 562566 568350
rect 562622 568294 562718 568350
rect 562098 568226 562718 568294
rect 562098 568170 562194 568226
rect 562250 568170 562318 568226
rect 562374 568170 562442 568226
rect 562498 568170 562566 568226
rect 562622 568170 562718 568226
rect 562098 568102 562718 568170
rect 562098 568046 562194 568102
rect 562250 568046 562318 568102
rect 562374 568046 562442 568102
rect 562498 568046 562566 568102
rect 562622 568046 562718 568102
rect 562098 567978 562718 568046
rect 562098 567922 562194 567978
rect 562250 567922 562318 567978
rect 562374 567922 562442 567978
rect 562498 567922 562566 567978
rect 562622 567922 562718 567978
rect 562098 550350 562718 567922
rect 562098 550294 562194 550350
rect 562250 550294 562318 550350
rect 562374 550294 562442 550350
rect 562498 550294 562566 550350
rect 562622 550294 562718 550350
rect 562098 550226 562718 550294
rect 562098 550170 562194 550226
rect 562250 550170 562318 550226
rect 562374 550170 562442 550226
rect 562498 550170 562566 550226
rect 562622 550170 562718 550226
rect 562098 550102 562718 550170
rect 562098 550046 562194 550102
rect 562250 550046 562318 550102
rect 562374 550046 562442 550102
rect 562498 550046 562566 550102
rect 562622 550046 562718 550102
rect 562098 549978 562718 550046
rect 562098 549922 562194 549978
rect 562250 549922 562318 549978
rect 562374 549922 562442 549978
rect 562498 549922 562566 549978
rect 562622 549922 562718 549978
rect 562098 532350 562718 549922
rect 562098 532294 562194 532350
rect 562250 532294 562318 532350
rect 562374 532294 562442 532350
rect 562498 532294 562566 532350
rect 562622 532294 562718 532350
rect 562098 532226 562718 532294
rect 562098 532170 562194 532226
rect 562250 532170 562318 532226
rect 562374 532170 562442 532226
rect 562498 532170 562566 532226
rect 562622 532170 562718 532226
rect 562098 532102 562718 532170
rect 562098 532046 562194 532102
rect 562250 532046 562318 532102
rect 562374 532046 562442 532102
rect 562498 532046 562566 532102
rect 562622 532046 562718 532102
rect 562098 531978 562718 532046
rect 562098 531922 562194 531978
rect 562250 531922 562318 531978
rect 562374 531922 562442 531978
rect 562498 531922 562566 531978
rect 562622 531922 562718 531978
rect 562098 514350 562718 531922
rect 562098 514294 562194 514350
rect 562250 514294 562318 514350
rect 562374 514294 562442 514350
rect 562498 514294 562566 514350
rect 562622 514294 562718 514350
rect 562098 514226 562718 514294
rect 562098 514170 562194 514226
rect 562250 514170 562318 514226
rect 562374 514170 562442 514226
rect 562498 514170 562566 514226
rect 562622 514170 562718 514226
rect 562098 514102 562718 514170
rect 562098 514046 562194 514102
rect 562250 514046 562318 514102
rect 562374 514046 562442 514102
rect 562498 514046 562566 514102
rect 562622 514046 562718 514102
rect 562098 513978 562718 514046
rect 562098 513922 562194 513978
rect 562250 513922 562318 513978
rect 562374 513922 562442 513978
rect 562498 513922 562566 513978
rect 562622 513922 562718 513978
rect 562098 496350 562718 513922
rect 562098 496294 562194 496350
rect 562250 496294 562318 496350
rect 562374 496294 562442 496350
rect 562498 496294 562566 496350
rect 562622 496294 562718 496350
rect 562098 496226 562718 496294
rect 562098 496170 562194 496226
rect 562250 496170 562318 496226
rect 562374 496170 562442 496226
rect 562498 496170 562566 496226
rect 562622 496170 562718 496226
rect 562098 496102 562718 496170
rect 562098 496046 562194 496102
rect 562250 496046 562318 496102
rect 562374 496046 562442 496102
rect 562498 496046 562566 496102
rect 562622 496046 562718 496102
rect 562098 495978 562718 496046
rect 562098 495922 562194 495978
rect 562250 495922 562318 495978
rect 562374 495922 562442 495978
rect 562498 495922 562566 495978
rect 562622 495922 562718 495978
rect 562098 478350 562718 495922
rect 562098 478294 562194 478350
rect 562250 478294 562318 478350
rect 562374 478294 562442 478350
rect 562498 478294 562566 478350
rect 562622 478294 562718 478350
rect 562098 478226 562718 478294
rect 562098 478170 562194 478226
rect 562250 478170 562318 478226
rect 562374 478170 562442 478226
rect 562498 478170 562566 478226
rect 562622 478170 562718 478226
rect 562098 478102 562718 478170
rect 562098 478046 562194 478102
rect 562250 478046 562318 478102
rect 562374 478046 562442 478102
rect 562498 478046 562566 478102
rect 562622 478046 562718 478102
rect 562098 477978 562718 478046
rect 562098 477922 562194 477978
rect 562250 477922 562318 477978
rect 562374 477922 562442 477978
rect 562498 477922 562566 477978
rect 562622 477922 562718 477978
rect 562098 460350 562718 477922
rect 562098 460294 562194 460350
rect 562250 460294 562318 460350
rect 562374 460294 562442 460350
rect 562498 460294 562566 460350
rect 562622 460294 562718 460350
rect 562098 460226 562718 460294
rect 562098 460170 562194 460226
rect 562250 460170 562318 460226
rect 562374 460170 562442 460226
rect 562498 460170 562566 460226
rect 562622 460170 562718 460226
rect 562098 460102 562718 460170
rect 562098 460046 562194 460102
rect 562250 460046 562318 460102
rect 562374 460046 562442 460102
rect 562498 460046 562566 460102
rect 562622 460046 562718 460102
rect 562098 459978 562718 460046
rect 562098 459922 562194 459978
rect 562250 459922 562318 459978
rect 562374 459922 562442 459978
rect 562498 459922 562566 459978
rect 562622 459922 562718 459978
rect 562098 442350 562718 459922
rect 562098 442294 562194 442350
rect 562250 442294 562318 442350
rect 562374 442294 562442 442350
rect 562498 442294 562566 442350
rect 562622 442294 562718 442350
rect 562098 442226 562718 442294
rect 562098 442170 562194 442226
rect 562250 442170 562318 442226
rect 562374 442170 562442 442226
rect 562498 442170 562566 442226
rect 562622 442170 562718 442226
rect 562098 442102 562718 442170
rect 562098 442046 562194 442102
rect 562250 442046 562318 442102
rect 562374 442046 562442 442102
rect 562498 442046 562566 442102
rect 562622 442046 562718 442102
rect 562098 441978 562718 442046
rect 562098 441922 562194 441978
rect 562250 441922 562318 441978
rect 562374 441922 562442 441978
rect 562498 441922 562566 441978
rect 562622 441922 562718 441978
rect 562098 424350 562718 441922
rect 562098 424294 562194 424350
rect 562250 424294 562318 424350
rect 562374 424294 562442 424350
rect 562498 424294 562566 424350
rect 562622 424294 562718 424350
rect 562098 424226 562718 424294
rect 562098 424170 562194 424226
rect 562250 424170 562318 424226
rect 562374 424170 562442 424226
rect 562498 424170 562566 424226
rect 562622 424170 562718 424226
rect 562098 424102 562718 424170
rect 562098 424046 562194 424102
rect 562250 424046 562318 424102
rect 562374 424046 562442 424102
rect 562498 424046 562566 424102
rect 562622 424046 562718 424102
rect 562098 423978 562718 424046
rect 562098 423922 562194 423978
rect 562250 423922 562318 423978
rect 562374 423922 562442 423978
rect 562498 423922 562566 423978
rect 562622 423922 562718 423978
rect 562098 406350 562718 423922
rect 562098 406294 562194 406350
rect 562250 406294 562318 406350
rect 562374 406294 562442 406350
rect 562498 406294 562566 406350
rect 562622 406294 562718 406350
rect 562098 406226 562718 406294
rect 562098 406170 562194 406226
rect 562250 406170 562318 406226
rect 562374 406170 562442 406226
rect 562498 406170 562566 406226
rect 562622 406170 562718 406226
rect 562098 406102 562718 406170
rect 562098 406046 562194 406102
rect 562250 406046 562318 406102
rect 562374 406046 562442 406102
rect 562498 406046 562566 406102
rect 562622 406046 562718 406102
rect 562098 405978 562718 406046
rect 562098 405922 562194 405978
rect 562250 405922 562318 405978
rect 562374 405922 562442 405978
rect 562498 405922 562566 405978
rect 562622 405922 562718 405978
rect 562098 388350 562718 405922
rect 589098 597212 589718 598268
rect 589098 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 589718 597212
rect 589098 597088 589718 597156
rect 589098 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 589718 597088
rect 589098 596964 589718 597032
rect 589098 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 589718 596964
rect 589098 596840 589718 596908
rect 589098 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 589718 596840
rect 589098 580350 589718 596784
rect 592818 598172 593438 598268
rect 592818 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 593438 598172
rect 592818 598048 593438 598116
rect 592818 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 593438 598048
rect 592818 597924 593438 597992
rect 592818 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 593438 597924
rect 592818 597800 593438 597868
rect 592818 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 593438 597800
rect 589098 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 589718 580350
rect 589098 580226 589718 580294
rect 589098 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 589718 580226
rect 589098 580102 589718 580170
rect 589098 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 589718 580102
rect 589098 579978 589718 580046
rect 589098 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 589718 579978
rect 589098 562350 589718 579922
rect 589098 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 589718 562350
rect 589098 562226 589718 562294
rect 589098 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 589718 562226
rect 589098 562102 589718 562170
rect 589098 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 589718 562102
rect 589098 561978 589718 562046
rect 589098 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 589718 561978
rect 589098 544350 589718 561922
rect 589098 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 589718 544350
rect 589098 544226 589718 544294
rect 589098 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 589718 544226
rect 589098 544102 589718 544170
rect 589098 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 589718 544102
rect 589098 543978 589718 544046
rect 589098 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 589718 543978
rect 589098 526350 589718 543922
rect 589098 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 589718 526350
rect 589098 526226 589718 526294
rect 589098 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 589718 526226
rect 589098 526102 589718 526170
rect 589098 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 589718 526102
rect 589098 525978 589718 526046
rect 589098 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 589718 525978
rect 589098 508350 589718 525922
rect 589098 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 589718 508350
rect 589098 508226 589718 508294
rect 589098 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 589718 508226
rect 589098 508102 589718 508170
rect 589098 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 589718 508102
rect 589098 507978 589718 508046
rect 589098 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 589718 507978
rect 589098 490350 589718 507922
rect 589098 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 589718 490350
rect 589098 490226 589718 490294
rect 589098 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 589718 490226
rect 589098 490102 589718 490170
rect 589098 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 589718 490102
rect 589098 489978 589718 490046
rect 589098 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 589718 489978
rect 589098 472350 589718 489922
rect 589098 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 589718 472350
rect 589098 472226 589718 472294
rect 589098 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 589718 472226
rect 589098 472102 589718 472170
rect 589098 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 589718 472102
rect 589098 471978 589718 472046
rect 589098 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 589718 471978
rect 589098 454350 589718 471922
rect 589098 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 589718 454350
rect 589098 454226 589718 454294
rect 589098 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 589718 454226
rect 589098 454102 589718 454170
rect 589098 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 589718 454102
rect 589098 453978 589718 454046
rect 589098 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 589718 453978
rect 589098 436350 589718 453922
rect 589098 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 589718 436350
rect 589098 436226 589718 436294
rect 589098 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 589718 436226
rect 589098 436102 589718 436170
rect 589098 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 589718 436102
rect 589098 435978 589718 436046
rect 589098 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 589718 435978
rect 589098 418350 589718 435922
rect 589098 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 589718 418350
rect 589098 418226 589718 418294
rect 589098 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 589718 418226
rect 589098 418102 589718 418170
rect 589098 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 589718 418102
rect 589098 417978 589718 418046
rect 589098 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 589718 417978
rect 589098 400350 589718 417922
rect 589098 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 589718 400350
rect 589098 400226 589718 400294
rect 589098 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 589718 400226
rect 589098 400102 589718 400170
rect 589098 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 589718 400102
rect 589098 399978 589718 400046
rect 589098 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 589718 399978
rect 562098 388294 562194 388350
rect 562250 388294 562318 388350
rect 562374 388294 562442 388350
rect 562498 388294 562566 388350
rect 562622 388294 562718 388350
rect 562098 388226 562718 388294
rect 562098 388170 562194 388226
rect 562250 388170 562318 388226
rect 562374 388170 562442 388226
rect 562498 388170 562566 388226
rect 562622 388170 562718 388226
rect 562098 388102 562718 388170
rect 562098 388046 562194 388102
rect 562250 388046 562318 388102
rect 562374 388046 562442 388102
rect 562498 388046 562566 388102
rect 562622 388046 562718 388102
rect 562098 387978 562718 388046
rect 562098 387922 562194 387978
rect 562250 387922 562318 387978
rect 562374 387922 562442 387978
rect 562498 387922 562566 387978
rect 562622 387922 562718 387978
rect 558378 364294 558474 364350
rect 558530 364294 558598 364350
rect 558654 364294 558722 364350
rect 558778 364294 558846 364350
rect 558902 364294 558998 364350
rect 558378 364226 558998 364294
rect 558378 364170 558474 364226
rect 558530 364170 558598 364226
rect 558654 364170 558722 364226
rect 558778 364170 558846 364226
rect 558902 364170 558998 364226
rect 558378 364102 558998 364170
rect 558378 364046 558474 364102
rect 558530 364046 558598 364102
rect 558654 364046 558722 364102
rect 558778 364046 558846 364102
rect 558902 364046 558998 364102
rect 558378 363978 558998 364046
rect 558378 363922 558474 363978
rect 558530 363922 558598 363978
rect 558654 363922 558722 363978
rect 558778 363922 558846 363978
rect 558902 363922 558998 363978
rect 558378 346350 558998 363922
rect 558378 346294 558474 346350
rect 558530 346294 558598 346350
rect 558654 346294 558722 346350
rect 558778 346294 558846 346350
rect 558902 346294 558998 346350
rect 558378 346226 558998 346294
rect 558378 346170 558474 346226
rect 558530 346170 558598 346226
rect 558654 346170 558722 346226
rect 558778 346170 558846 346226
rect 558902 346170 558998 346226
rect 558378 346102 558998 346170
rect 558378 346046 558474 346102
rect 558530 346046 558598 346102
rect 558654 346046 558722 346102
rect 558778 346046 558846 346102
rect 558902 346046 558998 346102
rect 558378 345978 558998 346046
rect 558378 345922 558474 345978
rect 558530 345922 558598 345978
rect 558654 345922 558722 345978
rect 558778 345922 558846 345978
rect 558902 345922 558998 345978
rect 531378 334294 531474 334350
rect 531530 334294 531598 334350
rect 531654 334294 531722 334350
rect 531778 334294 531846 334350
rect 531902 334294 531998 334350
rect 531378 334226 531998 334294
rect 531378 334170 531474 334226
rect 531530 334170 531598 334226
rect 531654 334170 531722 334226
rect 531778 334170 531846 334226
rect 531902 334170 531998 334226
rect 531378 334102 531998 334170
rect 531378 334046 531474 334102
rect 531530 334046 531598 334102
rect 531654 334046 531722 334102
rect 531778 334046 531846 334102
rect 531902 334046 531998 334102
rect 531378 333978 531998 334046
rect 531378 333922 531474 333978
rect 531530 333922 531598 333978
rect 531654 333922 531722 333978
rect 531778 333922 531846 333978
rect 531902 333922 531998 333978
rect 531378 316350 531998 333922
rect 531378 316294 531474 316350
rect 531530 316294 531598 316350
rect 531654 316294 531722 316350
rect 531778 316294 531846 316350
rect 531902 316294 531998 316350
rect 531378 316226 531998 316294
rect 531378 316170 531474 316226
rect 531530 316170 531598 316226
rect 531654 316170 531722 316226
rect 531778 316170 531846 316226
rect 531902 316170 531998 316226
rect 531378 316102 531998 316170
rect 531378 316046 531474 316102
rect 531530 316046 531598 316102
rect 531654 316046 531722 316102
rect 531778 316046 531846 316102
rect 531902 316046 531998 316102
rect 531378 315978 531998 316046
rect 531378 315922 531474 315978
rect 531530 315922 531598 315978
rect 531654 315922 531722 315978
rect 531778 315922 531846 315978
rect 531902 315922 531998 315978
rect 531378 298350 531998 315922
rect 531378 298294 531474 298350
rect 531530 298294 531598 298350
rect 531654 298294 531722 298350
rect 531778 298294 531846 298350
rect 531902 298294 531998 298350
rect 531378 298226 531998 298294
rect 531378 298170 531474 298226
rect 531530 298170 531598 298226
rect 531654 298170 531722 298226
rect 531778 298170 531846 298226
rect 531902 298170 531998 298226
rect 531378 298102 531998 298170
rect 531378 298046 531474 298102
rect 531530 298046 531598 298102
rect 531654 298046 531722 298102
rect 531778 298046 531846 298102
rect 531902 298046 531998 298102
rect 531378 297978 531998 298046
rect 531378 297922 531474 297978
rect 531530 297922 531598 297978
rect 531654 297922 531722 297978
rect 531778 297922 531846 297978
rect 531902 297922 531998 297978
rect 531378 280350 531998 297922
rect 531378 280294 531474 280350
rect 531530 280294 531598 280350
rect 531654 280294 531722 280350
rect 531778 280294 531846 280350
rect 531902 280294 531998 280350
rect 531378 280226 531998 280294
rect 531378 280170 531474 280226
rect 531530 280170 531598 280226
rect 531654 280170 531722 280226
rect 531778 280170 531846 280226
rect 531902 280170 531998 280226
rect 531378 280102 531998 280170
rect 531378 280046 531474 280102
rect 531530 280046 531598 280102
rect 531654 280046 531722 280102
rect 531778 280046 531846 280102
rect 531902 280046 531998 280102
rect 531378 279978 531998 280046
rect 531378 279922 531474 279978
rect 531530 279922 531598 279978
rect 531654 279922 531722 279978
rect 531778 279922 531846 279978
rect 531902 279922 531998 279978
rect 531378 262350 531998 279922
rect 531378 262294 531474 262350
rect 531530 262294 531598 262350
rect 531654 262294 531722 262350
rect 531778 262294 531846 262350
rect 531902 262294 531998 262350
rect 531378 262226 531998 262294
rect 531378 262170 531474 262226
rect 531530 262170 531598 262226
rect 531654 262170 531722 262226
rect 531778 262170 531846 262226
rect 531902 262170 531998 262226
rect 531378 262102 531998 262170
rect 531378 262046 531474 262102
rect 531530 262046 531598 262102
rect 531654 262046 531722 262102
rect 531778 262046 531846 262102
rect 531902 262046 531998 262102
rect 531378 261978 531998 262046
rect 531378 261922 531474 261978
rect 531530 261922 531598 261978
rect 531654 261922 531722 261978
rect 531778 261922 531846 261978
rect 531902 261922 531998 261978
rect 531378 244350 531998 261922
rect 531378 244294 531474 244350
rect 531530 244294 531598 244350
rect 531654 244294 531722 244350
rect 531778 244294 531846 244350
rect 531902 244294 531998 244350
rect 531378 244226 531998 244294
rect 531378 244170 531474 244226
rect 531530 244170 531598 244226
rect 531654 244170 531722 244226
rect 531778 244170 531846 244226
rect 531902 244170 531998 244226
rect 531378 244102 531998 244170
rect 531378 244046 531474 244102
rect 531530 244046 531598 244102
rect 531654 244046 531722 244102
rect 531778 244046 531846 244102
rect 531902 244046 531998 244102
rect 531378 243978 531998 244046
rect 531378 243922 531474 243978
rect 531530 243922 531598 243978
rect 531654 243922 531722 243978
rect 531778 243922 531846 243978
rect 531902 243922 531998 243978
rect 531378 226350 531998 243922
rect 531378 226294 531474 226350
rect 531530 226294 531598 226350
rect 531654 226294 531722 226350
rect 531778 226294 531846 226350
rect 531902 226294 531998 226350
rect 531378 226226 531998 226294
rect 531378 226170 531474 226226
rect 531530 226170 531598 226226
rect 531654 226170 531722 226226
rect 531778 226170 531846 226226
rect 531902 226170 531998 226226
rect 531378 226102 531998 226170
rect 531378 226046 531474 226102
rect 531530 226046 531598 226102
rect 531654 226046 531722 226102
rect 531778 226046 531846 226102
rect 531902 226046 531998 226102
rect 531378 225978 531998 226046
rect 531378 225922 531474 225978
rect 531530 225922 531598 225978
rect 531654 225922 531722 225978
rect 531778 225922 531846 225978
rect 531902 225922 531998 225978
rect 531378 208350 531998 225922
rect 531378 208294 531474 208350
rect 531530 208294 531598 208350
rect 531654 208294 531722 208350
rect 531778 208294 531846 208350
rect 531902 208294 531998 208350
rect 531378 208226 531998 208294
rect 531378 208170 531474 208226
rect 531530 208170 531598 208226
rect 531654 208170 531722 208226
rect 531778 208170 531846 208226
rect 531902 208170 531998 208226
rect 531378 208102 531998 208170
rect 531378 208046 531474 208102
rect 531530 208046 531598 208102
rect 531654 208046 531722 208102
rect 531778 208046 531846 208102
rect 531902 208046 531998 208102
rect 531378 207978 531998 208046
rect 531378 207922 531474 207978
rect 531530 207922 531598 207978
rect 531654 207922 531722 207978
rect 531778 207922 531846 207978
rect 531902 207922 531998 207978
rect 531378 190350 531998 207922
rect 531378 190294 531474 190350
rect 531530 190294 531598 190350
rect 531654 190294 531722 190350
rect 531778 190294 531846 190350
rect 531902 190294 531998 190350
rect 531378 190226 531998 190294
rect 531378 190170 531474 190226
rect 531530 190170 531598 190226
rect 531654 190170 531722 190226
rect 531778 190170 531846 190226
rect 531902 190170 531998 190226
rect 531378 190102 531998 190170
rect 531378 190046 531474 190102
rect 531530 190046 531598 190102
rect 531654 190046 531722 190102
rect 531778 190046 531846 190102
rect 531902 190046 531998 190102
rect 531378 189978 531998 190046
rect 531378 189922 531474 189978
rect 531530 189922 531598 189978
rect 531654 189922 531722 189978
rect 531778 189922 531846 189978
rect 531902 189922 531998 189978
rect 531378 172350 531998 189922
rect 531378 172294 531474 172350
rect 531530 172294 531598 172350
rect 531654 172294 531722 172350
rect 531778 172294 531846 172350
rect 531902 172294 531998 172350
rect 531378 172226 531998 172294
rect 531378 172170 531474 172226
rect 531530 172170 531598 172226
rect 531654 172170 531722 172226
rect 531778 172170 531846 172226
rect 531902 172170 531998 172226
rect 531378 172102 531998 172170
rect 531378 172046 531474 172102
rect 531530 172046 531598 172102
rect 531654 172046 531722 172102
rect 531778 172046 531846 172102
rect 531902 172046 531998 172102
rect 531378 171978 531998 172046
rect 531378 171922 531474 171978
rect 531530 171922 531598 171978
rect 531654 171922 531722 171978
rect 531778 171922 531846 171978
rect 531902 171922 531998 171978
rect 531378 154350 531998 171922
rect 531378 154294 531474 154350
rect 531530 154294 531598 154350
rect 531654 154294 531722 154350
rect 531778 154294 531846 154350
rect 531902 154294 531998 154350
rect 531378 154226 531998 154294
rect 531378 154170 531474 154226
rect 531530 154170 531598 154226
rect 531654 154170 531722 154226
rect 531778 154170 531846 154226
rect 531902 154170 531998 154226
rect 531378 154102 531998 154170
rect 531378 154046 531474 154102
rect 531530 154046 531598 154102
rect 531654 154046 531722 154102
rect 531778 154046 531846 154102
rect 531902 154046 531998 154102
rect 531378 153978 531998 154046
rect 531378 153922 531474 153978
rect 531530 153922 531598 153978
rect 531654 153922 531722 153978
rect 531778 153922 531846 153978
rect 531902 153922 531998 153978
rect 531378 149870 531998 153922
rect 540092 342132 540148 342142
rect 465500 149492 465556 149502
rect 465500 149156 465556 149436
rect 465500 149090 465556 149100
rect 509740 149492 509796 149502
rect 509740 149156 509796 149436
rect 509740 149090 509796 149100
rect 540092 148708 540148 342076
rect 540092 148642 540148 148652
rect 555212 341012 555268 341022
rect 555212 148148 555268 340956
rect 555212 148082 555268 148092
rect 556892 339892 556948 339902
rect 556892 148036 556948 339836
rect 558378 328350 558998 345922
rect 560252 371252 560308 371262
rect 559580 345492 559636 345502
rect 558378 328294 558474 328350
rect 558530 328294 558598 328350
rect 558654 328294 558722 328350
rect 558778 328294 558846 328350
rect 558902 328294 558998 328350
rect 558378 328226 558998 328294
rect 558378 328170 558474 328226
rect 558530 328170 558598 328226
rect 558654 328170 558722 328226
rect 558778 328170 558846 328226
rect 558902 328170 558998 328226
rect 558378 328102 558998 328170
rect 558378 328046 558474 328102
rect 558530 328046 558598 328102
rect 558654 328046 558722 328102
rect 558778 328046 558846 328102
rect 558902 328046 558998 328102
rect 558378 327978 558998 328046
rect 558378 327922 558474 327978
rect 558530 327922 558598 327978
rect 558654 327922 558722 327978
rect 558778 327922 558846 327978
rect 558902 327922 558998 327978
rect 558378 310350 558998 327922
rect 558378 310294 558474 310350
rect 558530 310294 558598 310350
rect 558654 310294 558722 310350
rect 558778 310294 558846 310350
rect 558902 310294 558998 310350
rect 558378 310226 558998 310294
rect 558378 310170 558474 310226
rect 558530 310170 558598 310226
rect 558654 310170 558722 310226
rect 558778 310170 558846 310226
rect 558902 310170 558998 310226
rect 558378 310102 558998 310170
rect 558378 310046 558474 310102
rect 558530 310046 558598 310102
rect 558654 310046 558722 310102
rect 558778 310046 558846 310102
rect 558902 310046 558998 310102
rect 558378 309978 558998 310046
rect 558378 309922 558474 309978
rect 558530 309922 558598 309978
rect 558654 309922 558722 309978
rect 558778 309922 558846 309978
rect 558902 309922 558998 309978
rect 558378 292350 558998 309922
rect 558378 292294 558474 292350
rect 558530 292294 558598 292350
rect 558654 292294 558722 292350
rect 558778 292294 558846 292350
rect 558902 292294 558998 292350
rect 558378 292226 558998 292294
rect 558378 292170 558474 292226
rect 558530 292170 558598 292226
rect 558654 292170 558722 292226
rect 558778 292170 558846 292226
rect 558902 292170 558998 292226
rect 558378 292102 558998 292170
rect 558378 292046 558474 292102
rect 558530 292046 558598 292102
rect 558654 292046 558722 292102
rect 558778 292046 558846 292102
rect 558902 292046 558998 292102
rect 558378 291978 558998 292046
rect 558378 291922 558474 291978
rect 558530 291922 558598 291978
rect 558654 291922 558722 291978
rect 558778 291922 558846 291978
rect 558902 291922 558998 291978
rect 558378 274350 558998 291922
rect 558378 274294 558474 274350
rect 558530 274294 558598 274350
rect 558654 274294 558722 274350
rect 558778 274294 558846 274350
rect 558902 274294 558998 274350
rect 558378 274226 558998 274294
rect 558378 274170 558474 274226
rect 558530 274170 558598 274226
rect 558654 274170 558722 274226
rect 558778 274170 558846 274226
rect 558902 274170 558998 274226
rect 558378 274102 558998 274170
rect 558378 274046 558474 274102
rect 558530 274046 558598 274102
rect 558654 274046 558722 274102
rect 558778 274046 558846 274102
rect 558902 274046 558998 274102
rect 558378 273978 558998 274046
rect 558378 273922 558474 273978
rect 558530 273922 558598 273978
rect 558654 273922 558722 273978
rect 558778 273922 558846 273978
rect 558902 273922 558998 273978
rect 558378 256350 558998 273922
rect 558378 256294 558474 256350
rect 558530 256294 558598 256350
rect 558654 256294 558722 256350
rect 558778 256294 558846 256350
rect 558902 256294 558998 256350
rect 558378 256226 558998 256294
rect 558378 256170 558474 256226
rect 558530 256170 558598 256226
rect 558654 256170 558722 256226
rect 558778 256170 558846 256226
rect 558902 256170 558998 256226
rect 558378 256102 558998 256170
rect 558378 256046 558474 256102
rect 558530 256046 558598 256102
rect 558654 256046 558722 256102
rect 558778 256046 558846 256102
rect 558902 256046 558998 256102
rect 558378 255978 558998 256046
rect 558378 255922 558474 255978
rect 558530 255922 558598 255978
rect 558654 255922 558722 255978
rect 558778 255922 558846 255978
rect 558902 255922 558998 255978
rect 558378 238350 558998 255922
rect 558378 238294 558474 238350
rect 558530 238294 558598 238350
rect 558654 238294 558722 238350
rect 558778 238294 558846 238350
rect 558902 238294 558998 238350
rect 558378 238226 558998 238294
rect 558378 238170 558474 238226
rect 558530 238170 558598 238226
rect 558654 238170 558722 238226
rect 558778 238170 558846 238226
rect 558902 238170 558998 238226
rect 558378 238102 558998 238170
rect 558378 238046 558474 238102
rect 558530 238046 558598 238102
rect 558654 238046 558722 238102
rect 558778 238046 558846 238102
rect 558902 238046 558998 238102
rect 558378 237978 558998 238046
rect 558378 237922 558474 237978
rect 558530 237922 558598 237978
rect 558654 237922 558722 237978
rect 558778 237922 558846 237978
rect 558902 237922 558998 237978
rect 558378 220350 558998 237922
rect 558378 220294 558474 220350
rect 558530 220294 558598 220350
rect 558654 220294 558722 220350
rect 558778 220294 558846 220350
rect 558902 220294 558998 220350
rect 558378 220226 558998 220294
rect 558378 220170 558474 220226
rect 558530 220170 558598 220226
rect 558654 220170 558722 220226
rect 558778 220170 558846 220226
rect 558902 220170 558998 220226
rect 558378 220102 558998 220170
rect 558378 220046 558474 220102
rect 558530 220046 558598 220102
rect 558654 220046 558722 220102
rect 558778 220046 558846 220102
rect 558902 220046 558998 220102
rect 558378 219978 558998 220046
rect 558378 219922 558474 219978
rect 558530 219922 558598 219978
rect 558654 219922 558722 219978
rect 558778 219922 558846 219978
rect 558902 219922 558998 219978
rect 558378 202350 558998 219922
rect 558378 202294 558474 202350
rect 558530 202294 558598 202350
rect 558654 202294 558722 202350
rect 558778 202294 558846 202350
rect 558902 202294 558998 202350
rect 558378 202226 558998 202294
rect 558378 202170 558474 202226
rect 558530 202170 558598 202226
rect 558654 202170 558722 202226
rect 558778 202170 558846 202226
rect 558902 202170 558998 202226
rect 558378 202102 558998 202170
rect 558378 202046 558474 202102
rect 558530 202046 558598 202102
rect 558654 202046 558722 202102
rect 558778 202046 558846 202102
rect 558902 202046 558998 202102
rect 558378 201978 558998 202046
rect 558378 201922 558474 201978
rect 558530 201922 558598 201978
rect 558654 201922 558722 201978
rect 558778 201922 558846 201978
rect 558902 201922 558998 201978
rect 558378 184350 558998 201922
rect 558378 184294 558474 184350
rect 558530 184294 558598 184350
rect 558654 184294 558722 184350
rect 558778 184294 558846 184350
rect 558902 184294 558998 184350
rect 558378 184226 558998 184294
rect 558378 184170 558474 184226
rect 558530 184170 558598 184226
rect 558654 184170 558722 184226
rect 558778 184170 558846 184226
rect 558902 184170 558998 184226
rect 558378 184102 558998 184170
rect 558378 184046 558474 184102
rect 558530 184046 558598 184102
rect 558654 184046 558722 184102
rect 558778 184046 558846 184102
rect 558902 184046 558998 184102
rect 558378 183978 558998 184046
rect 558378 183922 558474 183978
rect 558530 183922 558598 183978
rect 558654 183922 558722 183978
rect 558778 183922 558846 183978
rect 558902 183922 558998 183978
rect 558378 166350 558998 183922
rect 558378 166294 558474 166350
rect 558530 166294 558598 166350
rect 558654 166294 558722 166350
rect 558778 166294 558846 166350
rect 558902 166294 558998 166350
rect 558378 166226 558998 166294
rect 558378 166170 558474 166226
rect 558530 166170 558598 166226
rect 558654 166170 558722 166226
rect 558778 166170 558846 166226
rect 558902 166170 558998 166226
rect 558378 166102 558998 166170
rect 558378 166046 558474 166102
rect 558530 166046 558598 166102
rect 558654 166046 558722 166102
rect 558778 166046 558846 166102
rect 558902 166046 558998 166102
rect 558378 165978 558998 166046
rect 558378 165922 558474 165978
rect 558530 165922 558598 165978
rect 558654 165922 558722 165978
rect 558778 165922 558846 165978
rect 558902 165922 558998 165978
rect 558378 149870 558998 165922
rect 559468 343252 559524 343262
rect 556892 147970 556948 147980
rect 479808 136350 480128 136384
rect 479808 136294 479878 136350
rect 479934 136294 480002 136350
rect 480058 136294 480128 136350
rect 479808 136226 480128 136294
rect 479808 136170 479878 136226
rect 479934 136170 480002 136226
rect 480058 136170 480128 136226
rect 479808 136102 480128 136170
rect 479808 136046 479878 136102
rect 479934 136046 480002 136102
rect 480058 136046 480128 136102
rect 479808 135978 480128 136046
rect 479808 135922 479878 135978
rect 479934 135922 480002 135978
rect 480058 135922 480128 135978
rect 479808 135888 480128 135922
rect 510528 136350 510848 136384
rect 510528 136294 510598 136350
rect 510654 136294 510722 136350
rect 510778 136294 510848 136350
rect 510528 136226 510848 136294
rect 510528 136170 510598 136226
rect 510654 136170 510722 136226
rect 510778 136170 510848 136226
rect 510528 136102 510848 136170
rect 510528 136046 510598 136102
rect 510654 136046 510722 136102
rect 510778 136046 510848 136102
rect 510528 135978 510848 136046
rect 510528 135922 510598 135978
rect 510654 135922 510722 135978
rect 510778 135922 510848 135978
rect 510528 135888 510848 135922
rect 541248 136350 541568 136384
rect 541248 136294 541318 136350
rect 541374 136294 541442 136350
rect 541498 136294 541568 136350
rect 541248 136226 541568 136294
rect 541248 136170 541318 136226
rect 541374 136170 541442 136226
rect 541498 136170 541568 136226
rect 541248 136102 541568 136170
rect 541248 136046 541318 136102
rect 541374 136046 541442 136102
rect 541498 136046 541568 136102
rect 541248 135978 541568 136046
rect 541248 135922 541318 135978
rect 541374 135922 541442 135978
rect 541498 135922 541568 135978
rect 541248 135888 541568 135922
rect 464448 130350 464768 130384
rect 464448 130294 464518 130350
rect 464574 130294 464642 130350
rect 464698 130294 464768 130350
rect 464448 130226 464768 130294
rect 464448 130170 464518 130226
rect 464574 130170 464642 130226
rect 464698 130170 464768 130226
rect 464448 130102 464768 130170
rect 464448 130046 464518 130102
rect 464574 130046 464642 130102
rect 464698 130046 464768 130102
rect 464448 129978 464768 130046
rect 464448 129922 464518 129978
rect 464574 129922 464642 129978
rect 464698 129922 464768 129978
rect 464448 129888 464768 129922
rect 495168 130350 495488 130384
rect 495168 130294 495238 130350
rect 495294 130294 495362 130350
rect 495418 130294 495488 130350
rect 495168 130226 495488 130294
rect 495168 130170 495238 130226
rect 495294 130170 495362 130226
rect 495418 130170 495488 130226
rect 495168 130102 495488 130170
rect 495168 130046 495238 130102
rect 495294 130046 495362 130102
rect 495418 130046 495488 130102
rect 495168 129978 495488 130046
rect 495168 129922 495238 129978
rect 495294 129922 495362 129978
rect 495418 129922 495488 129978
rect 495168 129888 495488 129922
rect 525888 130350 526208 130384
rect 525888 130294 525958 130350
rect 526014 130294 526082 130350
rect 526138 130294 526208 130350
rect 525888 130226 526208 130294
rect 525888 130170 525958 130226
rect 526014 130170 526082 130226
rect 526138 130170 526208 130226
rect 525888 130102 526208 130170
rect 525888 130046 525958 130102
rect 526014 130046 526082 130102
rect 526138 130046 526208 130102
rect 525888 129978 526208 130046
rect 525888 129922 525958 129978
rect 526014 129922 526082 129978
rect 526138 129922 526208 129978
rect 525888 129888 526208 129922
rect 556608 130350 556928 130384
rect 556608 130294 556678 130350
rect 556734 130294 556802 130350
rect 556858 130294 556928 130350
rect 556608 130226 556928 130294
rect 556608 130170 556678 130226
rect 556734 130170 556802 130226
rect 556858 130170 556928 130226
rect 556608 130102 556928 130170
rect 556608 130046 556678 130102
rect 556734 130046 556802 130102
rect 556858 130046 556928 130102
rect 556608 129978 556928 130046
rect 556608 129922 556678 129978
rect 556734 129922 556802 129978
rect 556858 129922 556928 129978
rect 556608 129888 556928 129922
rect 457884 128548 457940 128558
rect 457884 83972 457940 128492
rect 457884 83906 457940 83916
rect 457996 120148 458052 120158
rect 457996 81060 458052 120092
rect 479808 118350 480128 118384
rect 479808 118294 479878 118350
rect 479934 118294 480002 118350
rect 480058 118294 480128 118350
rect 479808 118226 480128 118294
rect 479808 118170 479878 118226
rect 479934 118170 480002 118226
rect 480058 118170 480128 118226
rect 479808 118102 480128 118170
rect 479808 118046 479878 118102
rect 479934 118046 480002 118102
rect 480058 118046 480128 118102
rect 479808 117978 480128 118046
rect 479808 117922 479878 117978
rect 479934 117922 480002 117978
rect 480058 117922 480128 117978
rect 479808 117888 480128 117922
rect 510528 118350 510848 118384
rect 510528 118294 510598 118350
rect 510654 118294 510722 118350
rect 510778 118294 510848 118350
rect 510528 118226 510848 118294
rect 510528 118170 510598 118226
rect 510654 118170 510722 118226
rect 510778 118170 510848 118226
rect 510528 118102 510848 118170
rect 510528 118046 510598 118102
rect 510654 118046 510722 118102
rect 510778 118046 510848 118102
rect 510528 117978 510848 118046
rect 510528 117922 510598 117978
rect 510654 117922 510722 117978
rect 510778 117922 510848 117978
rect 510528 117888 510848 117922
rect 541248 118350 541568 118384
rect 541248 118294 541318 118350
rect 541374 118294 541442 118350
rect 541498 118294 541568 118350
rect 541248 118226 541568 118294
rect 541248 118170 541318 118226
rect 541374 118170 541442 118226
rect 541498 118170 541568 118226
rect 541248 118102 541568 118170
rect 541248 118046 541318 118102
rect 541374 118046 541442 118102
rect 541498 118046 541568 118102
rect 541248 117978 541568 118046
rect 541248 117922 541318 117978
rect 541374 117922 541442 117978
rect 541498 117922 541568 117978
rect 541248 117888 541568 117922
rect 464448 112350 464768 112384
rect 464448 112294 464518 112350
rect 464574 112294 464642 112350
rect 464698 112294 464768 112350
rect 464448 112226 464768 112294
rect 464448 112170 464518 112226
rect 464574 112170 464642 112226
rect 464698 112170 464768 112226
rect 464448 112102 464768 112170
rect 464448 112046 464518 112102
rect 464574 112046 464642 112102
rect 464698 112046 464768 112102
rect 464448 111978 464768 112046
rect 464448 111922 464518 111978
rect 464574 111922 464642 111978
rect 464698 111922 464768 111978
rect 464448 111888 464768 111922
rect 495168 112350 495488 112384
rect 495168 112294 495238 112350
rect 495294 112294 495362 112350
rect 495418 112294 495488 112350
rect 495168 112226 495488 112294
rect 495168 112170 495238 112226
rect 495294 112170 495362 112226
rect 495418 112170 495488 112226
rect 495168 112102 495488 112170
rect 495168 112046 495238 112102
rect 495294 112046 495362 112102
rect 495418 112046 495488 112102
rect 495168 111978 495488 112046
rect 495168 111922 495238 111978
rect 495294 111922 495362 111978
rect 495418 111922 495488 111978
rect 495168 111888 495488 111922
rect 525888 112350 526208 112384
rect 525888 112294 525958 112350
rect 526014 112294 526082 112350
rect 526138 112294 526208 112350
rect 525888 112226 526208 112294
rect 525888 112170 525958 112226
rect 526014 112170 526082 112226
rect 526138 112170 526208 112226
rect 525888 112102 526208 112170
rect 525888 112046 525958 112102
rect 526014 112046 526082 112102
rect 526138 112046 526208 112102
rect 525888 111978 526208 112046
rect 525888 111922 525958 111978
rect 526014 111922 526082 111978
rect 526138 111922 526208 111978
rect 525888 111888 526208 111922
rect 556608 112350 556928 112384
rect 556608 112294 556678 112350
rect 556734 112294 556802 112350
rect 556858 112294 556928 112350
rect 556608 112226 556928 112294
rect 556608 112170 556678 112226
rect 556734 112170 556802 112226
rect 556858 112170 556928 112226
rect 556608 112102 556928 112170
rect 556608 112046 556678 112102
rect 556734 112046 556802 112102
rect 556858 112046 556928 112102
rect 556608 111978 556928 112046
rect 556608 111922 556678 111978
rect 556734 111922 556802 111978
rect 556858 111922 556928 111978
rect 556608 111888 556928 111922
rect 479808 100350 480128 100384
rect 479808 100294 479878 100350
rect 479934 100294 480002 100350
rect 480058 100294 480128 100350
rect 479808 100226 480128 100294
rect 479808 100170 479878 100226
rect 479934 100170 480002 100226
rect 480058 100170 480128 100226
rect 479808 100102 480128 100170
rect 479808 100046 479878 100102
rect 479934 100046 480002 100102
rect 480058 100046 480128 100102
rect 479808 99978 480128 100046
rect 479808 99922 479878 99978
rect 479934 99922 480002 99978
rect 480058 99922 480128 99978
rect 479808 99888 480128 99922
rect 510528 100350 510848 100384
rect 510528 100294 510598 100350
rect 510654 100294 510722 100350
rect 510778 100294 510848 100350
rect 510528 100226 510848 100294
rect 510528 100170 510598 100226
rect 510654 100170 510722 100226
rect 510778 100170 510848 100226
rect 510528 100102 510848 100170
rect 510528 100046 510598 100102
rect 510654 100046 510722 100102
rect 510778 100046 510848 100102
rect 510528 99978 510848 100046
rect 510528 99922 510598 99978
rect 510654 99922 510722 99978
rect 510778 99922 510848 99978
rect 510528 99888 510848 99922
rect 541248 100350 541568 100384
rect 541248 100294 541318 100350
rect 541374 100294 541442 100350
rect 541498 100294 541568 100350
rect 541248 100226 541568 100294
rect 541248 100170 541318 100226
rect 541374 100170 541442 100226
rect 541498 100170 541568 100226
rect 541248 100102 541568 100170
rect 541248 100046 541318 100102
rect 541374 100046 541442 100102
rect 541498 100046 541568 100102
rect 541248 99978 541568 100046
rect 541248 99922 541318 99978
rect 541374 99922 541442 99978
rect 541498 99922 541568 99978
rect 541248 99888 541568 99922
rect 464448 94350 464768 94384
rect 464448 94294 464518 94350
rect 464574 94294 464642 94350
rect 464698 94294 464768 94350
rect 464448 94226 464768 94294
rect 464448 94170 464518 94226
rect 464574 94170 464642 94226
rect 464698 94170 464768 94226
rect 464448 94102 464768 94170
rect 464448 94046 464518 94102
rect 464574 94046 464642 94102
rect 464698 94046 464768 94102
rect 464448 93978 464768 94046
rect 464448 93922 464518 93978
rect 464574 93922 464642 93978
rect 464698 93922 464768 93978
rect 464448 93888 464768 93922
rect 495168 94350 495488 94384
rect 495168 94294 495238 94350
rect 495294 94294 495362 94350
rect 495418 94294 495488 94350
rect 495168 94226 495488 94294
rect 495168 94170 495238 94226
rect 495294 94170 495362 94226
rect 495418 94170 495488 94226
rect 495168 94102 495488 94170
rect 495168 94046 495238 94102
rect 495294 94046 495362 94102
rect 495418 94046 495488 94102
rect 495168 93978 495488 94046
rect 495168 93922 495238 93978
rect 495294 93922 495362 93978
rect 495418 93922 495488 93978
rect 495168 93888 495488 93922
rect 525888 94350 526208 94384
rect 525888 94294 525958 94350
rect 526014 94294 526082 94350
rect 526138 94294 526208 94350
rect 525888 94226 526208 94294
rect 525888 94170 525958 94226
rect 526014 94170 526082 94226
rect 526138 94170 526208 94226
rect 525888 94102 526208 94170
rect 525888 94046 525958 94102
rect 526014 94046 526082 94102
rect 526138 94046 526208 94102
rect 525888 93978 526208 94046
rect 525888 93922 525958 93978
rect 526014 93922 526082 93978
rect 526138 93922 526208 93978
rect 525888 93888 526208 93922
rect 556608 94350 556928 94384
rect 556608 94294 556678 94350
rect 556734 94294 556802 94350
rect 556858 94294 556928 94350
rect 556608 94226 556928 94294
rect 556608 94170 556678 94226
rect 556734 94170 556802 94226
rect 556858 94170 556928 94226
rect 556608 94102 556928 94170
rect 556608 94046 556678 94102
rect 556734 94046 556802 94102
rect 556858 94046 556928 94102
rect 556608 93978 556928 94046
rect 556608 93922 556678 93978
rect 556734 93922 556802 93978
rect 556858 93922 556928 93978
rect 556608 93888 556928 93922
rect 479808 82350 480128 82384
rect 479808 82294 479878 82350
rect 479934 82294 480002 82350
rect 480058 82294 480128 82350
rect 479808 82226 480128 82294
rect 479808 82170 479878 82226
rect 479934 82170 480002 82226
rect 480058 82170 480128 82226
rect 479808 82102 480128 82170
rect 479808 82046 479878 82102
rect 479934 82046 480002 82102
rect 480058 82046 480128 82102
rect 479808 81978 480128 82046
rect 479808 81922 479878 81978
rect 479934 81922 480002 81978
rect 480058 81922 480128 81978
rect 479808 81888 480128 81922
rect 510528 82350 510848 82384
rect 510528 82294 510598 82350
rect 510654 82294 510722 82350
rect 510778 82294 510848 82350
rect 510528 82226 510848 82294
rect 510528 82170 510598 82226
rect 510654 82170 510722 82226
rect 510778 82170 510848 82226
rect 510528 82102 510848 82170
rect 510528 82046 510598 82102
rect 510654 82046 510722 82102
rect 510778 82046 510848 82102
rect 510528 81978 510848 82046
rect 510528 81922 510598 81978
rect 510654 81922 510722 81978
rect 510778 81922 510848 81978
rect 510528 81888 510848 81922
rect 541248 82350 541568 82384
rect 541248 82294 541318 82350
rect 541374 82294 541442 82350
rect 541498 82294 541568 82350
rect 541248 82226 541568 82294
rect 541248 82170 541318 82226
rect 541374 82170 541442 82226
rect 541498 82170 541568 82226
rect 541248 82102 541568 82170
rect 541248 82046 541318 82102
rect 541374 82046 541442 82102
rect 541498 82046 541568 82102
rect 541248 81978 541568 82046
rect 541248 81922 541318 81978
rect 541374 81922 541442 81978
rect 541498 81922 541568 81978
rect 541248 81888 541568 81922
rect 457996 80994 458052 81004
rect 464448 76350 464768 76384
rect 464448 76294 464518 76350
rect 464574 76294 464642 76350
rect 464698 76294 464768 76350
rect 464448 76226 464768 76294
rect 464448 76170 464518 76226
rect 464574 76170 464642 76226
rect 464698 76170 464768 76226
rect 464448 76102 464768 76170
rect 464448 76046 464518 76102
rect 464574 76046 464642 76102
rect 464698 76046 464768 76102
rect 464448 75978 464768 76046
rect 464448 75922 464518 75978
rect 464574 75922 464642 75978
rect 464698 75922 464768 75978
rect 464448 75888 464768 75922
rect 495168 76350 495488 76384
rect 495168 76294 495238 76350
rect 495294 76294 495362 76350
rect 495418 76294 495488 76350
rect 495168 76226 495488 76294
rect 495168 76170 495238 76226
rect 495294 76170 495362 76226
rect 495418 76170 495488 76226
rect 495168 76102 495488 76170
rect 495168 76046 495238 76102
rect 495294 76046 495362 76102
rect 495418 76046 495488 76102
rect 495168 75978 495488 76046
rect 495168 75922 495238 75978
rect 495294 75922 495362 75978
rect 495418 75922 495488 75978
rect 495168 75888 495488 75922
rect 525888 76350 526208 76384
rect 525888 76294 525958 76350
rect 526014 76294 526082 76350
rect 526138 76294 526208 76350
rect 525888 76226 526208 76294
rect 525888 76170 525958 76226
rect 526014 76170 526082 76226
rect 526138 76170 526208 76226
rect 525888 76102 526208 76170
rect 525888 76046 525958 76102
rect 526014 76046 526082 76102
rect 526138 76046 526208 76102
rect 525888 75978 526208 76046
rect 525888 75922 525958 75978
rect 526014 75922 526082 75978
rect 526138 75922 526208 75978
rect 525888 75888 526208 75922
rect 556608 76350 556928 76384
rect 556608 76294 556678 76350
rect 556734 76294 556802 76350
rect 556858 76294 556928 76350
rect 556608 76226 556928 76294
rect 556608 76170 556678 76226
rect 556734 76170 556802 76226
rect 556858 76170 556928 76226
rect 556608 76102 556928 76170
rect 556608 76046 556678 76102
rect 556734 76046 556802 76102
rect 556858 76046 556928 76102
rect 556608 75978 556928 76046
rect 556608 75922 556678 75978
rect 556734 75922 556802 75978
rect 556858 75922 556928 75978
rect 556608 75888 556928 75922
rect 559468 67732 559524 343196
rect 559580 70868 559636 345436
rect 560252 120932 560308 371196
rect 560252 120866 560308 120876
rect 562098 370350 562718 387922
rect 562098 370294 562194 370350
rect 562250 370294 562318 370350
rect 562374 370294 562442 370350
rect 562498 370294 562566 370350
rect 562622 370294 562718 370350
rect 562098 370226 562718 370294
rect 562098 370170 562194 370226
rect 562250 370170 562318 370226
rect 562374 370170 562442 370226
rect 562498 370170 562566 370226
rect 562622 370170 562718 370226
rect 562098 370102 562718 370170
rect 562098 370046 562194 370102
rect 562250 370046 562318 370102
rect 562374 370046 562442 370102
rect 562498 370046 562566 370102
rect 562622 370046 562718 370102
rect 562098 369978 562718 370046
rect 562098 369922 562194 369978
rect 562250 369922 562318 369978
rect 562374 369922 562442 369978
rect 562498 369922 562566 369978
rect 562622 369922 562718 369978
rect 562098 352350 562718 369922
rect 577052 389818 577108 389828
rect 573132 369012 573188 369022
rect 571564 368788 571620 368798
rect 568204 366772 568260 366782
rect 564956 362068 565012 362078
rect 562098 352294 562194 352350
rect 562250 352294 562318 352350
rect 562374 352294 562442 352350
rect 562498 352294 562566 352350
rect 562622 352294 562718 352350
rect 562098 352226 562718 352294
rect 562098 352170 562194 352226
rect 562250 352170 562318 352226
rect 562374 352170 562442 352226
rect 562498 352170 562566 352226
rect 562622 352170 562718 352226
rect 562098 352102 562718 352170
rect 562098 352046 562194 352102
rect 562250 352046 562318 352102
rect 562374 352046 562442 352102
rect 562498 352046 562566 352102
rect 562622 352046 562718 352102
rect 562098 351978 562718 352046
rect 562098 351922 562194 351978
rect 562250 351922 562318 351978
rect 562374 351922 562442 351978
rect 562498 351922 562566 351978
rect 562622 351922 562718 351978
rect 562098 334350 562718 351922
rect 564844 353332 564900 353342
rect 564732 348852 564788 348862
rect 564620 346612 564676 346622
rect 562098 334294 562194 334350
rect 562250 334294 562318 334350
rect 562374 334294 562442 334350
rect 562498 334294 562566 334350
rect 562622 334294 562718 334350
rect 562098 334226 562718 334294
rect 562098 334170 562194 334226
rect 562250 334170 562318 334226
rect 562374 334170 562442 334226
rect 562498 334170 562566 334226
rect 562622 334170 562718 334226
rect 562098 334102 562718 334170
rect 562098 334046 562194 334102
rect 562250 334046 562318 334102
rect 562374 334046 562442 334102
rect 562498 334046 562566 334102
rect 562622 334046 562718 334102
rect 562098 333978 562718 334046
rect 562098 333922 562194 333978
rect 562250 333922 562318 333978
rect 562374 333922 562442 333978
rect 562498 333922 562566 333978
rect 562622 333922 562718 333978
rect 562098 316350 562718 333922
rect 564508 335412 564564 335422
rect 562098 316294 562194 316350
rect 562250 316294 562318 316350
rect 562374 316294 562442 316350
rect 562498 316294 562566 316350
rect 562622 316294 562718 316350
rect 562098 316226 562718 316294
rect 562098 316170 562194 316226
rect 562250 316170 562318 316226
rect 562374 316170 562442 316226
rect 562498 316170 562566 316226
rect 562622 316170 562718 316226
rect 562098 316102 562718 316170
rect 562098 316046 562194 316102
rect 562250 316046 562318 316102
rect 562374 316046 562442 316102
rect 562498 316046 562566 316102
rect 562622 316046 562718 316102
rect 562098 315978 562718 316046
rect 562098 315922 562194 315978
rect 562250 315922 562318 315978
rect 562374 315922 562442 315978
rect 562498 315922 562566 315978
rect 562622 315922 562718 315978
rect 562098 298350 562718 315922
rect 562098 298294 562194 298350
rect 562250 298294 562318 298350
rect 562374 298294 562442 298350
rect 562498 298294 562566 298350
rect 562622 298294 562718 298350
rect 562098 298226 562718 298294
rect 562098 298170 562194 298226
rect 562250 298170 562318 298226
rect 562374 298170 562442 298226
rect 562498 298170 562566 298226
rect 562622 298170 562718 298226
rect 562098 298102 562718 298170
rect 562098 298046 562194 298102
rect 562250 298046 562318 298102
rect 562374 298046 562442 298102
rect 562498 298046 562566 298102
rect 562622 298046 562718 298102
rect 562098 297978 562718 298046
rect 562098 297922 562194 297978
rect 562250 297922 562318 297978
rect 562374 297922 562442 297978
rect 562498 297922 562566 297978
rect 562622 297922 562718 297978
rect 562098 280350 562718 297922
rect 562098 280294 562194 280350
rect 562250 280294 562318 280350
rect 562374 280294 562442 280350
rect 562498 280294 562566 280350
rect 562622 280294 562718 280350
rect 562098 280226 562718 280294
rect 562098 280170 562194 280226
rect 562250 280170 562318 280226
rect 562374 280170 562442 280226
rect 562498 280170 562566 280226
rect 562622 280170 562718 280226
rect 562098 280102 562718 280170
rect 562098 280046 562194 280102
rect 562250 280046 562318 280102
rect 562374 280046 562442 280102
rect 562498 280046 562566 280102
rect 562622 280046 562718 280102
rect 562098 279978 562718 280046
rect 562098 279922 562194 279978
rect 562250 279922 562318 279978
rect 562374 279922 562442 279978
rect 562498 279922 562566 279978
rect 562622 279922 562718 279978
rect 562098 262350 562718 279922
rect 562098 262294 562194 262350
rect 562250 262294 562318 262350
rect 562374 262294 562442 262350
rect 562498 262294 562566 262350
rect 562622 262294 562718 262350
rect 562098 262226 562718 262294
rect 562098 262170 562194 262226
rect 562250 262170 562318 262226
rect 562374 262170 562442 262226
rect 562498 262170 562566 262226
rect 562622 262170 562718 262226
rect 562098 262102 562718 262170
rect 562098 262046 562194 262102
rect 562250 262046 562318 262102
rect 562374 262046 562442 262102
rect 562498 262046 562566 262102
rect 562622 262046 562718 262102
rect 562098 261978 562718 262046
rect 562098 261922 562194 261978
rect 562250 261922 562318 261978
rect 562374 261922 562442 261978
rect 562498 261922 562566 261978
rect 562622 261922 562718 261978
rect 562098 244350 562718 261922
rect 562098 244294 562194 244350
rect 562250 244294 562318 244350
rect 562374 244294 562442 244350
rect 562498 244294 562566 244350
rect 562622 244294 562718 244350
rect 562098 244226 562718 244294
rect 562098 244170 562194 244226
rect 562250 244170 562318 244226
rect 562374 244170 562442 244226
rect 562498 244170 562566 244226
rect 562622 244170 562718 244226
rect 562098 244102 562718 244170
rect 562098 244046 562194 244102
rect 562250 244046 562318 244102
rect 562374 244046 562442 244102
rect 562498 244046 562566 244102
rect 562622 244046 562718 244102
rect 562098 243978 562718 244046
rect 562098 243922 562194 243978
rect 562250 243922 562318 243978
rect 562374 243922 562442 243978
rect 562498 243922 562566 243978
rect 562622 243922 562718 243978
rect 562098 226350 562718 243922
rect 562098 226294 562194 226350
rect 562250 226294 562318 226350
rect 562374 226294 562442 226350
rect 562498 226294 562566 226350
rect 562622 226294 562718 226350
rect 562098 226226 562718 226294
rect 562098 226170 562194 226226
rect 562250 226170 562318 226226
rect 562374 226170 562442 226226
rect 562498 226170 562566 226226
rect 562622 226170 562718 226226
rect 562098 226102 562718 226170
rect 562098 226046 562194 226102
rect 562250 226046 562318 226102
rect 562374 226046 562442 226102
rect 562498 226046 562566 226102
rect 562622 226046 562718 226102
rect 562098 225978 562718 226046
rect 562098 225922 562194 225978
rect 562250 225922 562318 225978
rect 562374 225922 562442 225978
rect 562498 225922 562566 225978
rect 562622 225922 562718 225978
rect 562098 208350 562718 225922
rect 562098 208294 562194 208350
rect 562250 208294 562318 208350
rect 562374 208294 562442 208350
rect 562498 208294 562566 208350
rect 562622 208294 562718 208350
rect 562098 208226 562718 208294
rect 562098 208170 562194 208226
rect 562250 208170 562318 208226
rect 562374 208170 562442 208226
rect 562498 208170 562566 208226
rect 562622 208170 562718 208226
rect 562098 208102 562718 208170
rect 562098 208046 562194 208102
rect 562250 208046 562318 208102
rect 562374 208046 562442 208102
rect 562498 208046 562566 208102
rect 562622 208046 562718 208102
rect 562098 207978 562718 208046
rect 562098 207922 562194 207978
rect 562250 207922 562318 207978
rect 562374 207922 562442 207978
rect 562498 207922 562566 207978
rect 562622 207922 562718 207978
rect 562098 190350 562718 207922
rect 562098 190294 562194 190350
rect 562250 190294 562318 190350
rect 562374 190294 562442 190350
rect 562498 190294 562566 190350
rect 562622 190294 562718 190350
rect 562098 190226 562718 190294
rect 562098 190170 562194 190226
rect 562250 190170 562318 190226
rect 562374 190170 562442 190226
rect 562498 190170 562566 190226
rect 562622 190170 562718 190226
rect 562098 190102 562718 190170
rect 562098 190046 562194 190102
rect 562250 190046 562318 190102
rect 562374 190046 562442 190102
rect 562498 190046 562566 190102
rect 562622 190046 562718 190102
rect 562098 189978 562718 190046
rect 562098 189922 562194 189978
rect 562250 189922 562318 189978
rect 562374 189922 562442 189978
rect 562498 189922 562566 189978
rect 562622 189922 562718 189978
rect 562098 172350 562718 189922
rect 562098 172294 562194 172350
rect 562250 172294 562318 172350
rect 562374 172294 562442 172350
rect 562498 172294 562566 172350
rect 562622 172294 562718 172350
rect 562098 172226 562718 172294
rect 562098 172170 562194 172226
rect 562250 172170 562318 172226
rect 562374 172170 562442 172226
rect 562498 172170 562566 172226
rect 562622 172170 562718 172226
rect 562098 172102 562718 172170
rect 562098 172046 562194 172102
rect 562250 172046 562318 172102
rect 562374 172046 562442 172102
rect 562498 172046 562566 172102
rect 562622 172046 562718 172102
rect 562098 171978 562718 172046
rect 562098 171922 562194 171978
rect 562250 171922 562318 171978
rect 562374 171922 562442 171978
rect 562498 171922 562566 171978
rect 562622 171922 562718 171978
rect 562098 154350 562718 171922
rect 562098 154294 562194 154350
rect 562250 154294 562318 154350
rect 562374 154294 562442 154350
rect 562498 154294 562566 154350
rect 562622 154294 562718 154350
rect 562098 154226 562718 154294
rect 562098 154170 562194 154226
rect 562250 154170 562318 154226
rect 562374 154170 562442 154226
rect 562498 154170 562566 154226
rect 562622 154170 562718 154226
rect 562098 154102 562718 154170
rect 562098 154046 562194 154102
rect 562250 154046 562318 154102
rect 562374 154046 562442 154102
rect 562498 154046 562566 154102
rect 562622 154046 562718 154102
rect 562098 153978 562718 154046
rect 562098 153922 562194 153978
rect 562250 153922 562318 153978
rect 562374 153922 562442 153978
rect 562498 153922 562566 153978
rect 562622 153922 562718 153978
rect 562098 136350 562718 153922
rect 563276 331828 563332 331838
rect 563164 148708 563220 148718
rect 563052 148148 563108 148158
rect 562098 136294 562194 136350
rect 562250 136294 562318 136350
rect 562374 136294 562442 136350
rect 562498 136294 562566 136350
rect 562622 136294 562718 136350
rect 562098 136226 562718 136294
rect 562098 136170 562194 136226
rect 562250 136170 562318 136226
rect 562374 136170 562442 136226
rect 562498 136170 562566 136226
rect 562622 136170 562718 136226
rect 562098 136102 562718 136170
rect 562098 136046 562194 136102
rect 562250 136046 562318 136102
rect 562374 136046 562442 136102
rect 562498 136046 562566 136102
rect 562622 136046 562718 136102
rect 562098 135978 562718 136046
rect 562098 135922 562194 135978
rect 562250 135922 562318 135978
rect 562374 135922 562442 135978
rect 562498 135922 562566 135978
rect 562622 135922 562718 135978
rect 559580 70802 559636 70812
rect 562098 118350 562718 135922
rect 562940 148036 562996 148046
rect 562098 118294 562194 118350
rect 562250 118294 562318 118350
rect 562374 118294 562442 118350
rect 562498 118294 562566 118350
rect 562622 118294 562718 118350
rect 562098 118226 562718 118294
rect 562098 118170 562194 118226
rect 562250 118170 562318 118226
rect 562374 118170 562442 118226
rect 562498 118170 562566 118226
rect 562622 118170 562718 118226
rect 562098 118102 562718 118170
rect 562098 118046 562194 118102
rect 562250 118046 562318 118102
rect 562374 118046 562442 118102
rect 562498 118046 562566 118102
rect 562622 118046 562718 118102
rect 562098 117978 562718 118046
rect 562098 117922 562194 117978
rect 562250 117922 562318 117978
rect 562374 117922 562442 117978
rect 562498 117922 562566 117978
rect 562622 117922 562718 117978
rect 562098 100350 562718 117922
rect 562828 120932 562884 120942
rect 562828 106932 562884 120876
rect 562828 106866 562884 106876
rect 562098 100294 562194 100350
rect 562250 100294 562318 100350
rect 562374 100294 562442 100350
rect 562498 100294 562566 100350
rect 562622 100294 562718 100350
rect 562098 100226 562718 100294
rect 562098 100170 562194 100226
rect 562250 100170 562318 100226
rect 562374 100170 562442 100226
rect 562498 100170 562566 100226
rect 562622 100170 562718 100226
rect 562098 100102 562718 100170
rect 562098 100046 562194 100102
rect 562250 100046 562318 100102
rect 562374 100046 562442 100102
rect 562498 100046 562566 100102
rect 562622 100046 562718 100102
rect 562098 99978 562718 100046
rect 562098 99922 562194 99978
rect 562250 99922 562318 99978
rect 562374 99922 562442 99978
rect 562498 99922 562566 99978
rect 562622 99922 562718 99978
rect 562098 82350 562718 99922
rect 562098 82294 562194 82350
rect 562250 82294 562318 82350
rect 562374 82294 562442 82350
rect 562498 82294 562566 82350
rect 562622 82294 562718 82350
rect 562098 82226 562718 82294
rect 562098 82170 562194 82226
rect 562250 82170 562318 82226
rect 562374 82170 562442 82226
rect 562498 82170 562566 82226
rect 562622 82170 562718 82226
rect 562098 82102 562718 82170
rect 562098 82046 562194 82102
rect 562250 82046 562318 82102
rect 562374 82046 562442 82102
rect 562498 82046 562566 82102
rect 562622 82046 562718 82102
rect 562098 81978 562718 82046
rect 562098 81922 562194 81978
rect 562250 81922 562318 81978
rect 562374 81922 562442 81978
rect 562498 81922 562566 81978
rect 562622 81922 562718 81978
rect 559468 67666 559524 67676
rect 479808 64350 480128 64384
rect 479808 64294 479878 64350
rect 479934 64294 480002 64350
rect 480058 64294 480128 64350
rect 479808 64226 480128 64294
rect 479808 64170 479878 64226
rect 479934 64170 480002 64226
rect 480058 64170 480128 64226
rect 479808 64102 480128 64170
rect 479808 64046 479878 64102
rect 479934 64046 480002 64102
rect 480058 64046 480128 64102
rect 479808 63978 480128 64046
rect 479808 63922 479878 63978
rect 479934 63922 480002 63978
rect 480058 63922 480128 63978
rect 479808 63888 480128 63922
rect 510528 64350 510848 64384
rect 510528 64294 510598 64350
rect 510654 64294 510722 64350
rect 510778 64294 510848 64350
rect 510528 64226 510848 64294
rect 510528 64170 510598 64226
rect 510654 64170 510722 64226
rect 510778 64170 510848 64226
rect 510528 64102 510848 64170
rect 510528 64046 510598 64102
rect 510654 64046 510722 64102
rect 510778 64046 510848 64102
rect 510528 63978 510848 64046
rect 510528 63922 510598 63978
rect 510654 63922 510722 63978
rect 510778 63922 510848 63978
rect 510528 63888 510848 63922
rect 541248 64350 541568 64384
rect 541248 64294 541318 64350
rect 541374 64294 541442 64350
rect 541498 64294 541568 64350
rect 541248 64226 541568 64294
rect 541248 64170 541318 64226
rect 541374 64170 541442 64226
rect 541498 64170 541568 64226
rect 541248 64102 541568 64170
rect 541248 64046 541318 64102
rect 541374 64046 541442 64102
rect 541498 64046 541568 64102
rect 541248 63978 541568 64046
rect 541248 63922 541318 63978
rect 541374 63922 541442 63978
rect 541498 63922 541568 63978
rect 541248 63888 541568 63922
rect 562098 64350 562718 81922
rect 562098 64294 562194 64350
rect 562250 64294 562318 64350
rect 562374 64294 562442 64350
rect 562498 64294 562566 64350
rect 562622 64294 562718 64350
rect 562098 64226 562718 64294
rect 562098 64170 562194 64226
rect 562250 64170 562318 64226
rect 562374 64170 562442 64226
rect 562498 64170 562566 64226
rect 562622 64170 562718 64226
rect 562098 64102 562718 64170
rect 562098 64046 562194 64102
rect 562250 64046 562318 64102
rect 562374 64046 562442 64102
rect 562498 64046 562566 64102
rect 562622 64046 562718 64102
rect 562098 63978 562718 64046
rect 562098 63922 562194 63978
rect 562250 63922 562318 63978
rect 562374 63922 562442 63978
rect 562498 63922 562566 63978
rect 562622 63922 562718 63978
rect 464448 58350 464768 58384
rect 464448 58294 464518 58350
rect 464574 58294 464642 58350
rect 464698 58294 464768 58350
rect 464448 58226 464768 58294
rect 464448 58170 464518 58226
rect 464574 58170 464642 58226
rect 464698 58170 464768 58226
rect 464448 58102 464768 58170
rect 464448 58046 464518 58102
rect 464574 58046 464642 58102
rect 464698 58046 464768 58102
rect 464448 57978 464768 58046
rect 464448 57922 464518 57978
rect 464574 57922 464642 57978
rect 464698 57922 464768 57978
rect 464448 57888 464768 57922
rect 495168 58350 495488 58384
rect 495168 58294 495238 58350
rect 495294 58294 495362 58350
rect 495418 58294 495488 58350
rect 495168 58226 495488 58294
rect 495168 58170 495238 58226
rect 495294 58170 495362 58226
rect 495418 58170 495488 58226
rect 495168 58102 495488 58170
rect 495168 58046 495238 58102
rect 495294 58046 495362 58102
rect 495418 58046 495488 58102
rect 495168 57978 495488 58046
rect 495168 57922 495238 57978
rect 495294 57922 495362 57978
rect 495418 57922 495488 57978
rect 495168 57888 495488 57922
rect 525888 58350 526208 58384
rect 525888 58294 525958 58350
rect 526014 58294 526082 58350
rect 526138 58294 526208 58350
rect 525888 58226 526208 58294
rect 525888 58170 525958 58226
rect 526014 58170 526082 58226
rect 526138 58170 526208 58226
rect 525888 58102 526208 58170
rect 525888 58046 525958 58102
rect 526014 58046 526082 58102
rect 526138 58046 526208 58102
rect 525888 57978 526208 58046
rect 525888 57922 525958 57978
rect 526014 57922 526082 57978
rect 526138 57922 526208 57978
rect 525888 57888 526208 57922
rect 556608 58350 556928 58384
rect 556608 58294 556678 58350
rect 556734 58294 556802 58350
rect 556858 58294 556928 58350
rect 556608 58226 556928 58294
rect 556608 58170 556678 58226
rect 556734 58170 556802 58226
rect 556858 58170 556928 58226
rect 556608 58102 556928 58170
rect 556608 58046 556678 58102
rect 556734 58046 556802 58102
rect 556858 58046 556928 58102
rect 556608 57978 556928 58046
rect 556608 57922 556678 57978
rect 556734 57922 556802 57978
rect 556858 57922 556928 57978
rect 556608 57888 556928 57922
rect 457772 54786 457828 54796
rect 439218 46294 439314 46350
rect 439370 46294 439438 46350
rect 439494 46294 439562 46350
rect 439618 46294 439686 46350
rect 439742 46294 439838 46350
rect 439218 46226 439838 46294
rect 439218 46170 439314 46226
rect 439370 46170 439438 46226
rect 439494 46170 439562 46226
rect 439618 46170 439686 46226
rect 439742 46170 439838 46226
rect 439218 46102 439838 46170
rect 439218 46046 439314 46102
rect 439370 46046 439438 46102
rect 439494 46046 439562 46102
rect 439618 46046 439686 46102
rect 439742 46046 439838 46102
rect 439218 45978 439838 46046
rect 439218 45922 439314 45978
rect 439370 45922 439438 45978
rect 439494 45922 439562 45978
rect 439618 45922 439686 45978
rect 439742 45922 439838 45978
rect 439218 28350 439838 45922
rect 439218 28294 439314 28350
rect 439370 28294 439438 28350
rect 439494 28294 439562 28350
rect 439618 28294 439686 28350
rect 439742 28294 439838 28350
rect 439218 28226 439838 28294
rect 439218 28170 439314 28226
rect 439370 28170 439438 28226
rect 439494 28170 439562 28226
rect 439618 28170 439686 28226
rect 439742 28170 439838 28226
rect 439218 28102 439838 28170
rect 439218 28046 439314 28102
rect 439370 28046 439438 28102
rect 439494 28046 439562 28102
rect 439618 28046 439686 28102
rect 439742 28046 439838 28102
rect 439218 27978 439838 28046
rect 439218 27922 439314 27978
rect 439370 27922 439438 27978
rect 439494 27922 439562 27978
rect 439618 27922 439686 27978
rect 439742 27922 439838 27978
rect 439218 10350 439838 27922
rect 439218 10294 439314 10350
rect 439370 10294 439438 10350
rect 439494 10294 439562 10350
rect 439618 10294 439686 10350
rect 439742 10294 439838 10350
rect 439218 10226 439838 10294
rect 439218 10170 439314 10226
rect 439370 10170 439438 10226
rect 439494 10170 439562 10226
rect 439618 10170 439686 10226
rect 439742 10170 439838 10226
rect 439218 10102 439838 10170
rect 439218 10046 439314 10102
rect 439370 10046 439438 10102
rect 439494 10046 439562 10102
rect 439618 10046 439686 10102
rect 439742 10046 439838 10102
rect 439218 9978 439838 10046
rect 439218 9922 439314 9978
rect 439370 9922 439438 9978
rect 439494 9922 439562 9978
rect 439618 9922 439686 9978
rect 439742 9922 439838 9978
rect 439218 -1120 439838 9922
rect 439218 -1176 439314 -1120
rect 439370 -1176 439438 -1120
rect 439494 -1176 439562 -1120
rect 439618 -1176 439686 -1120
rect 439742 -1176 439838 -1120
rect 439218 -1244 439838 -1176
rect 439218 -1300 439314 -1244
rect 439370 -1300 439438 -1244
rect 439494 -1300 439562 -1244
rect 439618 -1300 439686 -1244
rect 439742 -1300 439838 -1244
rect 439218 -1368 439838 -1300
rect 439218 -1424 439314 -1368
rect 439370 -1424 439438 -1368
rect 439494 -1424 439562 -1368
rect 439618 -1424 439686 -1368
rect 439742 -1424 439838 -1368
rect 439218 -1492 439838 -1424
rect 439218 -1548 439314 -1492
rect 439370 -1548 439438 -1492
rect 439494 -1548 439562 -1492
rect 439618 -1548 439686 -1492
rect 439742 -1548 439838 -1492
rect 439218 -1644 439838 -1548
rect 466218 40350 466838 48690
rect 466218 40294 466314 40350
rect 466370 40294 466438 40350
rect 466494 40294 466562 40350
rect 466618 40294 466686 40350
rect 466742 40294 466838 40350
rect 466218 40226 466838 40294
rect 466218 40170 466314 40226
rect 466370 40170 466438 40226
rect 466494 40170 466562 40226
rect 466618 40170 466686 40226
rect 466742 40170 466838 40226
rect 466218 40102 466838 40170
rect 466218 40046 466314 40102
rect 466370 40046 466438 40102
rect 466494 40046 466562 40102
rect 466618 40046 466686 40102
rect 466742 40046 466838 40102
rect 466218 39978 466838 40046
rect 466218 39922 466314 39978
rect 466370 39922 466438 39978
rect 466494 39922 466562 39978
rect 466618 39922 466686 39978
rect 466742 39922 466838 39978
rect 466218 22350 466838 39922
rect 466218 22294 466314 22350
rect 466370 22294 466438 22350
rect 466494 22294 466562 22350
rect 466618 22294 466686 22350
rect 466742 22294 466838 22350
rect 466218 22226 466838 22294
rect 466218 22170 466314 22226
rect 466370 22170 466438 22226
rect 466494 22170 466562 22226
rect 466618 22170 466686 22226
rect 466742 22170 466838 22226
rect 466218 22102 466838 22170
rect 466218 22046 466314 22102
rect 466370 22046 466438 22102
rect 466494 22046 466562 22102
rect 466618 22046 466686 22102
rect 466742 22046 466838 22102
rect 466218 21978 466838 22046
rect 466218 21922 466314 21978
rect 466370 21922 466438 21978
rect 466494 21922 466562 21978
rect 466618 21922 466686 21978
rect 466742 21922 466838 21978
rect 466218 4350 466838 21922
rect 466218 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 466838 4350
rect 466218 4226 466838 4294
rect 466218 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 466838 4226
rect 466218 4102 466838 4170
rect 466218 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 466838 4102
rect 466218 3978 466838 4046
rect 466218 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 466838 3978
rect 466218 -160 466838 3922
rect 466218 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 466838 -160
rect 466218 -284 466838 -216
rect 466218 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 466838 -284
rect 466218 -408 466838 -340
rect 466218 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 466838 -408
rect 466218 -532 466838 -464
rect 466218 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 466838 -532
rect 466218 -1644 466838 -588
rect 469938 46350 470558 48690
rect 469938 46294 470034 46350
rect 470090 46294 470158 46350
rect 470214 46294 470282 46350
rect 470338 46294 470406 46350
rect 470462 46294 470558 46350
rect 469938 46226 470558 46294
rect 469938 46170 470034 46226
rect 470090 46170 470158 46226
rect 470214 46170 470282 46226
rect 470338 46170 470406 46226
rect 470462 46170 470558 46226
rect 469938 46102 470558 46170
rect 469938 46046 470034 46102
rect 470090 46046 470158 46102
rect 470214 46046 470282 46102
rect 470338 46046 470406 46102
rect 470462 46046 470558 46102
rect 469938 45978 470558 46046
rect 469938 45922 470034 45978
rect 470090 45922 470158 45978
rect 470214 45922 470282 45978
rect 470338 45922 470406 45978
rect 470462 45922 470558 45978
rect 469938 28350 470558 45922
rect 469938 28294 470034 28350
rect 470090 28294 470158 28350
rect 470214 28294 470282 28350
rect 470338 28294 470406 28350
rect 470462 28294 470558 28350
rect 469938 28226 470558 28294
rect 469938 28170 470034 28226
rect 470090 28170 470158 28226
rect 470214 28170 470282 28226
rect 470338 28170 470406 28226
rect 470462 28170 470558 28226
rect 469938 28102 470558 28170
rect 469938 28046 470034 28102
rect 470090 28046 470158 28102
rect 470214 28046 470282 28102
rect 470338 28046 470406 28102
rect 470462 28046 470558 28102
rect 469938 27978 470558 28046
rect 469938 27922 470034 27978
rect 470090 27922 470158 27978
rect 470214 27922 470282 27978
rect 470338 27922 470406 27978
rect 470462 27922 470558 27978
rect 469938 10350 470558 27922
rect 469938 10294 470034 10350
rect 470090 10294 470158 10350
rect 470214 10294 470282 10350
rect 470338 10294 470406 10350
rect 470462 10294 470558 10350
rect 469938 10226 470558 10294
rect 469938 10170 470034 10226
rect 470090 10170 470158 10226
rect 470214 10170 470282 10226
rect 470338 10170 470406 10226
rect 470462 10170 470558 10226
rect 469938 10102 470558 10170
rect 469938 10046 470034 10102
rect 470090 10046 470158 10102
rect 470214 10046 470282 10102
rect 470338 10046 470406 10102
rect 470462 10046 470558 10102
rect 469938 9978 470558 10046
rect 469938 9922 470034 9978
rect 470090 9922 470158 9978
rect 470214 9922 470282 9978
rect 470338 9922 470406 9978
rect 470462 9922 470558 9978
rect 469938 -1120 470558 9922
rect 469938 -1176 470034 -1120
rect 470090 -1176 470158 -1120
rect 470214 -1176 470282 -1120
rect 470338 -1176 470406 -1120
rect 470462 -1176 470558 -1120
rect 469938 -1244 470558 -1176
rect 469938 -1300 470034 -1244
rect 470090 -1300 470158 -1244
rect 470214 -1300 470282 -1244
rect 470338 -1300 470406 -1244
rect 470462 -1300 470558 -1244
rect 469938 -1368 470558 -1300
rect 469938 -1424 470034 -1368
rect 470090 -1424 470158 -1368
rect 470214 -1424 470282 -1368
rect 470338 -1424 470406 -1368
rect 470462 -1424 470558 -1368
rect 469938 -1492 470558 -1424
rect 469938 -1548 470034 -1492
rect 470090 -1548 470158 -1492
rect 470214 -1548 470282 -1492
rect 470338 -1548 470406 -1492
rect 470462 -1548 470558 -1492
rect 469938 -1644 470558 -1548
rect 496938 40350 497558 48690
rect 496938 40294 497034 40350
rect 497090 40294 497158 40350
rect 497214 40294 497282 40350
rect 497338 40294 497406 40350
rect 497462 40294 497558 40350
rect 496938 40226 497558 40294
rect 496938 40170 497034 40226
rect 497090 40170 497158 40226
rect 497214 40170 497282 40226
rect 497338 40170 497406 40226
rect 497462 40170 497558 40226
rect 496938 40102 497558 40170
rect 496938 40046 497034 40102
rect 497090 40046 497158 40102
rect 497214 40046 497282 40102
rect 497338 40046 497406 40102
rect 497462 40046 497558 40102
rect 496938 39978 497558 40046
rect 496938 39922 497034 39978
rect 497090 39922 497158 39978
rect 497214 39922 497282 39978
rect 497338 39922 497406 39978
rect 497462 39922 497558 39978
rect 496938 22350 497558 39922
rect 496938 22294 497034 22350
rect 497090 22294 497158 22350
rect 497214 22294 497282 22350
rect 497338 22294 497406 22350
rect 497462 22294 497558 22350
rect 496938 22226 497558 22294
rect 496938 22170 497034 22226
rect 497090 22170 497158 22226
rect 497214 22170 497282 22226
rect 497338 22170 497406 22226
rect 497462 22170 497558 22226
rect 496938 22102 497558 22170
rect 496938 22046 497034 22102
rect 497090 22046 497158 22102
rect 497214 22046 497282 22102
rect 497338 22046 497406 22102
rect 497462 22046 497558 22102
rect 496938 21978 497558 22046
rect 496938 21922 497034 21978
rect 497090 21922 497158 21978
rect 497214 21922 497282 21978
rect 497338 21922 497406 21978
rect 497462 21922 497558 21978
rect 496938 4350 497558 21922
rect 496938 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 497558 4350
rect 496938 4226 497558 4294
rect 496938 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 497558 4226
rect 496938 4102 497558 4170
rect 496938 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 497558 4102
rect 496938 3978 497558 4046
rect 496938 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 497558 3978
rect 496938 -160 497558 3922
rect 496938 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 497558 -160
rect 496938 -284 497558 -216
rect 496938 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 497558 -284
rect 496938 -408 497558 -340
rect 496938 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 497558 -408
rect 496938 -532 497558 -464
rect 496938 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 497558 -532
rect 496938 -1644 497558 -588
rect 500658 46350 501278 48690
rect 500658 46294 500754 46350
rect 500810 46294 500878 46350
rect 500934 46294 501002 46350
rect 501058 46294 501126 46350
rect 501182 46294 501278 46350
rect 500658 46226 501278 46294
rect 500658 46170 500754 46226
rect 500810 46170 500878 46226
rect 500934 46170 501002 46226
rect 501058 46170 501126 46226
rect 501182 46170 501278 46226
rect 500658 46102 501278 46170
rect 500658 46046 500754 46102
rect 500810 46046 500878 46102
rect 500934 46046 501002 46102
rect 501058 46046 501126 46102
rect 501182 46046 501278 46102
rect 500658 45978 501278 46046
rect 500658 45922 500754 45978
rect 500810 45922 500878 45978
rect 500934 45922 501002 45978
rect 501058 45922 501126 45978
rect 501182 45922 501278 45978
rect 500658 28350 501278 45922
rect 500658 28294 500754 28350
rect 500810 28294 500878 28350
rect 500934 28294 501002 28350
rect 501058 28294 501126 28350
rect 501182 28294 501278 28350
rect 500658 28226 501278 28294
rect 500658 28170 500754 28226
rect 500810 28170 500878 28226
rect 500934 28170 501002 28226
rect 501058 28170 501126 28226
rect 501182 28170 501278 28226
rect 500658 28102 501278 28170
rect 500658 28046 500754 28102
rect 500810 28046 500878 28102
rect 500934 28046 501002 28102
rect 501058 28046 501126 28102
rect 501182 28046 501278 28102
rect 500658 27978 501278 28046
rect 500658 27922 500754 27978
rect 500810 27922 500878 27978
rect 500934 27922 501002 27978
rect 501058 27922 501126 27978
rect 501182 27922 501278 27978
rect 500658 10350 501278 27922
rect 500658 10294 500754 10350
rect 500810 10294 500878 10350
rect 500934 10294 501002 10350
rect 501058 10294 501126 10350
rect 501182 10294 501278 10350
rect 500658 10226 501278 10294
rect 500658 10170 500754 10226
rect 500810 10170 500878 10226
rect 500934 10170 501002 10226
rect 501058 10170 501126 10226
rect 501182 10170 501278 10226
rect 500658 10102 501278 10170
rect 500658 10046 500754 10102
rect 500810 10046 500878 10102
rect 500934 10046 501002 10102
rect 501058 10046 501126 10102
rect 501182 10046 501278 10102
rect 500658 9978 501278 10046
rect 500658 9922 500754 9978
rect 500810 9922 500878 9978
rect 500934 9922 501002 9978
rect 501058 9922 501126 9978
rect 501182 9922 501278 9978
rect 500658 -1120 501278 9922
rect 500658 -1176 500754 -1120
rect 500810 -1176 500878 -1120
rect 500934 -1176 501002 -1120
rect 501058 -1176 501126 -1120
rect 501182 -1176 501278 -1120
rect 500658 -1244 501278 -1176
rect 500658 -1300 500754 -1244
rect 500810 -1300 500878 -1244
rect 500934 -1300 501002 -1244
rect 501058 -1300 501126 -1244
rect 501182 -1300 501278 -1244
rect 500658 -1368 501278 -1300
rect 500658 -1424 500754 -1368
rect 500810 -1424 500878 -1368
rect 500934 -1424 501002 -1368
rect 501058 -1424 501126 -1368
rect 501182 -1424 501278 -1368
rect 500658 -1492 501278 -1424
rect 500658 -1548 500754 -1492
rect 500810 -1548 500878 -1492
rect 500934 -1548 501002 -1492
rect 501058 -1548 501126 -1492
rect 501182 -1548 501278 -1492
rect 500658 -1644 501278 -1548
rect 527658 40350 528278 48690
rect 527658 40294 527754 40350
rect 527810 40294 527878 40350
rect 527934 40294 528002 40350
rect 528058 40294 528126 40350
rect 528182 40294 528278 40350
rect 527658 40226 528278 40294
rect 527658 40170 527754 40226
rect 527810 40170 527878 40226
rect 527934 40170 528002 40226
rect 528058 40170 528126 40226
rect 528182 40170 528278 40226
rect 527658 40102 528278 40170
rect 527658 40046 527754 40102
rect 527810 40046 527878 40102
rect 527934 40046 528002 40102
rect 528058 40046 528126 40102
rect 528182 40046 528278 40102
rect 527658 39978 528278 40046
rect 527658 39922 527754 39978
rect 527810 39922 527878 39978
rect 527934 39922 528002 39978
rect 528058 39922 528126 39978
rect 528182 39922 528278 39978
rect 527658 22350 528278 39922
rect 527658 22294 527754 22350
rect 527810 22294 527878 22350
rect 527934 22294 528002 22350
rect 528058 22294 528126 22350
rect 528182 22294 528278 22350
rect 527658 22226 528278 22294
rect 527658 22170 527754 22226
rect 527810 22170 527878 22226
rect 527934 22170 528002 22226
rect 528058 22170 528126 22226
rect 528182 22170 528278 22226
rect 527658 22102 528278 22170
rect 527658 22046 527754 22102
rect 527810 22046 527878 22102
rect 527934 22046 528002 22102
rect 528058 22046 528126 22102
rect 528182 22046 528278 22102
rect 527658 21978 528278 22046
rect 527658 21922 527754 21978
rect 527810 21922 527878 21978
rect 527934 21922 528002 21978
rect 528058 21922 528126 21978
rect 528182 21922 528278 21978
rect 527658 4350 528278 21922
rect 527658 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 528278 4350
rect 527658 4226 528278 4294
rect 527658 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 528278 4226
rect 527658 4102 528278 4170
rect 527658 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 528278 4102
rect 527658 3978 528278 4046
rect 527658 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 528278 3978
rect 527658 -160 528278 3922
rect 527658 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 528278 -160
rect 527658 -284 528278 -216
rect 527658 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 528278 -284
rect 527658 -408 528278 -340
rect 527658 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 528278 -408
rect 527658 -532 528278 -464
rect 527658 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 528278 -532
rect 527658 -1644 528278 -588
rect 531378 46350 531998 48690
rect 531378 46294 531474 46350
rect 531530 46294 531598 46350
rect 531654 46294 531722 46350
rect 531778 46294 531846 46350
rect 531902 46294 531998 46350
rect 531378 46226 531998 46294
rect 531378 46170 531474 46226
rect 531530 46170 531598 46226
rect 531654 46170 531722 46226
rect 531778 46170 531846 46226
rect 531902 46170 531998 46226
rect 531378 46102 531998 46170
rect 531378 46046 531474 46102
rect 531530 46046 531598 46102
rect 531654 46046 531722 46102
rect 531778 46046 531846 46102
rect 531902 46046 531998 46102
rect 531378 45978 531998 46046
rect 531378 45922 531474 45978
rect 531530 45922 531598 45978
rect 531654 45922 531722 45978
rect 531778 45922 531846 45978
rect 531902 45922 531998 45978
rect 531378 28350 531998 45922
rect 531378 28294 531474 28350
rect 531530 28294 531598 28350
rect 531654 28294 531722 28350
rect 531778 28294 531846 28350
rect 531902 28294 531998 28350
rect 531378 28226 531998 28294
rect 531378 28170 531474 28226
rect 531530 28170 531598 28226
rect 531654 28170 531722 28226
rect 531778 28170 531846 28226
rect 531902 28170 531998 28226
rect 531378 28102 531998 28170
rect 531378 28046 531474 28102
rect 531530 28046 531598 28102
rect 531654 28046 531722 28102
rect 531778 28046 531846 28102
rect 531902 28046 531998 28102
rect 531378 27978 531998 28046
rect 531378 27922 531474 27978
rect 531530 27922 531598 27978
rect 531654 27922 531722 27978
rect 531778 27922 531846 27978
rect 531902 27922 531998 27978
rect 531378 10350 531998 27922
rect 531378 10294 531474 10350
rect 531530 10294 531598 10350
rect 531654 10294 531722 10350
rect 531778 10294 531846 10350
rect 531902 10294 531998 10350
rect 531378 10226 531998 10294
rect 531378 10170 531474 10226
rect 531530 10170 531598 10226
rect 531654 10170 531722 10226
rect 531778 10170 531846 10226
rect 531902 10170 531998 10226
rect 531378 10102 531998 10170
rect 531378 10046 531474 10102
rect 531530 10046 531598 10102
rect 531654 10046 531722 10102
rect 531778 10046 531846 10102
rect 531902 10046 531998 10102
rect 531378 9978 531998 10046
rect 531378 9922 531474 9978
rect 531530 9922 531598 9978
rect 531654 9922 531722 9978
rect 531778 9922 531846 9978
rect 531902 9922 531998 9978
rect 531378 -1120 531998 9922
rect 531378 -1176 531474 -1120
rect 531530 -1176 531598 -1120
rect 531654 -1176 531722 -1120
rect 531778 -1176 531846 -1120
rect 531902 -1176 531998 -1120
rect 531378 -1244 531998 -1176
rect 531378 -1300 531474 -1244
rect 531530 -1300 531598 -1244
rect 531654 -1300 531722 -1244
rect 531778 -1300 531846 -1244
rect 531902 -1300 531998 -1244
rect 531378 -1368 531998 -1300
rect 531378 -1424 531474 -1368
rect 531530 -1424 531598 -1368
rect 531654 -1424 531722 -1368
rect 531778 -1424 531846 -1368
rect 531902 -1424 531998 -1368
rect 531378 -1492 531998 -1424
rect 531378 -1548 531474 -1492
rect 531530 -1548 531598 -1492
rect 531654 -1548 531722 -1492
rect 531778 -1548 531846 -1492
rect 531902 -1548 531998 -1492
rect 531378 -1644 531998 -1548
rect 558378 40350 558998 48690
rect 558378 40294 558474 40350
rect 558530 40294 558598 40350
rect 558654 40294 558722 40350
rect 558778 40294 558846 40350
rect 558902 40294 558998 40350
rect 558378 40226 558998 40294
rect 558378 40170 558474 40226
rect 558530 40170 558598 40226
rect 558654 40170 558722 40226
rect 558778 40170 558846 40226
rect 558902 40170 558998 40226
rect 558378 40102 558998 40170
rect 558378 40046 558474 40102
rect 558530 40046 558598 40102
rect 558654 40046 558722 40102
rect 558778 40046 558846 40102
rect 558902 40046 558998 40102
rect 558378 39978 558998 40046
rect 558378 39922 558474 39978
rect 558530 39922 558598 39978
rect 558654 39922 558722 39978
rect 558778 39922 558846 39978
rect 558902 39922 558998 39978
rect 558378 22350 558998 39922
rect 558378 22294 558474 22350
rect 558530 22294 558598 22350
rect 558654 22294 558722 22350
rect 558778 22294 558846 22350
rect 558902 22294 558998 22350
rect 558378 22226 558998 22294
rect 558378 22170 558474 22226
rect 558530 22170 558598 22226
rect 558654 22170 558722 22226
rect 558778 22170 558846 22226
rect 558902 22170 558998 22226
rect 558378 22102 558998 22170
rect 558378 22046 558474 22102
rect 558530 22046 558598 22102
rect 558654 22046 558722 22102
rect 558778 22046 558846 22102
rect 558902 22046 558998 22102
rect 558378 21978 558998 22046
rect 558378 21922 558474 21978
rect 558530 21922 558598 21978
rect 558654 21922 558722 21978
rect 558778 21922 558846 21978
rect 558902 21922 558998 21978
rect 558378 4350 558998 21922
rect 558378 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 558998 4350
rect 558378 4226 558998 4294
rect 558378 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 558998 4226
rect 558378 4102 558998 4170
rect 558378 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 558998 4102
rect 558378 3978 558998 4046
rect 558378 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 558998 3978
rect 558378 -160 558998 3922
rect 558378 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 558998 -160
rect 558378 -284 558998 -216
rect 558378 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 558998 -284
rect 558378 -408 558998 -340
rect 558378 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 558998 -408
rect 558378 -532 558998 -464
rect 558378 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 558998 -532
rect 558378 -1644 558998 -588
rect 562098 46350 562718 63922
rect 562940 63028 562996 147980
rect 563052 64596 563108 148092
rect 563164 66164 563220 148652
rect 563276 69300 563332 331772
rect 563276 69234 563332 69244
rect 563164 66098 563220 66108
rect 563052 64530 563108 64540
rect 562940 62962 562996 62972
rect 562828 59892 562884 59902
rect 562828 50372 562884 59836
rect 564508 58978 564564 335356
rect 564620 72436 564676 346556
rect 564732 75572 564788 348796
rect 564844 81844 564900 353276
rect 564956 97524 565012 362012
rect 566524 360052 566580 360062
rect 566412 354452 566468 354462
rect 564956 97458 565012 97468
rect 566188 349972 566244 349982
rect 564844 81778 564900 81788
rect 566188 77140 566244 349916
rect 566188 77074 566244 77084
rect 566300 347732 566356 347742
rect 564732 75506 564788 75516
rect 566300 74004 566356 347676
rect 566412 83412 566468 354396
rect 566524 91252 566580 359996
rect 567980 351092 568036 351102
rect 566524 91186 566580 91196
rect 567868 336532 567924 336542
rect 566412 83346 566468 83356
rect 566300 73938 566356 73948
rect 564620 72370 564676 72380
rect 564396 58922 564564 58978
rect 564396 56756 564452 58922
rect 567868 58884 567924 336476
rect 567980 78708 568036 351036
rect 568092 350308 568148 350318
rect 568092 80276 568148 350252
rect 568204 100660 568260 366716
rect 571452 363412 571508 363422
rect 571340 358932 571396 358942
rect 569772 358708 569828 358718
rect 568204 100594 568260 100604
rect 569548 356692 569604 356702
rect 569548 86548 569604 356636
rect 569548 86482 569604 86492
rect 569660 355572 569716 355582
rect 569660 84980 569716 355516
rect 569772 92820 569828 358652
rect 569772 92754 569828 92764
rect 571228 357812 571284 357822
rect 571228 88116 571284 357756
rect 571340 89684 571396 358876
rect 571452 95956 571508 363356
rect 571564 105364 571620 368732
rect 573020 365652 573076 365662
rect 571564 105298 571620 105308
rect 572908 362292 572964 362302
rect 571452 95890 571508 95900
rect 572908 94388 572964 362236
rect 573020 99092 573076 365596
rect 573132 103796 573188 368956
rect 574700 367892 574756 367902
rect 573132 103730 573188 103740
rect 574588 338772 574644 338782
rect 573020 99026 573076 99036
rect 572908 94322 572964 94332
rect 571340 89618 571396 89628
rect 571228 88050 571284 88060
rect 569660 84914 569716 84924
rect 568092 80210 568148 80220
rect 567980 78642 568036 78652
rect 574588 61460 574644 338716
rect 574700 102228 574756 367836
rect 574700 102162 574756 102172
rect 574588 61394 574644 61404
rect 577052 60004 577108 389762
rect 582988 385498 583044 385508
rect 577052 59938 577108 59948
rect 579628 385318 579684 385328
rect 567868 58818 567924 58828
rect 564396 56690 564452 56700
rect 562828 50306 562884 50316
rect 562098 46294 562194 46350
rect 562250 46294 562318 46350
rect 562374 46294 562442 46350
rect 562498 46294 562566 46350
rect 562622 46294 562718 46350
rect 562098 46226 562718 46294
rect 562098 46170 562194 46226
rect 562250 46170 562318 46226
rect 562374 46170 562442 46226
rect 562498 46170 562566 46226
rect 562622 46170 562718 46226
rect 562098 46102 562718 46170
rect 562098 46046 562194 46102
rect 562250 46046 562318 46102
rect 562374 46046 562442 46102
rect 562498 46046 562566 46102
rect 562622 46046 562718 46102
rect 562098 45978 562718 46046
rect 562098 45922 562194 45978
rect 562250 45922 562318 45978
rect 562374 45922 562442 45978
rect 562498 45922 562566 45978
rect 562622 45922 562718 45978
rect 562098 28350 562718 45922
rect 562098 28294 562194 28350
rect 562250 28294 562318 28350
rect 562374 28294 562442 28350
rect 562498 28294 562566 28350
rect 562622 28294 562718 28350
rect 562098 28226 562718 28294
rect 562098 28170 562194 28226
rect 562250 28170 562318 28226
rect 562374 28170 562442 28226
rect 562498 28170 562566 28226
rect 562622 28170 562718 28226
rect 562098 28102 562718 28170
rect 562098 28046 562194 28102
rect 562250 28046 562318 28102
rect 562374 28046 562442 28102
rect 562498 28046 562566 28102
rect 562622 28046 562718 28102
rect 562098 27978 562718 28046
rect 562098 27922 562194 27978
rect 562250 27922 562318 27978
rect 562374 27922 562442 27978
rect 562498 27922 562566 27978
rect 562622 27922 562718 27978
rect 562098 10350 562718 27922
rect 562098 10294 562194 10350
rect 562250 10294 562318 10350
rect 562374 10294 562442 10350
rect 562498 10294 562566 10350
rect 562622 10294 562718 10350
rect 562098 10226 562718 10294
rect 562098 10170 562194 10226
rect 562250 10170 562318 10226
rect 562374 10170 562442 10226
rect 562498 10170 562566 10226
rect 562622 10170 562718 10226
rect 562098 10102 562718 10170
rect 562098 10046 562194 10102
rect 562250 10046 562318 10102
rect 562374 10046 562442 10102
rect 562498 10046 562566 10102
rect 562622 10046 562718 10102
rect 562098 9978 562718 10046
rect 562098 9922 562194 9978
rect 562250 9922 562318 9978
rect 562374 9922 562442 9978
rect 562498 9922 562566 9978
rect 562622 9922 562718 9978
rect 562098 -1120 562718 9922
rect 579628 4228 579684 385262
rect 579628 4162 579684 4172
rect 582988 4228 583044 385442
rect 582988 4162 583044 4172
rect 589098 382350 589718 399922
rect 590492 588644 590548 588654
rect 590492 399028 590548 588588
rect 592818 586350 593438 597744
rect 597360 598172 597980 598268
rect 597360 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect 597360 598048 597980 598116
rect 597360 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect 597360 597924 597980 597992
rect 597360 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect 597360 597800 597980 597868
rect 597360 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect 592818 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 593438 586350
rect 592818 586226 593438 586294
rect 592818 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 593438 586226
rect 592818 586102 593438 586170
rect 592818 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 593438 586102
rect 592818 585978 593438 586046
rect 592818 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 593438 585978
rect 592818 568350 593438 585922
rect 592818 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 593438 568350
rect 592818 568226 593438 568294
rect 592818 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 593438 568226
rect 592818 568102 593438 568170
rect 592818 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 593438 568102
rect 592818 567978 593438 568046
rect 592818 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 593438 567978
rect 592818 550350 593438 567922
rect 592818 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 593438 550350
rect 592818 550226 593438 550294
rect 592818 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 593438 550226
rect 592818 550102 593438 550170
rect 592818 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 593438 550102
rect 592818 549978 593438 550046
rect 592818 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 593438 549978
rect 590604 548996 590660 549006
rect 590604 402500 590660 548940
rect 592818 532350 593438 549922
rect 592818 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 593438 532350
rect 592818 532226 593438 532294
rect 592818 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 593438 532226
rect 592818 532102 593438 532170
rect 592818 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 593438 532102
rect 592818 531978 593438 532046
rect 592818 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 593438 531978
rect 592818 514350 593438 531922
rect 592818 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 593438 514350
rect 592818 514226 593438 514294
rect 592818 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 593438 514226
rect 592818 514102 593438 514170
rect 592818 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 593438 514102
rect 592818 513978 593438 514046
rect 592818 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 593438 513978
rect 590604 402434 590660 402444
rect 590716 509348 590772 509358
rect 590492 398962 590548 398972
rect 590716 397348 590772 509292
rect 592818 496350 593438 513922
rect 592818 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 593438 496350
rect 592818 496226 593438 496294
rect 592818 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 593438 496226
rect 592818 496102 593438 496170
rect 592818 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 593438 496102
rect 592818 495978 593438 496046
rect 592818 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 593438 495978
rect 592818 478350 593438 495922
rect 592818 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 593438 478350
rect 592818 478226 593438 478294
rect 592818 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 593438 478226
rect 592818 478102 593438 478170
rect 592818 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 593438 478102
rect 592818 477978 593438 478046
rect 592818 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 593438 477978
rect 590828 469700 590884 469710
rect 590828 404038 590884 469644
rect 592818 460350 593438 477922
rect 592818 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 593438 460350
rect 592818 460226 593438 460294
rect 592818 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 593438 460226
rect 592818 460102 593438 460170
rect 592818 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 593438 460102
rect 592818 459978 593438 460046
rect 592818 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 593438 459978
rect 592818 442350 593438 459922
rect 592818 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 593438 442350
rect 592818 442226 593438 442294
rect 592818 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 593438 442226
rect 592818 442102 593438 442170
rect 592818 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 593438 442102
rect 592818 441978 593438 442046
rect 592818 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 593438 441978
rect 590828 403972 590884 403982
rect 590940 430164 590996 430174
rect 590940 402388 590996 430108
rect 590940 402322 590996 402332
rect 592818 424350 593438 441922
rect 592818 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 593438 424350
rect 592818 424226 593438 424294
rect 592818 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 593438 424226
rect 592818 424102 593438 424170
rect 592818 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 593438 424102
rect 592818 423978 593438 424046
rect 592818 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 593438 423978
rect 592818 406350 593438 423922
rect 592818 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 593438 406350
rect 592818 406226 593438 406294
rect 592818 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 593438 406226
rect 592818 406102 593438 406170
rect 592818 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 593438 406102
rect 592818 405978 593438 406046
rect 592818 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 593438 405978
rect 590716 397282 590772 397292
rect 590156 390404 590212 390414
rect 590156 387268 590212 390348
rect 590156 387202 590212 387212
rect 592818 388350 593438 405922
rect 592818 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 593438 388350
rect 592818 388226 593438 388294
rect 592818 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 593438 388226
rect 592818 388102 593438 388170
rect 592818 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 593438 388102
rect 592818 387978 593438 388046
rect 592818 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 593438 387978
rect 589098 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 589718 382350
rect 589098 382226 589718 382294
rect 589098 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 589718 382226
rect 589098 382102 589718 382170
rect 589098 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 589718 382102
rect 589098 381978 589718 382046
rect 589098 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 589718 381978
rect 589098 364350 589718 381922
rect 589098 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 589718 364350
rect 589098 364226 589718 364294
rect 589098 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 589718 364226
rect 589098 364102 589718 364170
rect 589098 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 589718 364102
rect 589098 363978 589718 364046
rect 589098 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 589718 363978
rect 589098 346350 589718 363922
rect 592818 370350 593438 387922
rect 592818 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 593438 370350
rect 592818 370226 593438 370294
rect 592818 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 593438 370226
rect 592818 370102 593438 370170
rect 592818 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 593438 370102
rect 592818 369978 593438 370046
rect 592818 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 593438 369978
rect 592818 352350 593438 369922
rect 592818 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 593438 352350
rect 592818 352226 593438 352294
rect 592818 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 593438 352226
rect 592818 352102 593438 352170
rect 592818 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 593438 352102
rect 592818 351978 593438 352046
rect 592818 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 593438 351978
rect 589098 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 589718 346350
rect 589098 346226 589718 346294
rect 589098 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 589718 346226
rect 589098 346102 589718 346170
rect 589098 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 589718 346102
rect 589098 345978 589718 346046
rect 589098 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 589718 345978
rect 589098 328350 589718 345922
rect 589098 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 589718 328350
rect 589098 328226 589718 328294
rect 589098 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 589718 328226
rect 589098 328102 589718 328170
rect 589098 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 589718 328102
rect 589098 327978 589718 328046
rect 589098 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 589718 327978
rect 589098 310350 589718 327922
rect 589098 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 589718 310350
rect 589098 310226 589718 310294
rect 589098 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 589718 310226
rect 589098 310102 589718 310170
rect 589098 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 589718 310102
rect 589098 309978 589718 310046
rect 589098 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 589718 309978
rect 589098 292350 589718 309922
rect 589098 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 589718 292350
rect 589098 292226 589718 292294
rect 589098 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 589718 292226
rect 589098 292102 589718 292170
rect 589098 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 589718 292102
rect 589098 291978 589718 292046
rect 589098 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 589718 291978
rect 589098 274350 589718 291922
rect 589098 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 589718 274350
rect 589098 274226 589718 274294
rect 589098 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 589718 274226
rect 589098 274102 589718 274170
rect 589098 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 589718 274102
rect 589098 273978 589718 274046
rect 589098 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 589718 273978
rect 589098 256350 589718 273922
rect 590492 350756 590548 350766
rect 590492 256564 590548 350700
rect 592818 334350 593438 351922
rect 592818 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 593438 334350
rect 592818 334226 593438 334294
rect 592818 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 593438 334226
rect 592818 334102 593438 334170
rect 592818 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 593438 334102
rect 592818 333978 593438 334046
rect 592818 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 593438 333978
rect 592818 316350 593438 333922
rect 592818 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 593438 316350
rect 592818 316226 593438 316294
rect 592818 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 593438 316226
rect 592818 316102 593438 316170
rect 592818 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 593438 316102
rect 592818 315978 593438 316046
rect 592818 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 593438 315978
rect 590492 256498 590548 256508
rect 590604 311108 590660 311118
rect 589098 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 589718 256350
rect 589098 256226 589718 256294
rect 589098 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 589718 256226
rect 589098 256102 589718 256170
rect 589098 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 589718 256102
rect 589098 255978 589718 256046
rect 589098 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 589718 255978
rect 589098 238350 589718 255922
rect 590604 255332 590660 311052
rect 592818 298350 593438 315922
rect 592818 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 593438 298350
rect 592818 298226 593438 298294
rect 592818 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 593438 298226
rect 592818 298102 593438 298170
rect 592818 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 593438 298102
rect 592818 297978 593438 298046
rect 592818 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 593438 297978
rect 592818 280350 593438 297922
rect 592818 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 593438 280350
rect 592818 280226 593438 280294
rect 592818 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 593438 280226
rect 592818 280102 593438 280170
rect 592818 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 593438 280102
rect 592818 279978 593438 280046
rect 592818 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 593438 279978
rect 590604 255266 590660 255276
rect 590828 271460 590884 271470
rect 590828 255220 590884 271404
rect 590828 255154 590884 255164
rect 592818 262350 593438 279922
rect 592818 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 593438 262350
rect 592818 262226 593438 262294
rect 592818 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 593438 262226
rect 592818 262102 593438 262170
rect 592818 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 593438 262102
rect 592818 261978 593438 262046
rect 592818 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 593438 261978
rect 592818 244350 593438 261922
rect 592818 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 593438 244350
rect 592818 244226 593438 244294
rect 592818 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 593438 244226
rect 592818 244102 593438 244170
rect 592818 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 593438 244102
rect 592818 243978 593438 244046
rect 592818 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 593438 243978
rect 590828 241108 590884 241118
rect 589098 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 589718 238350
rect 589098 238226 589718 238294
rect 589098 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 589718 238226
rect 589098 238102 589718 238170
rect 589098 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 589718 238102
rect 589098 237978 589718 238046
rect 589098 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 589718 237978
rect 589098 220350 589718 237922
rect 590156 239540 590212 239550
rect 590156 232036 590212 239484
rect 590604 239428 590660 239438
rect 590156 231970 590212 231980
rect 590492 236516 590548 236526
rect 589098 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 589718 220350
rect 589098 220226 589718 220294
rect 589098 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 589718 220226
rect 589098 220102 589718 220170
rect 589098 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 589718 220102
rect 589098 219978 589718 220046
rect 589098 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 589718 219978
rect 589098 202350 589718 219922
rect 589098 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 589718 202350
rect 589098 202226 589718 202294
rect 589098 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 589718 202226
rect 589098 202102 589718 202170
rect 589098 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 589718 202102
rect 589098 201978 589718 202046
rect 589098 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 589718 201978
rect 589098 184350 589718 201922
rect 589098 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 589718 184350
rect 589098 184226 589718 184294
rect 589098 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 589718 184226
rect 589098 184102 589718 184170
rect 589098 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 589718 184102
rect 589098 183978 589718 184046
rect 589098 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 589718 183978
rect 589098 166350 589718 183922
rect 589098 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 589718 166350
rect 589098 166226 589718 166294
rect 589098 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 589718 166226
rect 589098 166102 589718 166170
rect 589098 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 589718 166102
rect 589098 165978 589718 166046
rect 589098 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 589718 165978
rect 589098 148350 589718 165922
rect 589098 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 589718 148350
rect 589098 148226 589718 148294
rect 589098 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 589718 148226
rect 589098 148102 589718 148170
rect 589098 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 589718 148102
rect 589098 147978 589718 148046
rect 589098 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 589718 147978
rect 589098 130350 589718 147922
rect 589098 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 589718 130350
rect 589098 130226 589718 130294
rect 589098 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 589718 130226
rect 589098 130102 589718 130170
rect 589098 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 589718 130102
rect 589098 129978 589718 130046
rect 589098 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 589718 129978
rect 589098 112350 589718 129922
rect 589098 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 589718 112350
rect 589098 112226 589718 112294
rect 589098 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 589718 112226
rect 589098 112102 589718 112170
rect 589098 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 589718 112102
rect 589098 111978 589718 112046
rect 589098 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 589718 111978
rect 589098 94350 589718 111922
rect 589098 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 589718 94350
rect 589098 94226 589718 94294
rect 589098 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 589718 94226
rect 589098 94102 589718 94170
rect 589098 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 589718 94102
rect 589098 93978 589718 94046
rect 589098 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 589718 93978
rect 589098 76350 589718 93922
rect 589098 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 589718 76350
rect 589098 76226 589718 76294
rect 589098 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 589718 76226
rect 589098 76102 589718 76170
rect 589098 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 589718 76102
rect 589098 75978 589718 76046
rect 589098 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 589718 75978
rect 589098 58350 589718 75922
rect 590492 73444 590548 236460
rect 590604 113092 590660 239372
rect 590716 236404 590772 236414
rect 590716 152740 590772 236348
rect 590828 192388 590884 241052
rect 590828 192322 590884 192332
rect 592818 226350 593438 243922
rect 592818 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 593438 226350
rect 592818 226226 593438 226294
rect 592818 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 593438 226226
rect 592818 226102 593438 226170
rect 592818 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 593438 226102
rect 592818 225978 593438 226046
rect 592818 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 593438 225978
rect 592818 208350 593438 225922
rect 592818 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 593438 208350
rect 592818 208226 593438 208294
rect 592818 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 593438 208226
rect 592818 208102 593438 208170
rect 592818 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 593438 208102
rect 592818 207978 593438 208046
rect 592818 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 593438 207978
rect 590716 152674 590772 152684
rect 592818 190350 593438 207922
rect 592818 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 593438 190350
rect 592818 190226 593438 190294
rect 592818 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 593438 190226
rect 592818 190102 593438 190170
rect 592818 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 593438 190102
rect 592818 189978 593438 190046
rect 592818 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 593438 189978
rect 592818 172350 593438 189922
rect 592818 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 593438 172350
rect 592818 172226 593438 172294
rect 592818 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 593438 172226
rect 592818 172102 593438 172170
rect 592818 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 593438 172102
rect 592818 171978 593438 172046
rect 592818 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 593438 171978
rect 592818 154350 593438 171922
rect 592818 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 593438 154350
rect 592818 154226 593438 154294
rect 592818 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 593438 154226
rect 592818 154102 593438 154170
rect 592818 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 593438 154102
rect 592818 153978 593438 154046
rect 592818 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 593438 153978
rect 590604 113026 590660 113036
rect 592818 136350 593438 153922
rect 592818 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 593438 136350
rect 592818 136226 593438 136294
rect 592818 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 593438 136226
rect 592818 136102 593438 136170
rect 592818 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 593438 136102
rect 592818 135978 593438 136046
rect 592818 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 593438 135978
rect 592818 118350 593438 135922
rect 592818 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 593438 118350
rect 592818 118226 593438 118294
rect 592818 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 593438 118226
rect 592818 118102 593438 118170
rect 592818 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 593438 118102
rect 592818 117978 593438 118046
rect 592818 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 593438 117978
rect 590492 73378 590548 73388
rect 592818 100350 593438 117922
rect 592818 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 593438 100350
rect 592818 100226 593438 100294
rect 592818 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 593438 100226
rect 592818 100102 593438 100170
rect 592818 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 593438 100102
rect 592818 99978 593438 100046
rect 592818 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 593438 99978
rect 592818 82350 593438 99922
rect 592818 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 593438 82350
rect 592818 82226 593438 82294
rect 592818 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 593438 82226
rect 592818 82102 593438 82170
rect 592818 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 593438 82102
rect 592818 81978 593438 82046
rect 592818 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 593438 81978
rect 589098 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 589718 58350
rect 589098 58226 589718 58294
rect 589098 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 589718 58226
rect 589098 58102 589718 58170
rect 589098 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 589718 58102
rect 589098 57978 589718 58046
rect 589098 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 589718 57978
rect 589098 40350 589718 57922
rect 589098 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 589718 40350
rect 589098 40226 589718 40294
rect 589098 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 589718 40226
rect 589098 40102 589718 40170
rect 589098 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 589718 40102
rect 589098 39978 589718 40046
rect 589098 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 589718 39978
rect 589098 22350 589718 39922
rect 589098 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 589718 22350
rect 589098 22226 589718 22294
rect 589098 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 589718 22226
rect 589098 22102 589718 22170
rect 589098 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 589718 22102
rect 589098 21978 589718 22046
rect 589098 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 589718 21978
rect 589098 4350 589718 21922
rect 589098 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 589718 4350
rect 589098 4226 589718 4294
rect 589098 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 589718 4226
rect 562098 -1176 562194 -1120
rect 562250 -1176 562318 -1120
rect 562374 -1176 562442 -1120
rect 562498 -1176 562566 -1120
rect 562622 -1176 562718 -1120
rect 562098 -1244 562718 -1176
rect 562098 -1300 562194 -1244
rect 562250 -1300 562318 -1244
rect 562374 -1300 562442 -1244
rect 562498 -1300 562566 -1244
rect 562622 -1300 562718 -1244
rect 562098 -1368 562718 -1300
rect 562098 -1424 562194 -1368
rect 562250 -1424 562318 -1368
rect 562374 -1424 562442 -1368
rect 562498 -1424 562566 -1368
rect 562622 -1424 562718 -1368
rect 562098 -1492 562718 -1424
rect 562098 -1548 562194 -1492
rect 562250 -1548 562318 -1492
rect 562374 -1548 562442 -1492
rect 562498 -1548 562566 -1492
rect 562622 -1548 562718 -1492
rect 562098 -1644 562718 -1548
rect 589098 4102 589718 4170
rect 589098 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 589718 4102
rect 589098 3978 589718 4046
rect 589098 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 589718 3978
rect 589098 -160 589718 3922
rect 589098 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 589718 -160
rect 589098 -284 589718 -216
rect 589098 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 589718 -284
rect 589098 -408 589718 -340
rect 589098 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 589718 -408
rect 589098 -532 589718 -464
rect 589098 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 589718 -532
rect 589098 -1644 589718 -588
rect 592818 64350 593438 81922
rect 592818 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 593438 64350
rect 592818 64226 593438 64294
rect 592818 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 593438 64226
rect 592818 64102 593438 64170
rect 592818 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 593438 64102
rect 592818 63978 593438 64046
rect 592818 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 593438 63978
rect 592818 46350 593438 63922
rect 592818 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 593438 46350
rect 592818 46226 593438 46294
rect 592818 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 593438 46226
rect 592818 46102 593438 46170
rect 592818 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 593438 46102
rect 592818 45978 593438 46046
rect 592818 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 593438 45978
rect 592818 28350 593438 45922
rect 592818 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 593438 28350
rect 592818 28226 593438 28294
rect 592818 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 593438 28226
rect 592818 28102 593438 28170
rect 592818 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 593438 28102
rect 592818 27978 593438 28046
rect 592818 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 593438 27978
rect 592818 10350 593438 27922
rect 592818 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 593438 10350
rect 592818 10226 593438 10294
rect 592818 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 593438 10226
rect 592818 10102 593438 10170
rect 592818 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 593438 10102
rect 592818 9978 593438 10046
rect 592818 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 593438 9978
rect 592818 -1120 593438 9922
rect 596400 597212 597020 597308
rect 596400 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect 596400 597088 597020 597156
rect 596400 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect 596400 596964 597020 597032
rect 596400 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect 596400 596840 597020 596908
rect 596400 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect 596400 580350 597020 596784
rect 596400 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597020 580350
rect 596400 580226 597020 580294
rect 596400 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597020 580226
rect 596400 580102 597020 580170
rect 596400 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597020 580102
rect 596400 579978 597020 580046
rect 596400 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597020 579978
rect 596400 562350 597020 579922
rect 596400 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597020 562350
rect 596400 562226 597020 562294
rect 596400 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597020 562226
rect 596400 562102 597020 562170
rect 596400 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597020 562102
rect 596400 561978 597020 562046
rect 596400 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597020 561978
rect 596400 544350 597020 561922
rect 596400 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597020 544350
rect 596400 544226 597020 544294
rect 596400 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597020 544226
rect 596400 544102 597020 544170
rect 596400 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597020 544102
rect 596400 543978 597020 544046
rect 596400 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597020 543978
rect 596400 526350 597020 543922
rect 596400 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597020 526350
rect 596400 526226 597020 526294
rect 596400 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597020 526226
rect 596400 526102 597020 526170
rect 596400 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597020 526102
rect 596400 525978 597020 526046
rect 596400 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597020 525978
rect 596400 508350 597020 525922
rect 596400 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597020 508350
rect 596400 508226 597020 508294
rect 596400 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597020 508226
rect 596400 508102 597020 508170
rect 596400 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597020 508102
rect 596400 507978 597020 508046
rect 596400 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597020 507978
rect 596400 490350 597020 507922
rect 596400 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597020 490350
rect 596400 490226 597020 490294
rect 596400 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597020 490226
rect 596400 490102 597020 490170
rect 596400 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597020 490102
rect 596400 489978 597020 490046
rect 596400 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597020 489978
rect 596400 472350 597020 489922
rect 596400 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597020 472350
rect 596400 472226 597020 472294
rect 596400 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597020 472226
rect 596400 472102 597020 472170
rect 596400 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597020 472102
rect 596400 471978 597020 472046
rect 596400 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597020 471978
rect 596400 454350 597020 471922
rect 596400 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597020 454350
rect 596400 454226 597020 454294
rect 596400 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597020 454226
rect 596400 454102 597020 454170
rect 596400 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597020 454102
rect 596400 453978 597020 454046
rect 596400 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597020 453978
rect 596400 436350 597020 453922
rect 596400 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597020 436350
rect 596400 436226 597020 436294
rect 596400 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597020 436226
rect 596400 436102 597020 436170
rect 596400 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597020 436102
rect 596400 435978 597020 436046
rect 596400 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597020 435978
rect 596400 418350 597020 435922
rect 596400 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597020 418350
rect 596400 418226 597020 418294
rect 596400 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597020 418226
rect 596400 418102 597020 418170
rect 596400 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597020 418102
rect 596400 417978 597020 418046
rect 596400 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597020 417978
rect 596400 400350 597020 417922
rect 596400 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597020 400350
rect 596400 400226 597020 400294
rect 596400 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597020 400226
rect 596400 400102 597020 400170
rect 596400 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597020 400102
rect 596400 399978 597020 400046
rect 596400 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597020 399978
rect 596400 382350 597020 399922
rect 596400 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597020 382350
rect 596400 382226 597020 382294
rect 596400 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597020 382226
rect 596400 382102 597020 382170
rect 596400 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597020 382102
rect 596400 381978 597020 382046
rect 596400 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597020 381978
rect 596400 364350 597020 381922
rect 596400 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597020 364350
rect 596400 364226 597020 364294
rect 596400 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597020 364226
rect 596400 364102 597020 364170
rect 596400 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597020 364102
rect 596400 363978 597020 364046
rect 596400 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597020 363978
rect 596400 346350 597020 363922
rect 596400 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597020 346350
rect 596400 346226 597020 346294
rect 596400 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597020 346226
rect 596400 346102 597020 346170
rect 596400 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597020 346102
rect 596400 345978 597020 346046
rect 596400 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597020 345978
rect 596400 328350 597020 345922
rect 596400 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597020 328350
rect 596400 328226 597020 328294
rect 596400 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597020 328226
rect 596400 328102 597020 328170
rect 596400 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597020 328102
rect 596400 327978 597020 328046
rect 596400 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597020 327978
rect 596400 310350 597020 327922
rect 596400 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597020 310350
rect 596400 310226 597020 310294
rect 596400 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597020 310226
rect 596400 310102 597020 310170
rect 596400 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597020 310102
rect 596400 309978 597020 310046
rect 596400 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597020 309978
rect 596400 292350 597020 309922
rect 596400 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597020 292350
rect 596400 292226 597020 292294
rect 596400 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597020 292226
rect 596400 292102 597020 292170
rect 596400 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597020 292102
rect 596400 291978 597020 292046
rect 596400 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597020 291978
rect 596400 274350 597020 291922
rect 596400 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597020 274350
rect 596400 274226 597020 274294
rect 596400 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597020 274226
rect 596400 274102 597020 274170
rect 596400 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597020 274102
rect 596400 273978 597020 274046
rect 596400 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597020 273978
rect 596400 256350 597020 273922
rect 596400 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597020 256350
rect 596400 256226 597020 256294
rect 596400 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597020 256226
rect 596400 256102 597020 256170
rect 596400 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597020 256102
rect 596400 255978 597020 256046
rect 596400 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597020 255978
rect 596400 238350 597020 255922
rect 596400 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597020 238350
rect 596400 238226 597020 238294
rect 596400 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597020 238226
rect 596400 238102 597020 238170
rect 596400 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597020 238102
rect 596400 237978 597020 238046
rect 596400 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597020 237978
rect 596400 220350 597020 237922
rect 596400 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597020 220350
rect 596400 220226 597020 220294
rect 596400 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597020 220226
rect 596400 220102 597020 220170
rect 596400 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597020 220102
rect 596400 219978 597020 220046
rect 596400 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597020 219978
rect 596400 202350 597020 219922
rect 596400 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597020 202350
rect 596400 202226 597020 202294
rect 596400 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597020 202226
rect 596400 202102 597020 202170
rect 596400 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597020 202102
rect 596400 201978 597020 202046
rect 596400 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597020 201978
rect 596400 184350 597020 201922
rect 596400 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597020 184350
rect 596400 184226 597020 184294
rect 596400 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597020 184226
rect 596400 184102 597020 184170
rect 596400 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597020 184102
rect 596400 183978 597020 184046
rect 596400 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597020 183978
rect 596400 166350 597020 183922
rect 596400 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597020 166350
rect 596400 166226 597020 166294
rect 596400 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597020 166226
rect 596400 166102 597020 166170
rect 596400 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597020 166102
rect 596400 165978 597020 166046
rect 596400 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597020 165978
rect 596400 148350 597020 165922
rect 596400 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597020 148350
rect 596400 148226 597020 148294
rect 596400 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597020 148226
rect 596400 148102 597020 148170
rect 596400 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597020 148102
rect 596400 147978 597020 148046
rect 596400 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597020 147978
rect 596400 130350 597020 147922
rect 596400 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597020 130350
rect 596400 130226 597020 130294
rect 596400 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597020 130226
rect 596400 130102 597020 130170
rect 596400 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597020 130102
rect 596400 129978 597020 130046
rect 596400 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597020 129978
rect 596400 112350 597020 129922
rect 596400 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597020 112350
rect 596400 112226 597020 112294
rect 596400 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597020 112226
rect 596400 112102 597020 112170
rect 596400 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597020 112102
rect 596400 111978 597020 112046
rect 596400 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597020 111978
rect 596400 94350 597020 111922
rect 596400 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597020 94350
rect 596400 94226 597020 94294
rect 596400 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597020 94226
rect 596400 94102 597020 94170
rect 596400 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597020 94102
rect 596400 93978 597020 94046
rect 596400 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597020 93978
rect 596400 76350 597020 93922
rect 596400 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597020 76350
rect 596400 76226 597020 76294
rect 596400 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597020 76226
rect 596400 76102 597020 76170
rect 596400 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597020 76102
rect 596400 75978 597020 76046
rect 596400 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597020 75978
rect 596400 58350 597020 75922
rect 596400 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597020 58350
rect 596400 58226 597020 58294
rect 596400 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597020 58226
rect 596400 58102 597020 58170
rect 596400 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597020 58102
rect 596400 57978 597020 58046
rect 596400 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597020 57978
rect 596400 40350 597020 57922
rect 596400 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597020 40350
rect 596400 40226 597020 40294
rect 596400 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597020 40226
rect 596400 40102 597020 40170
rect 596400 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597020 40102
rect 596400 39978 597020 40046
rect 596400 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597020 39978
rect 596400 22350 597020 39922
rect 596400 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597020 22350
rect 596400 22226 597020 22294
rect 596400 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597020 22226
rect 596400 22102 597020 22170
rect 596400 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597020 22102
rect 596400 21978 597020 22046
rect 596400 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597020 21978
rect 596400 4350 597020 21922
rect 596400 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597020 4350
rect 596400 4226 597020 4294
rect 596400 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597020 4226
rect 596400 4102 597020 4170
rect 596400 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597020 4102
rect 596400 3978 597020 4046
rect 596400 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597020 3978
rect 596400 -160 597020 3922
rect 596400 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect 596400 -284 597020 -216
rect 596400 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect 596400 -408 597020 -340
rect 596400 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect 596400 -532 597020 -464
rect 596400 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect 596400 -684 597020 -588
rect 597360 586350 597980 597744
rect 597360 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect 597360 586226 597980 586294
rect 597360 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect 597360 586102 597980 586170
rect 597360 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect 597360 585978 597980 586046
rect 597360 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect 597360 568350 597980 585922
rect 597360 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect 597360 568226 597980 568294
rect 597360 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect 597360 568102 597980 568170
rect 597360 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect 597360 567978 597980 568046
rect 597360 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect 597360 550350 597980 567922
rect 597360 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect 597360 550226 597980 550294
rect 597360 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect 597360 550102 597980 550170
rect 597360 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect 597360 549978 597980 550046
rect 597360 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect 597360 532350 597980 549922
rect 597360 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect 597360 532226 597980 532294
rect 597360 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect 597360 532102 597980 532170
rect 597360 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect 597360 531978 597980 532046
rect 597360 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect 597360 514350 597980 531922
rect 597360 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect 597360 514226 597980 514294
rect 597360 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect 597360 514102 597980 514170
rect 597360 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect 597360 513978 597980 514046
rect 597360 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect 597360 496350 597980 513922
rect 597360 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect 597360 496226 597980 496294
rect 597360 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect 597360 496102 597980 496170
rect 597360 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 597360 495978 597980 496046
rect 597360 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect 597360 478350 597980 495922
rect 597360 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect 597360 478226 597980 478294
rect 597360 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect 597360 478102 597980 478170
rect 597360 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect 597360 477978 597980 478046
rect 597360 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect 597360 460350 597980 477922
rect 597360 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect 597360 460226 597980 460294
rect 597360 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect 597360 460102 597980 460170
rect 597360 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect 597360 459978 597980 460046
rect 597360 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect 597360 442350 597980 459922
rect 597360 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect 597360 442226 597980 442294
rect 597360 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect 597360 442102 597980 442170
rect 597360 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect 597360 441978 597980 442046
rect 597360 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect 597360 424350 597980 441922
rect 597360 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect 597360 424226 597980 424294
rect 597360 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect 597360 424102 597980 424170
rect 597360 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect 597360 423978 597980 424046
rect 597360 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect 597360 406350 597980 423922
rect 597360 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect 597360 406226 597980 406294
rect 597360 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect 597360 406102 597980 406170
rect 597360 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect 597360 405978 597980 406046
rect 597360 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect 597360 388350 597980 405922
rect 597360 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect 597360 388226 597980 388294
rect 597360 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect 597360 388102 597980 388170
rect 597360 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect 597360 387978 597980 388046
rect 597360 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect 597360 370350 597980 387922
rect 597360 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect 597360 370226 597980 370294
rect 597360 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect 597360 370102 597980 370170
rect 597360 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect 597360 369978 597980 370046
rect 597360 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect 597360 352350 597980 369922
rect 597360 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect 597360 352226 597980 352294
rect 597360 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect 597360 352102 597980 352170
rect 597360 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect 597360 351978 597980 352046
rect 597360 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect 597360 334350 597980 351922
rect 597360 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect 597360 334226 597980 334294
rect 597360 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect 597360 334102 597980 334170
rect 597360 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect 597360 333978 597980 334046
rect 597360 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect 597360 316350 597980 333922
rect 597360 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect 597360 316226 597980 316294
rect 597360 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect 597360 316102 597980 316170
rect 597360 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect 597360 315978 597980 316046
rect 597360 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect 597360 298350 597980 315922
rect 597360 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect 597360 298226 597980 298294
rect 597360 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect 597360 298102 597980 298170
rect 597360 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect 597360 297978 597980 298046
rect 597360 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect 597360 280350 597980 297922
rect 597360 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect 597360 280226 597980 280294
rect 597360 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect 597360 280102 597980 280170
rect 597360 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect 597360 279978 597980 280046
rect 597360 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect 597360 262350 597980 279922
rect 597360 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect 597360 262226 597980 262294
rect 597360 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect 597360 262102 597980 262170
rect 597360 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect 597360 261978 597980 262046
rect 597360 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect 597360 244350 597980 261922
rect 597360 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect 597360 244226 597980 244294
rect 597360 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect 597360 244102 597980 244170
rect 597360 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect 597360 243978 597980 244046
rect 597360 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect 597360 226350 597980 243922
rect 597360 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect 597360 226226 597980 226294
rect 597360 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect 597360 226102 597980 226170
rect 597360 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect 597360 225978 597980 226046
rect 597360 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect 597360 208350 597980 225922
rect 597360 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect 597360 208226 597980 208294
rect 597360 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect 597360 208102 597980 208170
rect 597360 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect 597360 207978 597980 208046
rect 597360 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect 597360 190350 597980 207922
rect 597360 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect 597360 190226 597980 190294
rect 597360 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect 597360 190102 597980 190170
rect 597360 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect 597360 189978 597980 190046
rect 597360 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect 597360 172350 597980 189922
rect 597360 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect 597360 172226 597980 172294
rect 597360 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect 597360 172102 597980 172170
rect 597360 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect 597360 171978 597980 172046
rect 597360 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect 597360 154350 597980 171922
rect 597360 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect 597360 154226 597980 154294
rect 597360 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect 597360 154102 597980 154170
rect 597360 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect 597360 153978 597980 154046
rect 597360 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect 597360 136350 597980 153922
rect 597360 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect 597360 136226 597980 136294
rect 597360 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect 597360 136102 597980 136170
rect 597360 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect 597360 135978 597980 136046
rect 597360 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect 597360 118350 597980 135922
rect 597360 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect 597360 118226 597980 118294
rect 597360 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect 597360 118102 597980 118170
rect 597360 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect 597360 117978 597980 118046
rect 597360 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect 597360 100350 597980 117922
rect 597360 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect 597360 100226 597980 100294
rect 597360 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect 597360 100102 597980 100170
rect 597360 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect 597360 99978 597980 100046
rect 597360 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect 597360 82350 597980 99922
rect 597360 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect 597360 82226 597980 82294
rect 597360 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect 597360 82102 597980 82170
rect 597360 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect 597360 81978 597980 82046
rect 597360 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 597360 64350 597980 81922
rect 597360 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect 597360 64226 597980 64294
rect 597360 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect 597360 64102 597980 64170
rect 597360 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect 597360 63978 597980 64046
rect 597360 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect 597360 46350 597980 63922
rect 597360 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect 597360 46226 597980 46294
rect 597360 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect 597360 46102 597980 46170
rect 597360 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect 597360 45978 597980 46046
rect 597360 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect 597360 28350 597980 45922
rect 597360 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect 597360 28226 597980 28294
rect 597360 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect 597360 28102 597980 28170
rect 597360 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect 597360 27978 597980 28046
rect 597360 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect 597360 10350 597980 27922
rect 597360 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect 597360 10226 597980 10294
rect 597360 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect 597360 10102 597980 10170
rect 597360 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect 597360 9978 597980 10046
rect 597360 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect 592818 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 593438 -1120
rect 592818 -1244 593438 -1176
rect 592818 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 593438 -1244
rect 592818 -1368 593438 -1300
rect 592818 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 593438 -1368
rect 592818 -1492 593438 -1424
rect 592818 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 593438 -1492
rect 592818 -1644 593438 -1548
rect 597360 -1120 597980 9922
rect 597360 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect 597360 -1244 597980 -1176
rect 597360 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect 597360 -1368 597980 -1300
rect 597360 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect 597360 -1492 597980 -1424
rect 597360 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect 597360 -1644 597980 -1548
<< via4 >>
rect -1820 598116 -1764 598172
rect -1696 598116 -1640 598172
rect -1572 598116 -1516 598172
rect -1448 598116 -1392 598172
rect -1820 597992 -1764 598048
rect -1696 597992 -1640 598048
rect -1572 597992 -1516 598048
rect -1448 597992 -1392 598048
rect -1820 597868 -1764 597924
rect -1696 597868 -1640 597924
rect -1572 597868 -1516 597924
rect -1448 597868 -1392 597924
rect -1820 597744 -1764 597800
rect -1696 597744 -1640 597800
rect -1572 597744 -1516 597800
rect -1448 597744 -1392 597800
rect -1820 586294 -1764 586350
rect -1696 586294 -1640 586350
rect -1572 586294 -1516 586350
rect -1448 586294 -1392 586350
rect -1820 586170 -1764 586226
rect -1696 586170 -1640 586226
rect -1572 586170 -1516 586226
rect -1448 586170 -1392 586226
rect -1820 586046 -1764 586102
rect -1696 586046 -1640 586102
rect -1572 586046 -1516 586102
rect -1448 586046 -1392 586102
rect -1820 585922 -1764 585978
rect -1696 585922 -1640 585978
rect -1572 585922 -1516 585978
rect -1448 585922 -1392 585978
rect -1820 568294 -1764 568350
rect -1696 568294 -1640 568350
rect -1572 568294 -1516 568350
rect -1448 568294 -1392 568350
rect -1820 568170 -1764 568226
rect -1696 568170 -1640 568226
rect -1572 568170 -1516 568226
rect -1448 568170 -1392 568226
rect -1820 568046 -1764 568102
rect -1696 568046 -1640 568102
rect -1572 568046 -1516 568102
rect -1448 568046 -1392 568102
rect -1820 567922 -1764 567978
rect -1696 567922 -1640 567978
rect -1572 567922 -1516 567978
rect -1448 567922 -1392 567978
rect -1820 550294 -1764 550350
rect -1696 550294 -1640 550350
rect -1572 550294 -1516 550350
rect -1448 550294 -1392 550350
rect -1820 550170 -1764 550226
rect -1696 550170 -1640 550226
rect -1572 550170 -1516 550226
rect -1448 550170 -1392 550226
rect -1820 550046 -1764 550102
rect -1696 550046 -1640 550102
rect -1572 550046 -1516 550102
rect -1448 550046 -1392 550102
rect -1820 549922 -1764 549978
rect -1696 549922 -1640 549978
rect -1572 549922 -1516 549978
rect -1448 549922 -1392 549978
rect -1820 532294 -1764 532350
rect -1696 532294 -1640 532350
rect -1572 532294 -1516 532350
rect -1448 532294 -1392 532350
rect -1820 532170 -1764 532226
rect -1696 532170 -1640 532226
rect -1572 532170 -1516 532226
rect -1448 532170 -1392 532226
rect -1820 532046 -1764 532102
rect -1696 532046 -1640 532102
rect -1572 532046 -1516 532102
rect -1448 532046 -1392 532102
rect -1820 531922 -1764 531978
rect -1696 531922 -1640 531978
rect -1572 531922 -1516 531978
rect -1448 531922 -1392 531978
rect -1820 514294 -1764 514350
rect -1696 514294 -1640 514350
rect -1572 514294 -1516 514350
rect -1448 514294 -1392 514350
rect -1820 514170 -1764 514226
rect -1696 514170 -1640 514226
rect -1572 514170 -1516 514226
rect -1448 514170 -1392 514226
rect -1820 514046 -1764 514102
rect -1696 514046 -1640 514102
rect -1572 514046 -1516 514102
rect -1448 514046 -1392 514102
rect -1820 513922 -1764 513978
rect -1696 513922 -1640 513978
rect -1572 513922 -1516 513978
rect -1448 513922 -1392 513978
rect -1820 496294 -1764 496350
rect -1696 496294 -1640 496350
rect -1572 496294 -1516 496350
rect -1448 496294 -1392 496350
rect -1820 496170 -1764 496226
rect -1696 496170 -1640 496226
rect -1572 496170 -1516 496226
rect -1448 496170 -1392 496226
rect -1820 496046 -1764 496102
rect -1696 496046 -1640 496102
rect -1572 496046 -1516 496102
rect -1448 496046 -1392 496102
rect -1820 495922 -1764 495978
rect -1696 495922 -1640 495978
rect -1572 495922 -1516 495978
rect -1448 495922 -1392 495978
rect -1820 478294 -1764 478350
rect -1696 478294 -1640 478350
rect -1572 478294 -1516 478350
rect -1448 478294 -1392 478350
rect -1820 478170 -1764 478226
rect -1696 478170 -1640 478226
rect -1572 478170 -1516 478226
rect -1448 478170 -1392 478226
rect -1820 478046 -1764 478102
rect -1696 478046 -1640 478102
rect -1572 478046 -1516 478102
rect -1448 478046 -1392 478102
rect -1820 477922 -1764 477978
rect -1696 477922 -1640 477978
rect -1572 477922 -1516 477978
rect -1448 477922 -1392 477978
rect -1820 460294 -1764 460350
rect -1696 460294 -1640 460350
rect -1572 460294 -1516 460350
rect -1448 460294 -1392 460350
rect -1820 460170 -1764 460226
rect -1696 460170 -1640 460226
rect -1572 460170 -1516 460226
rect -1448 460170 -1392 460226
rect -1820 460046 -1764 460102
rect -1696 460046 -1640 460102
rect -1572 460046 -1516 460102
rect -1448 460046 -1392 460102
rect -1820 459922 -1764 459978
rect -1696 459922 -1640 459978
rect -1572 459922 -1516 459978
rect -1448 459922 -1392 459978
rect -1820 442294 -1764 442350
rect -1696 442294 -1640 442350
rect -1572 442294 -1516 442350
rect -1448 442294 -1392 442350
rect -1820 442170 -1764 442226
rect -1696 442170 -1640 442226
rect -1572 442170 -1516 442226
rect -1448 442170 -1392 442226
rect -1820 442046 -1764 442102
rect -1696 442046 -1640 442102
rect -1572 442046 -1516 442102
rect -1448 442046 -1392 442102
rect -1820 441922 -1764 441978
rect -1696 441922 -1640 441978
rect -1572 441922 -1516 441978
rect -1448 441922 -1392 441978
rect -1820 424294 -1764 424350
rect -1696 424294 -1640 424350
rect -1572 424294 -1516 424350
rect -1448 424294 -1392 424350
rect -1820 424170 -1764 424226
rect -1696 424170 -1640 424226
rect -1572 424170 -1516 424226
rect -1448 424170 -1392 424226
rect -1820 424046 -1764 424102
rect -1696 424046 -1640 424102
rect -1572 424046 -1516 424102
rect -1448 424046 -1392 424102
rect -1820 423922 -1764 423978
rect -1696 423922 -1640 423978
rect -1572 423922 -1516 423978
rect -1448 423922 -1392 423978
rect -1820 406294 -1764 406350
rect -1696 406294 -1640 406350
rect -1572 406294 -1516 406350
rect -1448 406294 -1392 406350
rect -1820 406170 -1764 406226
rect -1696 406170 -1640 406226
rect -1572 406170 -1516 406226
rect -1448 406170 -1392 406226
rect -1820 406046 -1764 406102
rect -1696 406046 -1640 406102
rect -1572 406046 -1516 406102
rect -1448 406046 -1392 406102
rect -1820 405922 -1764 405978
rect -1696 405922 -1640 405978
rect -1572 405922 -1516 405978
rect -1448 405922 -1392 405978
rect -1820 388294 -1764 388350
rect -1696 388294 -1640 388350
rect -1572 388294 -1516 388350
rect -1448 388294 -1392 388350
rect -1820 388170 -1764 388226
rect -1696 388170 -1640 388226
rect -1572 388170 -1516 388226
rect -1448 388170 -1392 388226
rect -1820 388046 -1764 388102
rect -1696 388046 -1640 388102
rect -1572 388046 -1516 388102
rect -1448 388046 -1392 388102
rect -1820 387922 -1764 387978
rect -1696 387922 -1640 387978
rect -1572 387922 -1516 387978
rect -1448 387922 -1392 387978
rect -1820 370294 -1764 370350
rect -1696 370294 -1640 370350
rect -1572 370294 -1516 370350
rect -1448 370294 -1392 370350
rect -1820 370170 -1764 370226
rect -1696 370170 -1640 370226
rect -1572 370170 -1516 370226
rect -1448 370170 -1392 370226
rect -1820 370046 -1764 370102
rect -1696 370046 -1640 370102
rect -1572 370046 -1516 370102
rect -1448 370046 -1392 370102
rect -1820 369922 -1764 369978
rect -1696 369922 -1640 369978
rect -1572 369922 -1516 369978
rect -1448 369922 -1392 369978
rect -1820 352294 -1764 352350
rect -1696 352294 -1640 352350
rect -1572 352294 -1516 352350
rect -1448 352294 -1392 352350
rect -1820 352170 -1764 352226
rect -1696 352170 -1640 352226
rect -1572 352170 -1516 352226
rect -1448 352170 -1392 352226
rect -1820 352046 -1764 352102
rect -1696 352046 -1640 352102
rect -1572 352046 -1516 352102
rect -1448 352046 -1392 352102
rect -1820 351922 -1764 351978
rect -1696 351922 -1640 351978
rect -1572 351922 -1516 351978
rect -1448 351922 -1392 351978
rect -1820 334294 -1764 334350
rect -1696 334294 -1640 334350
rect -1572 334294 -1516 334350
rect -1448 334294 -1392 334350
rect -1820 334170 -1764 334226
rect -1696 334170 -1640 334226
rect -1572 334170 -1516 334226
rect -1448 334170 -1392 334226
rect -1820 334046 -1764 334102
rect -1696 334046 -1640 334102
rect -1572 334046 -1516 334102
rect -1448 334046 -1392 334102
rect -1820 333922 -1764 333978
rect -1696 333922 -1640 333978
rect -1572 333922 -1516 333978
rect -1448 333922 -1392 333978
rect -1820 316294 -1764 316350
rect -1696 316294 -1640 316350
rect -1572 316294 -1516 316350
rect -1448 316294 -1392 316350
rect -1820 316170 -1764 316226
rect -1696 316170 -1640 316226
rect -1572 316170 -1516 316226
rect -1448 316170 -1392 316226
rect -1820 316046 -1764 316102
rect -1696 316046 -1640 316102
rect -1572 316046 -1516 316102
rect -1448 316046 -1392 316102
rect -1820 315922 -1764 315978
rect -1696 315922 -1640 315978
rect -1572 315922 -1516 315978
rect -1448 315922 -1392 315978
rect -1820 298294 -1764 298350
rect -1696 298294 -1640 298350
rect -1572 298294 -1516 298350
rect -1448 298294 -1392 298350
rect -1820 298170 -1764 298226
rect -1696 298170 -1640 298226
rect -1572 298170 -1516 298226
rect -1448 298170 -1392 298226
rect -1820 298046 -1764 298102
rect -1696 298046 -1640 298102
rect -1572 298046 -1516 298102
rect -1448 298046 -1392 298102
rect -1820 297922 -1764 297978
rect -1696 297922 -1640 297978
rect -1572 297922 -1516 297978
rect -1448 297922 -1392 297978
rect -1820 280294 -1764 280350
rect -1696 280294 -1640 280350
rect -1572 280294 -1516 280350
rect -1448 280294 -1392 280350
rect -1820 280170 -1764 280226
rect -1696 280170 -1640 280226
rect -1572 280170 -1516 280226
rect -1448 280170 -1392 280226
rect -1820 280046 -1764 280102
rect -1696 280046 -1640 280102
rect -1572 280046 -1516 280102
rect -1448 280046 -1392 280102
rect -1820 279922 -1764 279978
rect -1696 279922 -1640 279978
rect -1572 279922 -1516 279978
rect -1448 279922 -1392 279978
rect -1820 262294 -1764 262350
rect -1696 262294 -1640 262350
rect -1572 262294 -1516 262350
rect -1448 262294 -1392 262350
rect -1820 262170 -1764 262226
rect -1696 262170 -1640 262226
rect -1572 262170 -1516 262226
rect -1448 262170 -1392 262226
rect -1820 262046 -1764 262102
rect -1696 262046 -1640 262102
rect -1572 262046 -1516 262102
rect -1448 262046 -1392 262102
rect -1820 261922 -1764 261978
rect -1696 261922 -1640 261978
rect -1572 261922 -1516 261978
rect -1448 261922 -1392 261978
rect -1820 244294 -1764 244350
rect -1696 244294 -1640 244350
rect -1572 244294 -1516 244350
rect -1448 244294 -1392 244350
rect -1820 244170 -1764 244226
rect -1696 244170 -1640 244226
rect -1572 244170 -1516 244226
rect -1448 244170 -1392 244226
rect -1820 244046 -1764 244102
rect -1696 244046 -1640 244102
rect -1572 244046 -1516 244102
rect -1448 244046 -1392 244102
rect -1820 243922 -1764 243978
rect -1696 243922 -1640 243978
rect -1572 243922 -1516 243978
rect -1448 243922 -1392 243978
rect -1820 226294 -1764 226350
rect -1696 226294 -1640 226350
rect -1572 226294 -1516 226350
rect -1448 226294 -1392 226350
rect -1820 226170 -1764 226226
rect -1696 226170 -1640 226226
rect -1572 226170 -1516 226226
rect -1448 226170 -1392 226226
rect -1820 226046 -1764 226102
rect -1696 226046 -1640 226102
rect -1572 226046 -1516 226102
rect -1448 226046 -1392 226102
rect -1820 225922 -1764 225978
rect -1696 225922 -1640 225978
rect -1572 225922 -1516 225978
rect -1448 225922 -1392 225978
rect -1820 208294 -1764 208350
rect -1696 208294 -1640 208350
rect -1572 208294 -1516 208350
rect -1448 208294 -1392 208350
rect -1820 208170 -1764 208226
rect -1696 208170 -1640 208226
rect -1572 208170 -1516 208226
rect -1448 208170 -1392 208226
rect -1820 208046 -1764 208102
rect -1696 208046 -1640 208102
rect -1572 208046 -1516 208102
rect -1448 208046 -1392 208102
rect -1820 207922 -1764 207978
rect -1696 207922 -1640 207978
rect -1572 207922 -1516 207978
rect -1448 207922 -1392 207978
rect -1820 190294 -1764 190350
rect -1696 190294 -1640 190350
rect -1572 190294 -1516 190350
rect -1448 190294 -1392 190350
rect -1820 190170 -1764 190226
rect -1696 190170 -1640 190226
rect -1572 190170 -1516 190226
rect -1448 190170 -1392 190226
rect -1820 190046 -1764 190102
rect -1696 190046 -1640 190102
rect -1572 190046 -1516 190102
rect -1448 190046 -1392 190102
rect -1820 189922 -1764 189978
rect -1696 189922 -1640 189978
rect -1572 189922 -1516 189978
rect -1448 189922 -1392 189978
rect -1820 172294 -1764 172350
rect -1696 172294 -1640 172350
rect -1572 172294 -1516 172350
rect -1448 172294 -1392 172350
rect -1820 172170 -1764 172226
rect -1696 172170 -1640 172226
rect -1572 172170 -1516 172226
rect -1448 172170 -1392 172226
rect -1820 172046 -1764 172102
rect -1696 172046 -1640 172102
rect -1572 172046 -1516 172102
rect -1448 172046 -1392 172102
rect -1820 171922 -1764 171978
rect -1696 171922 -1640 171978
rect -1572 171922 -1516 171978
rect -1448 171922 -1392 171978
rect -1820 154294 -1764 154350
rect -1696 154294 -1640 154350
rect -1572 154294 -1516 154350
rect -1448 154294 -1392 154350
rect -1820 154170 -1764 154226
rect -1696 154170 -1640 154226
rect -1572 154170 -1516 154226
rect -1448 154170 -1392 154226
rect -1820 154046 -1764 154102
rect -1696 154046 -1640 154102
rect -1572 154046 -1516 154102
rect -1448 154046 -1392 154102
rect -1820 153922 -1764 153978
rect -1696 153922 -1640 153978
rect -1572 153922 -1516 153978
rect -1448 153922 -1392 153978
rect -1820 136294 -1764 136350
rect -1696 136294 -1640 136350
rect -1572 136294 -1516 136350
rect -1448 136294 -1392 136350
rect -1820 136170 -1764 136226
rect -1696 136170 -1640 136226
rect -1572 136170 -1516 136226
rect -1448 136170 -1392 136226
rect -1820 136046 -1764 136102
rect -1696 136046 -1640 136102
rect -1572 136046 -1516 136102
rect -1448 136046 -1392 136102
rect -1820 135922 -1764 135978
rect -1696 135922 -1640 135978
rect -1572 135922 -1516 135978
rect -1448 135922 -1392 135978
rect -1820 118294 -1764 118350
rect -1696 118294 -1640 118350
rect -1572 118294 -1516 118350
rect -1448 118294 -1392 118350
rect -1820 118170 -1764 118226
rect -1696 118170 -1640 118226
rect -1572 118170 -1516 118226
rect -1448 118170 -1392 118226
rect -1820 118046 -1764 118102
rect -1696 118046 -1640 118102
rect -1572 118046 -1516 118102
rect -1448 118046 -1392 118102
rect -1820 117922 -1764 117978
rect -1696 117922 -1640 117978
rect -1572 117922 -1516 117978
rect -1448 117922 -1392 117978
rect -1820 100294 -1764 100350
rect -1696 100294 -1640 100350
rect -1572 100294 -1516 100350
rect -1448 100294 -1392 100350
rect -1820 100170 -1764 100226
rect -1696 100170 -1640 100226
rect -1572 100170 -1516 100226
rect -1448 100170 -1392 100226
rect -1820 100046 -1764 100102
rect -1696 100046 -1640 100102
rect -1572 100046 -1516 100102
rect -1448 100046 -1392 100102
rect -1820 99922 -1764 99978
rect -1696 99922 -1640 99978
rect -1572 99922 -1516 99978
rect -1448 99922 -1392 99978
rect -1820 82294 -1764 82350
rect -1696 82294 -1640 82350
rect -1572 82294 -1516 82350
rect -1448 82294 -1392 82350
rect -1820 82170 -1764 82226
rect -1696 82170 -1640 82226
rect -1572 82170 -1516 82226
rect -1448 82170 -1392 82226
rect -1820 82046 -1764 82102
rect -1696 82046 -1640 82102
rect -1572 82046 -1516 82102
rect -1448 82046 -1392 82102
rect -1820 81922 -1764 81978
rect -1696 81922 -1640 81978
rect -1572 81922 -1516 81978
rect -1448 81922 -1392 81978
rect -1820 64294 -1764 64350
rect -1696 64294 -1640 64350
rect -1572 64294 -1516 64350
rect -1448 64294 -1392 64350
rect -1820 64170 -1764 64226
rect -1696 64170 -1640 64226
rect -1572 64170 -1516 64226
rect -1448 64170 -1392 64226
rect -1820 64046 -1764 64102
rect -1696 64046 -1640 64102
rect -1572 64046 -1516 64102
rect -1448 64046 -1392 64102
rect -1820 63922 -1764 63978
rect -1696 63922 -1640 63978
rect -1572 63922 -1516 63978
rect -1448 63922 -1392 63978
rect -1820 46294 -1764 46350
rect -1696 46294 -1640 46350
rect -1572 46294 -1516 46350
rect -1448 46294 -1392 46350
rect -1820 46170 -1764 46226
rect -1696 46170 -1640 46226
rect -1572 46170 -1516 46226
rect -1448 46170 -1392 46226
rect -1820 46046 -1764 46102
rect -1696 46046 -1640 46102
rect -1572 46046 -1516 46102
rect -1448 46046 -1392 46102
rect -1820 45922 -1764 45978
rect -1696 45922 -1640 45978
rect -1572 45922 -1516 45978
rect -1448 45922 -1392 45978
rect -1820 28294 -1764 28350
rect -1696 28294 -1640 28350
rect -1572 28294 -1516 28350
rect -1448 28294 -1392 28350
rect -1820 28170 -1764 28226
rect -1696 28170 -1640 28226
rect -1572 28170 -1516 28226
rect -1448 28170 -1392 28226
rect -1820 28046 -1764 28102
rect -1696 28046 -1640 28102
rect -1572 28046 -1516 28102
rect -1448 28046 -1392 28102
rect -1820 27922 -1764 27978
rect -1696 27922 -1640 27978
rect -1572 27922 -1516 27978
rect -1448 27922 -1392 27978
rect -1820 10294 -1764 10350
rect -1696 10294 -1640 10350
rect -1572 10294 -1516 10350
rect -1448 10294 -1392 10350
rect -1820 10170 -1764 10226
rect -1696 10170 -1640 10226
rect -1572 10170 -1516 10226
rect -1448 10170 -1392 10226
rect -1820 10046 -1764 10102
rect -1696 10046 -1640 10102
rect -1572 10046 -1516 10102
rect -1448 10046 -1392 10102
rect -1820 9922 -1764 9978
rect -1696 9922 -1640 9978
rect -1572 9922 -1516 9978
rect -1448 9922 -1392 9978
rect -860 597156 -804 597212
rect -736 597156 -680 597212
rect -612 597156 -556 597212
rect -488 597156 -432 597212
rect -860 597032 -804 597088
rect -736 597032 -680 597088
rect -612 597032 -556 597088
rect -488 597032 -432 597088
rect -860 596908 -804 596964
rect -736 596908 -680 596964
rect -612 596908 -556 596964
rect -488 596908 -432 596964
rect -860 596784 -804 596840
rect -736 596784 -680 596840
rect -612 596784 -556 596840
rect -488 596784 -432 596840
rect -860 580294 -804 580350
rect -736 580294 -680 580350
rect -612 580294 -556 580350
rect -488 580294 -432 580350
rect -860 580170 -804 580226
rect -736 580170 -680 580226
rect -612 580170 -556 580226
rect -488 580170 -432 580226
rect -860 580046 -804 580102
rect -736 580046 -680 580102
rect -612 580046 -556 580102
rect -488 580046 -432 580102
rect -860 579922 -804 579978
rect -736 579922 -680 579978
rect -612 579922 -556 579978
rect -488 579922 -432 579978
rect -860 562294 -804 562350
rect -736 562294 -680 562350
rect -612 562294 -556 562350
rect -488 562294 -432 562350
rect -860 562170 -804 562226
rect -736 562170 -680 562226
rect -612 562170 -556 562226
rect -488 562170 -432 562226
rect -860 562046 -804 562102
rect -736 562046 -680 562102
rect -612 562046 -556 562102
rect -488 562046 -432 562102
rect -860 561922 -804 561978
rect -736 561922 -680 561978
rect -612 561922 -556 561978
rect -488 561922 -432 561978
rect 5514 597156 5570 597212
rect 5638 597156 5694 597212
rect 5762 597156 5818 597212
rect 5886 597156 5942 597212
rect 5514 597032 5570 597088
rect 5638 597032 5694 597088
rect 5762 597032 5818 597088
rect 5886 597032 5942 597088
rect 5514 596908 5570 596964
rect 5638 596908 5694 596964
rect 5762 596908 5818 596964
rect 5886 596908 5942 596964
rect 5514 596784 5570 596840
rect 5638 596784 5694 596840
rect 5762 596784 5818 596840
rect 5886 596784 5942 596840
rect 5514 580294 5570 580350
rect 5638 580294 5694 580350
rect 5762 580294 5818 580350
rect 5886 580294 5942 580350
rect 5514 580170 5570 580226
rect 5638 580170 5694 580226
rect 5762 580170 5818 580226
rect 5886 580170 5942 580226
rect 5514 580046 5570 580102
rect 5638 580046 5694 580102
rect 5762 580046 5818 580102
rect 5886 580046 5942 580102
rect 5514 579922 5570 579978
rect 5638 579922 5694 579978
rect 5762 579922 5818 579978
rect 5886 579922 5942 579978
rect 5514 562294 5570 562350
rect 5638 562294 5694 562350
rect 5762 562294 5818 562350
rect 5886 562294 5942 562350
rect 5514 562170 5570 562226
rect 5638 562170 5694 562226
rect 5762 562170 5818 562226
rect 5886 562170 5942 562226
rect 5514 562046 5570 562102
rect 5638 562046 5694 562102
rect 5762 562046 5818 562102
rect 5886 562046 5942 562102
rect 5514 561922 5570 561978
rect 5638 561922 5694 561978
rect 5762 561922 5818 561978
rect 5886 561922 5942 561978
rect -860 544294 -804 544350
rect -736 544294 -680 544350
rect -612 544294 -556 544350
rect -488 544294 -432 544350
rect -860 544170 -804 544226
rect -736 544170 -680 544226
rect -612 544170 -556 544226
rect -488 544170 -432 544226
rect -860 544046 -804 544102
rect -736 544046 -680 544102
rect -612 544046 -556 544102
rect -488 544046 -432 544102
rect -860 543922 -804 543978
rect -736 543922 -680 543978
rect -612 543922 -556 543978
rect -488 543922 -432 543978
rect -860 526294 -804 526350
rect -736 526294 -680 526350
rect -612 526294 -556 526350
rect -488 526294 -432 526350
rect -860 526170 -804 526226
rect -736 526170 -680 526226
rect -612 526170 -556 526226
rect -488 526170 -432 526226
rect -860 526046 -804 526102
rect -736 526046 -680 526102
rect -612 526046 -556 526102
rect -488 526046 -432 526102
rect -860 525922 -804 525978
rect -736 525922 -680 525978
rect -612 525922 -556 525978
rect -488 525922 -432 525978
rect -860 508294 -804 508350
rect -736 508294 -680 508350
rect -612 508294 -556 508350
rect -488 508294 -432 508350
rect -860 508170 -804 508226
rect -736 508170 -680 508226
rect -612 508170 -556 508226
rect -488 508170 -432 508226
rect -860 508046 -804 508102
rect -736 508046 -680 508102
rect -612 508046 -556 508102
rect -488 508046 -432 508102
rect -860 507922 -804 507978
rect -736 507922 -680 507978
rect -612 507922 -556 507978
rect -488 507922 -432 507978
rect -860 490294 -804 490350
rect -736 490294 -680 490350
rect -612 490294 -556 490350
rect -488 490294 -432 490350
rect -860 490170 -804 490226
rect -736 490170 -680 490226
rect -612 490170 -556 490226
rect -488 490170 -432 490226
rect -860 490046 -804 490102
rect -736 490046 -680 490102
rect -612 490046 -556 490102
rect -488 490046 -432 490102
rect -860 489922 -804 489978
rect -736 489922 -680 489978
rect -612 489922 -556 489978
rect -488 489922 -432 489978
rect 9234 598116 9290 598172
rect 9358 598116 9414 598172
rect 9482 598116 9538 598172
rect 9606 598116 9662 598172
rect 9234 597992 9290 598048
rect 9358 597992 9414 598048
rect 9482 597992 9538 598048
rect 9606 597992 9662 598048
rect 9234 597868 9290 597924
rect 9358 597868 9414 597924
rect 9482 597868 9538 597924
rect 9606 597868 9662 597924
rect 9234 597744 9290 597800
rect 9358 597744 9414 597800
rect 9482 597744 9538 597800
rect 9606 597744 9662 597800
rect 9234 586294 9290 586350
rect 9358 586294 9414 586350
rect 9482 586294 9538 586350
rect 9606 586294 9662 586350
rect 9234 586170 9290 586226
rect 9358 586170 9414 586226
rect 9482 586170 9538 586226
rect 9606 586170 9662 586226
rect 9234 586046 9290 586102
rect 9358 586046 9414 586102
rect 9482 586046 9538 586102
rect 9606 586046 9662 586102
rect 9234 585922 9290 585978
rect 9358 585922 9414 585978
rect 9482 585922 9538 585978
rect 9606 585922 9662 585978
rect 9234 568294 9290 568350
rect 9358 568294 9414 568350
rect 9482 568294 9538 568350
rect 9606 568294 9662 568350
rect 9234 568170 9290 568226
rect 9358 568170 9414 568226
rect 9482 568170 9538 568226
rect 9606 568170 9662 568226
rect 9234 568046 9290 568102
rect 9358 568046 9414 568102
rect 9482 568046 9538 568102
rect 9606 568046 9662 568102
rect 9234 567922 9290 567978
rect 9358 567922 9414 567978
rect 9482 567922 9538 567978
rect 9606 567922 9662 567978
rect 9234 550294 9290 550350
rect 9358 550294 9414 550350
rect 9482 550294 9538 550350
rect 9606 550294 9662 550350
rect 9234 550170 9290 550226
rect 9358 550170 9414 550226
rect 9482 550170 9538 550226
rect 9606 550170 9662 550226
rect 9234 550046 9290 550102
rect 9358 550046 9414 550102
rect 9482 550046 9538 550102
rect 9606 550046 9662 550102
rect 9234 549922 9290 549978
rect 9358 549922 9414 549978
rect 9482 549922 9538 549978
rect 9606 549922 9662 549978
rect 5514 544294 5570 544350
rect 5638 544294 5694 544350
rect 5762 544294 5818 544350
rect 5886 544294 5942 544350
rect 5514 544170 5570 544226
rect 5638 544170 5694 544226
rect 5762 544170 5818 544226
rect 5886 544170 5942 544226
rect 5514 544046 5570 544102
rect 5638 544046 5694 544102
rect 5762 544046 5818 544102
rect 5886 544046 5942 544102
rect 5514 543922 5570 543978
rect 5638 543922 5694 543978
rect 5762 543922 5818 543978
rect 5886 543922 5942 543978
rect 5514 526294 5570 526350
rect 5638 526294 5694 526350
rect 5762 526294 5818 526350
rect 5886 526294 5942 526350
rect 5514 526170 5570 526226
rect 5638 526170 5694 526226
rect 5762 526170 5818 526226
rect 5886 526170 5942 526226
rect 5514 526046 5570 526102
rect 5638 526046 5694 526102
rect 5762 526046 5818 526102
rect 5886 526046 5942 526102
rect 5514 525922 5570 525978
rect 5638 525922 5694 525978
rect 5762 525922 5818 525978
rect 5886 525922 5942 525978
rect -860 472294 -804 472350
rect -736 472294 -680 472350
rect -612 472294 -556 472350
rect -488 472294 -432 472350
rect -860 472170 -804 472226
rect -736 472170 -680 472226
rect -612 472170 -556 472226
rect -488 472170 -432 472226
rect -860 472046 -804 472102
rect -736 472046 -680 472102
rect -612 472046 -556 472102
rect -488 472046 -432 472102
rect -860 471922 -804 471978
rect -736 471922 -680 471978
rect -612 471922 -556 471978
rect -488 471922 -432 471978
rect 5514 508294 5570 508350
rect 5638 508294 5694 508350
rect 5762 508294 5818 508350
rect 5886 508294 5942 508350
rect 5514 508170 5570 508226
rect 5638 508170 5694 508226
rect 5762 508170 5818 508226
rect 5886 508170 5942 508226
rect 5514 508046 5570 508102
rect 5638 508046 5694 508102
rect 5762 508046 5818 508102
rect 5886 508046 5942 508102
rect 5514 507922 5570 507978
rect 5638 507922 5694 507978
rect 5762 507922 5818 507978
rect 5886 507922 5942 507978
rect 5514 490294 5570 490350
rect 5638 490294 5694 490350
rect 5762 490294 5818 490350
rect 5886 490294 5942 490350
rect 5514 490170 5570 490226
rect 5638 490170 5694 490226
rect 5762 490170 5818 490226
rect 5886 490170 5942 490226
rect 5514 490046 5570 490102
rect 5638 490046 5694 490102
rect 5762 490046 5818 490102
rect 5886 490046 5942 490102
rect 5514 489922 5570 489978
rect 5638 489922 5694 489978
rect 5762 489922 5818 489978
rect 5886 489922 5942 489978
rect 5514 472294 5570 472350
rect 5638 472294 5694 472350
rect 5762 472294 5818 472350
rect 5886 472294 5942 472350
rect 5514 472170 5570 472226
rect 5638 472170 5694 472226
rect 5762 472170 5818 472226
rect 5886 472170 5942 472226
rect 5514 472046 5570 472102
rect 5638 472046 5694 472102
rect 5762 472046 5818 472102
rect 5886 472046 5942 472102
rect 5514 471922 5570 471978
rect 5638 471922 5694 471978
rect 5762 471922 5818 471978
rect 5886 471922 5942 471978
rect -860 454294 -804 454350
rect -736 454294 -680 454350
rect -612 454294 -556 454350
rect -488 454294 -432 454350
rect -860 454170 -804 454226
rect -736 454170 -680 454226
rect -612 454170 -556 454226
rect -488 454170 -432 454226
rect -860 454046 -804 454102
rect -736 454046 -680 454102
rect -612 454046 -556 454102
rect -488 454046 -432 454102
rect -860 453922 -804 453978
rect -736 453922 -680 453978
rect -612 453922 -556 453978
rect -488 453922 -432 453978
rect -860 436294 -804 436350
rect -736 436294 -680 436350
rect -612 436294 -556 436350
rect -488 436294 -432 436350
rect -860 436170 -804 436226
rect -736 436170 -680 436226
rect -612 436170 -556 436226
rect -488 436170 -432 436226
rect -860 436046 -804 436102
rect -736 436046 -680 436102
rect -612 436046 -556 436102
rect -488 436046 -432 436102
rect -860 435922 -804 435978
rect -736 435922 -680 435978
rect -612 435922 -556 435978
rect -488 435922 -432 435978
rect -860 418294 -804 418350
rect -736 418294 -680 418350
rect -612 418294 -556 418350
rect -488 418294 -432 418350
rect -860 418170 -804 418226
rect -736 418170 -680 418226
rect -612 418170 -556 418226
rect -488 418170 -432 418226
rect -860 418046 -804 418102
rect -736 418046 -680 418102
rect -612 418046 -556 418102
rect -488 418046 -432 418102
rect -860 417922 -804 417978
rect -736 417922 -680 417978
rect -612 417922 -556 417978
rect -488 417922 -432 417978
rect -860 400294 -804 400350
rect -736 400294 -680 400350
rect -612 400294 -556 400350
rect -488 400294 -432 400350
rect -860 400170 -804 400226
rect -736 400170 -680 400226
rect -612 400170 -556 400226
rect -488 400170 -432 400226
rect -860 400046 -804 400102
rect -736 400046 -680 400102
rect -612 400046 -556 400102
rect -488 400046 -432 400102
rect -860 399922 -804 399978
rect -736 399922 -680 399978
rect -612 399922 -556 399978
rect -488 399922 -432 399978
rect 5514 454294 5570 454350
rect 5638 454294 5694 454350
rect 5762 454294 5818 454350
rect 5886 454294 5942 454350
rect 5514 454170 5570 454226
rect 5638 454170 5694 454226
rect 5762 454170 5818 454226
rect 5886 454170 5942 454226
rect 5514 454046 5570 454102
rect 5638 454046 5694 454102
rect 5762 454046 5818 454102
rect 5886 454046 5942 454102
rect 5514 453922 5570 453978
rect 5638 453922 5694 453978
rect 5762 453922 5818 453978
rect 5886 453922 5942 453978
rect 5514 436294 5570 436350
rect 5638 436294 5694 436350
rect 5762 436294 5818 436350
rect 5886 436294 5942 436350
rect 5514 436170 5570 436226
rect 5638 436170 5694 436226
rect 5762 436170 5818 436226
rect 5886 436170 5942 436226
rect 5514 436046 5570 436102
rect 5638 436046 5694 436102
rect 5762 436046 5818 436102
rect 5886 436046 5942 436102
rect 5514 435922 5570 435978
rect 5638 435922 5694 435978
rect 5762 435922 5818 435978
rect 5886 435922 5942 435978
rect 5514 418294 5570 418350
rect 5638 418294 5694 418350
rect 5762 418294 5818 418350
rect 5886 418294 5942 418350
rect 5514 418170 5570 418226
rect 5638 418170 5694 418226
rect 5762 418170 5818 418226
rect 5886 418170 5942 418226
rect 5514 418046 5570 418102
rect 5638 418046 5694 418102
rect 5762 418046 5818 418102
rect 5886 418046 5942 418102
rect 5514 417922 5570 417978
rect 5638 417922 5694 417978
rect 5762 417922 5818 417978
rect 5886 417922 5942 417978
rect 7532 409022 7588 409078
rect 9234 532294 9290 532350
rect 9358 532294 9414 532350
rect 9482 532294 9538 532350
rect 9606 532294 9662 532350
rect 9234 532170 9290 532226
rect 9358 532170 9414 532226
rect 9482 532170 9538 532226
rect 9606 532170 9662 532226
rect 9234 532046 9290 532102
rect 9358 532046 9414 532102
rect 9482 532046 9538 532102
rect 9606 532046 9662 532102
rect 9234 531922 9290 531978
rect 9358 531922 9414 531978
rect 9482 531922 9538 531978
rect 9606 531922 9662 531978
rect 9234 514294 9290 514350
rect 9358 514294 9414 514350
rect 9482 514294 9538 514350
rect 9606 514294 9662 514350
rect 9234 514170 9290 514226
rect 9358 514170 9414 514226
rect 9482 514170 9538 514226
rect 9606 514170 9662 514226
rect 9234 514046 9290 514102
rect 9358 514046 9414 514102
rect 9482 514046 9538 514102
rect 9606 514046 9662 514102
rect 9234 513922 9290 513978
rect 9358 513922 9414 513978
rect 9482 513922 9538 513978
rect 9606 513922 9662 513978
rect 9234 496294 9290 496350
rect 9358 496294 9414 496350
rect 9482 496294 9538 496350
rect 9606 496294 9662 496350
rect 9234 496170 9290 496226
rect 9358 496170 9414 496226
rect 9482 496170 9538 496226
rect 9606 496170 9662 496226
rect 9234 496046 9290 496102
rect 9358 496046 9414 496102
rect 9482 496046 9538 496102
rect 9606 496046 9662 496102
rect 9234 495922 9290 495978
rect 9358 495922 9414 495978
rect 9482 495922 9538 495978
rect 9606 495922 9662 495978
rect 9234 478294 9290 478350
rect 9358 478294 9414 478350
rect 9482 478294 9538 478350
rect 9606 478294 9662 478350
rect 9234 478170 9290 478226
rect 9358 478170 9414 478226
rect 9482 478170 9538 478226
rect 9606 478170 9662 478226
rect 9234 478046 9290 478102
rect 9358 478046 9414 478102
rect 9482 478046 9538 478102
rect 9606 478046 9662 478102
rect 9234 477922 9290 477978
rect 9358 477922 9414 477978
rect 9482 477922 9538 477978
rect 9606 477922 9662 477978
rect 9234 460294 9290 460350
rect 9358 460294 9414 460350
rect 9482 460294 9538 460350
rect 9606 460294 9662 460350
rect 9234 460170 9290 460226
rect 9358 460170 9414 460226
rect 9482 460170 9538 460226
rect 9606 460170 9662 460226
rect 9234 460046 9290 460102
rect 9358 460046 9414 460102
rect 9482 460046 9538 460102
rect 9606 460046 9662 460102
rect 9234 459922 9290 459978
rect 9358 459922 9414 459978
rect 9482 459922 9538 459978
rect 9606 459922 9662 459978
rect 9234 442294 9290 442350
rect 9358 442294 9414 442350
rect 9482 442294 9538 442350
rect 9606 442294 9662 442350
rect 9234 442170 9290 442226
rect 9358 442170 9414 442226
rect 9482 442170 9538 442226
rect 9606 442170 9662 442226
rect 9234 442046 9290 442102
rect 9358 442046 9414 442102
rect 9482 442046 9538 442102
rect 9606 442046 9662 442102
rect 9234 441922 9290 441978
rect 9358 441922 9414 441978
rect 9482 441922 9538 441978
rect 9606 441922 9662 441978
rect 9234 424294 9290 424350
rect 9358 424294 9414 424350
rect 9482 424294 9538 424350
rect 9606 424294 9662 424350
rect 9234 424170 9290 424226
rect 9358 424170 9414 424226
rect 9482 424170 9538 424226
rect 9606 424170 9662 424226
rect 9234 424046 9290 424102
rect 9358 424046 9414 424102
rect 9482 424046 9538 424102
rect 9606 424046 9662 424102
rect 9234 423922 9290 423978
rect 9358 423922 9414 423978
rect 9482 423922 9538 423978
rect 9606 423922 9662 423978
rect 5514 400294 5570 400350
rect 5638 400294 5694 400350
rect 5762 400294 5818 400350
rect 5886 400294 5942 400350
rect 5514 400170 5570 400226
rect 5638 400170 5694 400226
rect 5762 400170 5818 400226
rect 5886 400170 5942 400226
rect 5514 400046 5570 400102
rect 5638 400046 5694 400102
rect 5762 400046 5818 400102
rect 5886 400046 5942 400102
rect 5514 399922 5570 399978
rect 5638 399922 5694 399978
rect 5762 399922 5818 399978
rect 5886 399922 5942 399978
rect -860 382294 -804 382350
rect -736 382294 -680 382350
rect -612 382294 -556 382350
rect -488 382294 -432 382350
rect -860 382170 -804 382226
rect -736 382170 -680 382226
rect -612 382170 -556 382226
rect -488 382170 -432 382226
rect -860 382046 -804 382102
rect -736 382046 -680 382102
rect -612 382046 -556 382102
rect -488 382046 -432 382102
rect -860 381922 -804 381978
rect -736 381922 -680 381978
rect -612 381922 -556 381978
rect -488 381922 -432 381978
rect 9234 406294 9290 406350
rect 9358 406294 9414 406350
rect 9482 406294 9538 406350
rect 9606 406294 9662 406350
rect 9234 406170 9290 406226
rect 9358 406170 9414 406226
rect 9482 406170 9538 406226
rect 9606 406170 9662 406226
rect 9234 406046 9290 406102
rect 9358 406046 9414 406102
rect 9482 406046 9538 406102
rect 9606 406046 9662 406102
rect 9234 405922 9290 405978
rect 9358 405922 9414 405978
rect 9482 405922 9538 405978
rect 9606 405922 9662 405978
rect 9234 388294 9290 388350
rect 9358 388294 9414 388350
rect 9482 388294 9538 388350
rect 9606 388294 9662 388350
rect 9234 388170 9290 388226
rect 9358 388170 9414 388226
rect 9482 388170 9538 388226
rect 9606 388170 9662 388226
rect 9234 388046 9290 388102
rect 9358 388046 9414 388102
rect 9482 388046 9538 388102
rect 9606 388046 9662 388102
rect 9234 387922 9290 387978
rect 9358 387922 9414 387978
rect 9482 387922 9538 387978
rect 9606 387922 9662 387978
rect 5514 382294 5570 382350
rect 5638 382294 5694 382350
rect 5762 382294 5818 382350
rect 5886 382294 5942 382350
rect 5514 382170 5570 382226
rect 5638 382170 5694 382226
rect 5762 382170 5818 382226
rect 5886 382170 5942 382226
rect 5514 382046 5570 382102
rect 5638 382046 5694 382102
rect 5762 382046 5818 382102
rect 5886 382046 5942 382102
rect 5514 381922 5570 381978
rect 5638 381922 5694 381978
rect 5762 381922 5818 381978
rect 5886 381922 5942 381978
rect -860 364294 -804 364350
rect -736 364294 -680 364350
rect -612 364294 -556 364350
rect -488 364294 -432 364350
rect -860 364170 -804 364226
rect -736 364170 -680 364226
rect -612 364170 -556 364226
rect -488 364170 -432 364226
rect -860 364046 -804 364102
rect -736 364046 -680 364102
rect -612 364046 -556 364102
rect -488 364046 -432 364102
rect -860 363922 -804 363978
rect -736 363922 -680 363978
rect -612 363922 -556 363978
rect -488 363922 -432 363978
rect 5514 364294 5570 364350
rect 5638 364294 5694 364350
rect 5762 364294 5818 364350
rect 5886 364294 5942 364350
rect 5514 364170 5570 364226
rect 5638 364170 5694 364226
rect 5762 364170 5818 364226
rect 5886 364170 5942 364226
rect 5514 364046 5570 364102
rect 5638 364046 5694 364102
rect 5762 364046 5818 364102
rect 5886 364046 5942 364102
rect 5514 363922 5570 363978
rect 5638 363922 5694 363978
rect 5762 363922 5818 363978
rect 5886 363922 5942 363978
rect -860 346294 -804 346350
rect -736 346294 -680 346350
rect -612 346294 -556 346350
rect -488 346294 -432 346350
rect -860 346170 -804 346226
rect -736 346170 -680 346226
rect -612 346170 -556 346226
rect -488 346170 -432 346226
rect -860 346046 -804 346102
rect -736 346046 -680 346102
rect -612 346046 -556 346102
rect -488 346046 -432 346102
rect -860 345922 -804 345978
rect -736 345922 -680 345978
rect -612 345922 -556 345978
rect -488 345922 -432 345978
rect 5514 346294 5570 346350
rect 5638 346294 5694 346350
rect 5762 346294 5818 346350
rect 5886 346294 5942 346350
rect 5514 346170 5570 346226
rect 5638 346170 5694 346226
rect 5762 346170 5818 346226
rect 5886 346170 5942 346226
rect 5514 346046 5570 346102
rect 5638 346046 5694 346102
rect 5762 346046 5818 346102
rect 5886 346046 5942 346102
rect 5514 345922 5570 345978
rect 5638 345922 5694 345978
rect 5762 345922 5818 345978
rect 5886 345922 5942 345978
rect -860 328294 -804 328350
rect -736 328294 -680 328350
rect -612 328294 -556 328350
rect -488 328294 -432 328350
rect -860 328170 -804 328226
rect -736 328170 -680 328226
rect -612 328170 -556 328226
rect -488 328170 -432 328226
rect -860 328046 -804 328102
rect -736 328046 -680 328102
rect -612 328046 -556 328102
rect -488 328046 -432 328102
rect -860 327922 -804 327978
rect -736 327922 -680 327978
rect -612 327922 -556 327978
rect -488 327922 -432 327978
rect -860 310294 -804 310350
rect -736 310294 -680 310350
rect -612 310294 -556 310350
rect -488 310294 -432 310350
rect -860 310170 -804 310226
rect -736 310170 -680 310226
rect -612 310170 -556 310226
rect -488 310170 -432 310226
rect -860 310046 -804 310102
rect -736 310046 -680 310102
rect -612 310046 -556 310102
rect -488 310046 -432 310102
rect -860 309922 -804 309978
rect -736 309922 -680 309978
rect -612 309922 -556 309978
rect -488 309922 -432 309978
rect 5514 328294 5570 328350
rect 5638 328294 5694 328350
rect 5762 328294 5818 328350
rect 5886 328294 5942 328350
rect 5514 328170 5570 328226
rect 5638 328170 5694 328226
rect 5762 328170 5818 328226
rect 5886 328170 5942 328226
rect 5514 328046 5570 328102
rect 5638 328046 5694 328102
rect 5762 328046 5818 328102
rect 5886 328046 5942 328102
rect 5514 327922 5570 327978
rect 5638 327922 5694 327978
rect 5762 327922 5818 327978
rect 5886 327922 5942 327978
rect 5514 310294 5570 310350
rect 5638 310294 5694 310350
rect 5762 310294 5818 310350
rect 5886 310294 5942 310350
rect 5514 310170 5570 310226
rect 5638 310170 5694 310226
rect 5762 310170 5818 310226
rect 5886 310170 5942 310226
rect 5514 310046 5570 310102
rect 5638 310046 5694 310102
rect 5762 310046 5818 310102
rect 5886 310046 5942 310102
rect 5514 309922 5570 309978
rect 5638 309922 5694 309978
rect 5762 309922 5818 309978
rect 5886 309922 5942 309978
rect -860 292294 -804 292350
rect -736 292294 -680 292350
rect -612 292294 -556 292350
rect -488 292294 -432 292350
rect -860 292170 -804 292226
rect -736 292170 -680 292226
rect -612 292170 -556 292226
rect -488 292170 -432 292226
rect -860 292046 -804 292102
rect -736 292046 -680 292102
rect -612 292046 -556 292102
rect -488 292046 -432 292102
rect -860 291922 -804 291978
rect -736 291922 -680 291978
rect -612 291922 -556 291978
rect -488 291922 -432 291978
rect -860 274294 -804 274350
rect -736 274294 -680 274350
rect -612 274294 -556 274350
rect -488 274294 -432 274350
rect -860 274170 -804 274226
rect -736 274170 -680 274226
rect -612 274170 -556 274226
rect -488 274170 -432 274226
rect -860 274046 -804 274102
rect -736 274046 -680 274102
rect -612 274046 -556 274102
rect -488 274046 -432 274102
rect -860 273922 -804 273978
rect -736 273922 -680 273978
rect -612 273922 -556 273978
rect -488 273922 -432 273978
rect -860 256294 -804 256350
rect -736 256294 -680 256350
rect -612 256294 -556 256350
rect -488 256294 -432 256350
rect -860 256170 -804 256226
rect -736 256170 -680 256226
rect -612 256170 -556 256226
rect -488 256170 -432 256226
rect -860 256046 -804 256102
rect -736 256046 -680 256102
rect -612 256046 -556 256102
rect -488 256046 -432 256102
rect -860 255922 -804 255978
rect -736 255922 -680 255978
rect -612 255922 -556 255978
rect -488 255922 -432 255978
rect 4060 247022 4116 247078
rect -860 238294 -804 238350
rect -736 238294 -680 238350
rect -612 238294 -556 238350
rect -488 238294 -432 238350
rect -860 238170 -804 238226
rect -736 238170 -680 238226
rect -612 238170 -556 238226
rect -488 238170 -432 238226
rect -860 238046 -804 238102
rect -736 238046 -680 238102
rect -612 238046 -556 238102
rect -488 238046 -432 238102
rect -860 237922 -804 237978
rect -736 237922 -680 237978
rect -612 237922 -556 237978
rect -488 237922 -432 237978
rect -860 220294 -804 220350
rect -736 220294 -680 220350
rect -612 220294 -556 220350
rect -488 220294 -432 220350
rect -860 220170 -804 220226
rect -736 220170 -680 220226
rect -612 220170 -556 220226
rect -488 220170 -432 220226
rect -860 220046 -804 220102
rect -736 220046 -680 220102
rect -612 220046 -556 220102
rect -488 220046 -432 220102
rect -860 219922 -804 219978
rect -736 219922 -680 219978
rect -612 219922 -556 219978
rect -488 219922 -432 219978
rect -860 202294 -804 202350
rect -736 202294 -680 202350
rect -612 202294 -556 202350
rect -488 202294 -432 202350
rect -860 202170 -804 202226
rect -736 202170 -680 202226
rect -612 202170 -556 202226
rect -488 202170 -432 202226
rect -860 202046 -804 202102
rect -736 202046 -680 202102
rect -612 202046 -556 202102
rect -488 202046 -432 202102
rect -860 201922 -804 201978
rect -736 201922 -680 201978
rect -612 201922 -556 201978
rect -488 201922 -432 201978
rect 4172 206522 4228 206578
rect -860 184294 -804 184350
rect -736 184294 -680 184350
rect -612 184294 -556 184350
rect -488 184294 -432 184350
rect -860 184170 -804 184226
rect -736 184170 -680 184226
rect -612 184170 -556 184226
rect -488 184170 -432 184226
rect -860 184046 -804 184102
rect -736 184046 -680 184102
rect -612 184046 -556 184102
rect -488 184046 -432 184102
rect -860 183922 -804 183978
rect -736 183922 -680 183978
rect -612 183922 -556 183978
rect -488 183922 -432 183978
rect -860 166294 -804 166350
rect -736 166294 -680 166350
rect -612 166294 -556 166350
rect -488 166294 -432 166350
rect -860 166170 -804 166226
rect -736 166170 -680 166226
rect -612 166170 -556 166226
rect -488 166170 -432 166226
rect -860 166046 -804 166102
rect -736 166046 -680 166102
rect -612 166046 -556 166102
rect -488 166046 -432 166102
rect -860 165922 -804 165978
rect -736 165922 -680 165978
rect -612 165922 -556 165978
rect -488 165922 -432 165978
rect 4172 164582 4228 164638
rect -860 148294 -804 148350
rect -736 148294 -680 148350
rect -612 148294 -556 148350
rect -488 148294 -432 148350
rect -860 148170 -804 148226
rect -736 148170 -680 148226
rect -612 148170 -556 148226
rect -488 148170 -432 148226
rect -860 148046 -804 148102
rect -736 148046 -680 148102
rect -612 148046 -556 148102
rect -488 148046 -432 148102
rect -860 147922 -804 147978
rect -736 147922 -680 147978
rect -612 147922 -556 147978
rect -488 147922 -432 147978
rect -860 130294 -804 130350
rect -736 130294 -680 130350
rect -612 130294 -556 130350
rect -488 130294 -432 130350
rect -860 130170 -804 130226
rect -736 130170 -680 130226
rect -612 130170 -556 130226
rect -488 130170 -432 130226
rect -860 130046 -804 130102
rect -736 130046 -680 130102
rect -612 130046 -556 130102
rect -488 130046 -432 130102
rect -860 129922 -804 129978
rect -736 129922 -680 129978
rect -612 129922 -556 129978
rect -488 129922 -432 129978
rect -860 112294 -804 112350
rect -736 112294 -680 112350
rect -612 112294 -556 112350
rect -488 112294 -432 112350
rect -860 112170 -804 112226
rect -736 112170 -680 112226
rect -612 112170 -556 112226
rect -488 112170 -432 112226
rect -860 112046 -804 112102
rect -736 112046 -680 112102
rect -612 112046 -556 112102
rect -488 112046 -432 112102
rect -860 111922 -804 111978
rect -736 111922 -680 111978
rect -612 111922 -556 111978
rect -488 111922 -432 111978
rect -860 94294 -804 94350
rect -736 94294 -680 94350
rect -612 94294 -556 94350
rect -488 94294 -432 94350
rect -860 94170 -804 94226
rect -736 94170 -680 94226
rect -612 94170 -556 94226
rect -488 94170 -432 94226
rect -860 94046 -804 94102
rect -736 94046 -680 94102
rect -612 94046 -556 94102
rect -488 94046 -432 94102
rect -860 93922 -804 93978
rect -736 93922 -680 93978
rect -612 93922 -556 93978
rect -488 93922 -432 93978
rect -860 76294 -804 76350
rect -736 76294 -680 76350
rect -612 76294 -556 76350
rect -488 76294 -432 76350
rect -860 76170 -804 76226
rect -736 76170 -680 76226
rect -612 76170 -556 76226
rect -488 76170 -432 76226
rect -860 76046 -804 76102
rect -736 76046 -680 76102
rect -612 76046 -556 76102
rect -488 76046 -432 76102
rect -860 75922 -804 75978
rect -736 75922 -680 75978
rect -612 75922 -556 75978
rect -488 75922 -432 75978
rect -860 58294 -804 58350
rect -736 58294 -680 58350
rect -612 58294 -556 58350
rect -488 58294 -432 58350
rect -860 58170 -804 58226
rect -736 58170 -680 58226
rect -612 58170 -556 58226
rect -488 58170 -432 58226
rect -860 58046 -804 58102
rect -736 58046 -680 58102
rect -612 58046 -556 58102
rect -488 58046 -432 58102
rect -860 57922 -804 57978
rect -736 57922 -680 57978
rect -612 57922 -556 57978
rect -488 57922 -432 57978
rect -860 40294 -804 40350
rect -736 40294 -680 40350
rect -612 40294 -556 40350
rect -488 40294 -432 40350
rect -860 40170 -804 40226
rect -736 40170 -680 40226
rect -612 40170 -556 40226
rect -488 40170 -432 40226
rect -860 40046 -804 40102
rect -736 40046 -680 40102
rect -612 40046 -556 40102
rect -488 40046 -432 40102
rect -860 39922 -804 39978
rect -736 39922 -680 39978
rect -612 39922 -556 39978
rect -488 39922 -432 39978
rect -860 22294 -804 22350
rect -736 22294 -680 22350
rect -612 22294 -556 22350
rect -488 22294 -432 22350
rect -860 22170 -804 22226
rect -736 22170 -680 22226
rect -612 22170 -556 22226
rect -488 22170 -432 22226
rect -860 22046 -804 22102
rect -736 22046 -680 22102
rect -612 22046 -556 22102
rect -488 22046 -432 22102
rect -860 21922 -804 21978
rect -736 21922 -680 21978
rect -612 21922 -556 21978
rect -488 21922 -432 21978
rect 5514 292294 5570 292350
rect 5638 292294 5694 292350
rect 5762 292294 5818 292350
rect 5886 292294 5942 292350
rect 5514 292170 5570 292226
rect 5638 292170 5694 292226
rect 5762 292170 5818 292226
rect 5886 292170 5942 292226
rect 5514 292046 5570 292102
rect 5638 292046 5694 292102
rect 5762 292046 5818 292102
rect 5886 292046 5942 292102
rect 5514 291922 5570 291978
rect 5638 291922 5694 291978
rect 5762 291922 5818 291978
rect 5886 291922 5942 291978
rect 5514 274294 5570 274350
rect 5638 274294 5694 274350
rect 5762 274294 5818 274350
rect 5886 274294 5942 274350
rect 5514 274170 5570 274226
rect 5638 274170 5694 274226
rect 5762 274170 5818 274226
rect 5886 274170 5942 274226
rect 5514 274046 5570 274102
rect 5638 274046 5694 274102
rect 5762 274046 5818 274102
rect 5886 274046 5942 274102
rect 5514 273922 5570 273978
rect 5638 273922 5694 273978
rect 5762 273922 5818 273978
rect 5886 273922 5942 273978
rect 5514 256294 5570 256350
rect 5638 256294 5694 256350
rect 5762 256294 5818 256350
rect 5886 256294 5942 256350
rect 5514 256170 5570 256226
rect 5638 256170 5694 256226
rect 5762 256170 5818 256226
rect 5886 256170 5942 256226
rect 5514 256046 5570 256102
rect 5638 256046 5694 256102
rect 5762 256046 5818 256102
rect 5886 256046 5942 256102
rect 5514 255922 5570 255978
rect 5638 255922 5694 255978
rect 5762 255922 5818 255978
rect 5886 255922 5942 255978
rect 5514 238294 5570 238350
rect 5638 238294 5694 238350
rect 5762 238294 5818 238350
rect 5886 238294 5942 238350
rect 5514 238170 5570 238226
rect 5638 238170 5694 238226
rect 5762 238170 5818 238226
rect 5886 238170 5942 238226
rect 5514 238046 5570 238102
rect 5638 238046 5694 238102
rect 5762 238046 5818 238102
rect 5886 238046 5942 238102
rect 5514 237922 5570 237978
rect 5638 237922 5694 237978
rect 5762 237922 5818 237978
rect 5886 237922 5942 237978
rect 5514 220294 5570 220350
rect 5638 220294 5694 220350
rect 5762 220294 5818 220350
rect 5886 220294 5942 220350
rect 5514 220170 5570 220226
rect 5638 220170 5694 220226
rect 5762 220170 5818 220226
rect 5886 220170 5942 220226
rect 5514 220046 5570 220102
rect 5638 220046 5694 220102
rect 5762 220046 5818 220102
rect 5886 220046 5942 220102
rect 5514 219922 5570 219978
rect 5638 219922 5694 219978
rect 5762 219922 5818 219978
rect 5886 219922 5942 219978
rect 5514 202294 5570 202350
rect 5638 202294 5694 202350
rect 5762 202294 5818 202350
rect 5886 202294 5942 202350
rect 5514 202170 5570 202226
rect 5638 202170 5694 202226
rect 5762 202170 5818 202226
rect 5886 202170 5942 202226
rect 5514 202046 5570 202102
rect 5638 202046 5694 202102
rect 5762 202046 5818 202102
rect 5886 202046 5942 202102
rect 5514 201922 5570 201978
rect 5638 201922 5694 201978
rect 5762 201922 5818 201978
rect 5886 201922 5942 201978
rect 5514 184294 5570 184350
rect 5638 184294 5694 184350
rect 5762 184294 5818 184350
rect 5886 184294 5942 184350
rect 5514 184170 5570 184226
rect 5638 184170 5694 184226
rect 5762 184170 5818 184226
rect 5886 184170 5942 184226
rect 5514 184046 5570 184102
rect 5638 184046 5694 184102
rect 5762 184046 5818 184102
rect 5886 184046 5942 184102
rect 5514 183922 5570 183978
rect 5638 183922 5694 183978
rect 5762 183922 5818 183978
rect 5886 183922 5942 183978
rect 5514 166294 5570 166350
rect 5638 166294 5694 166350
rect 5762 166294 5818 166350
rect 5886 166294 5942 166350
rect 5514 166170 5570 166226
rect 5638 166170 5694 166226
rect 5762 166170 5818 166226
rect 5886 166170 5942 166226
rect 5514 166046 5570 166102
rect 5638 166046 5694 166102
rect 5762 166046 5818 166102
rect 5886 166046 5942 166102
rect 5514 165922 5570 165978
rect 5638 165922 5694 165978
rect 5762 165922 5818 165978
rect 5886 165922 5942 165978
rect 7532 385442 7588 385498
rect 36234 597156 36290 597212
rect 36358 597156 36414 597212
rect 36482 597156 36538 597212
rect 36606 597156 36662 597212
rect 36234 597032 36290 597088
rect 36358 597032 36414 597088
rect 36482 597032 36538 597088
rect 36606 597032 36662 597088
rect 36234 596908 36290 596964
rect 36358 596908 36414 596964
rect 36482 596908 36538 596964
rect 36606 596908 36662 596964
rect 36234 596784 36290 596840
rect 36358 596784 36414 596840
rect 36482 596784 36538 596840
rect 36606 596784 36662 596840
rect 36234 580294 36290 580350
rect 36358 580294 36414 580350
rect 36482 580294 36538 580350
rect 36606 580294 36662 580350
rect 36234 580170 36290 580226
rect 36358 580170 36414 580226
rect 36482 580170 36538 580226
rect 36606 580170 36662 580226
rect 36234 580046 36290 580102
rect 36358 580046 36414 580102
rect 36482 580046 36538 580102
rect 36606 580046 36662 580102
rect 36234 579922 36290 579978
rect 36358 579922 36414 579978
rect 36482 579922 36538 579978
rect 36606 579922 36662 579978
rect 36234 562294 36290 562350
rect 36358 562294 36414 562350
rect 36482 562294 36538 562350
rect 36606 562294 36662 562350
rect 36234 562170 36290 562226
rect 36358 562170 36414 562226
rect 36482 562170 36538 562226
rect 36606 562170 36662 562226
rect 36234 562046 36290 562102
rect 36358 562046 36414 562102
rect 36482 562046 36538 562102
rect 36606 562046 36662 562102
rect 36234 561922 36290 561978
rect 36358 561922 36414 561978
rect 36482 561922 36538 561978
rect 36606 561922 36662 561978
rect 36234 544294 36290 544350
rect 36358 544294 36414 544350
rect 36482 544294 36538 544350
rect 36606 544294 36662 544350
rect 36234 544170 36290 544226
rect 36358 544170 36414 544226
rect 36482 544170 36538 544226
rect 36606 544170 36662 544226
rect 36234 544046 36290 544102
rect 36358 544046 36414 544102
rect 36482 544046 36538 544102
rect 36606 544046 36662 544102
rect 36234 543922 36290 543978
rect 36358 543922 36414 543978
rect 36482 543922 36538 543978
rect 36606 543922 36662 543978
rect 36234 526294 36290 526350
rect 36358 526294 36414 526350
rect 36482 526294 36538 526350
rect 36606 526294 36662 526350
rect 36234 526170 36290 526226
rect 36358 526170 36414 526226
rect 36482 526170 36538 526226
rect 36606 526170 36662 526226
rect 36234 526046 36290 526102
rect 36358 526046 36414 526102
rect 36482 526046 36538 526102
rect 36606 526046 36662 526102
rect 36234 525922 36290 525978
rect 36358 525922 36414 525978
rect 36482 525922 36538 525978
rect 36606 525922 36662 525978
rect 36234 508294 36290 508350
rect 36358 508294 36414 508350
rect 36482 508294 36538 508350
rect 36606 508294 36662 508350
rect 36234 508170 36290 508226
rect 36358 508170 36414 508226
rect 36482 508170 36538 508226
rect 36606 508170 36662 508226
rect 36234 508046 36290 508102
rect 36358 508046 36414 508102
rect 36482 508046 36538 508102
rect 36606 508046 36662 508102
rect 36234 507922 36290 507978
rect 36358 507922 36414 507978
rect 36482 507922 36538 507978
rect 36606 507922 36662 507978
rect 36234 490294 36290 490350
rect 36358 490294 36414 490350
rect 36482 490294 36538 490350
rect 36606 490294 36662 490350
rect 36234 490170 36290 490226
rect 36358 490170 36414 490226
rect 36482 490170 36538 490226
rect 36606 490170 36662 490226
rect 36234 490046 36290 490102
rect 36358 490046 36414 490102
rect 36482 490046 36538 490102
rect 36606 490046 36662 490102
rect 36234 489922 36290 489978
rect 36358 489922 36414 489978
rect 36482 489922 36538 489978
rect 36606 489922 36662 489978
rect 36234 472294 36290 472350
rect 36358 472294 36414 472350
rect 36482 472294 36538 472350
rect 36606 472294 36662 472350
rect 36234 472170 36290 472226
rect 36358 472170 36414 472226
rect 36482 472170 36538 472226
rect 36606 472170 36662 472226
rect 36234 472046 36290 472102
rect 36358 472046 36414 472102
rect 36482 472046 36538 472102
rect 36606 472046 36662 472102
rect 36234 471922 36290 471978
rect 36358 471922 36414 471978
rect 36482 471922 36538 471978
rect 36606 471922 36662 471978
rect 36234 454294 36290 454350
rect 36358 454294 36414 454350
rect 36482 454294 36538 454350
rect 36606 454294 36662 454350
rect 36234 454170 36290 454226
rect 36358 454170 36414 454226
rect 36482 454170 36538 454226
rect 36606 454170 36662 454226
rect 36234 454046 36290 454102
rect 36358 454046 36414 454102
rect 36482 454046 36538 454102
rect 36606 454046 36662 454102
rect 36234 453922 36290 453978
rect 36358 453922 36414 453978
rect 36482 453922 36538 453978
rect 36606 453922 36662 453978
rect 36234 436294 36290 436350
rect 36358 436294 36414 436350
rect 36482 436294 36538 436350
rect 36606 436294 36662 436350
rect 36234 436170 36290 436226
rect 36358 436170 36414 436226
rect 36482 436170 36538 436226
rect 36606 436170 36662 436226
rect 36234 436046 36290 436102
rect 36358 436046 36414 436102
rect 36482 436046 36538 436102
rect 36606 436046 36662 436102
rect 36234 435922 36290 435978
rect 36358 435922 36414 435978
rect 36482 435922 36538 435978
rect 36606 435922 36662 435978
rect 36234 418294 36290 418350
rect 36358 418294 36414 418350
rect 36482 418294 36538 418350
rect 36606 418294 36662 418350
rect 36234 418170 36290 418226
rect 36358 418170 36414 418226
rect 36482 418170 36538 418226
rect 36606 418170 36662 418226
rect 36234 418046 36290 418102
rect 36358 418046 36414 418102
rect 36482 418046 36538 418102
rect 36606 418046 36662 418102
rect 36234 417922 36290 417978
rect 36358 417922 36414 417978
rect 36482 417922 36538 417978
rect 36606 417922 36662 417978
rect 36234 400294 36290 400350
rect 36358 400294 36414 400350
rect 36482 400294 36538 400350
rect 36606 400294 36662 400350
rect 36234 400170 36290 400226
rect 36358 400170 36414 400226
rect 36482 400170 36538 400226
rect 36606 400170 36662 400226
rect 36234 400046 36290 400102
rect 36358 400046 36414 400102
rect 36482 400046 36538 400102
rect 36606 400046 36662 400102
rect 36234 399922 36290 399978
rect 36358 399922 36414 399978
rect 36482 399922 36538 399978
rect 36606 399922 36662 399978
rect 9234 370294 9290 370350
rect 9358 370294 9414 370350
rect 9482 370294 9538 370350
rect 9606 370294 9662 370350
rect 9234 370170 9290 370226
rect 9358 370170 9414 370226
rect 9482 370170 9538 370226
rect 9606 370170 9662 370226
rect 9234 370046 9290 370102
rect 9358 370046 9414 370102
rect 9482 370046 9538 370102
rect 9606 370046 9662 370102
rect 9234 369922 9290 369978
rect 9358 369922 9414 369978
rect 9482 369922 9538 369978
rect 9606 369922 9662 369978
rect 9234 352294 9290 352350
rect 9358 352294 9414 352350
rect 9482 352294 9538 352350
rect 9606 352294 9662 352350
rect 9234 352170 9290 352226
rect 9358 352170 9414 352226
rect 9482 352170 9538 352226
rect 9606 352170 9662 352226
rect 9234 352046 9290 352102
rect 9358 352046 9414 352102
rect 9482 352046 9538 352102
rect 9606 352046 9662 352102
rect 9234 351922 9290 351978
rect 9358 351922 9414 351978
rect 9482 351922 9538 351978
rect 9606 351922 9662 351978
rect 9234 334294 9290 334350
rect 9358 334294 9414 334350
rect 9482 334294 9538 334350
rect 9606 334294 9662 334350
rect 9234 334170 9290 334226
rect 9358 334170 9414 334226
rect 9482 334170 9538 334226
rect 9606 334170 9662 334226
rect 9234 334046 9290 334102
rect 9358 334046 9414 334102
rect 9482 334046 9538 334102
rect 9606 334046 9662 334102
rect 9234 333922 9290 333978
rect 9358 333922 9414 333978
rect 9482 333922 9538 333978
rect 9606 333922 9662 333978
rect 9234 316294 9290 316350
rect 9358 316294 9414 316350
rect 9482 316294 9538 316350
rect 9606 316294 9662 316350
rect 9234 316170 9290 316226
rect 9358 316170 9414 316226
rect 9482 316170 9538 316226
rect 9606 316170 9662 316226
rect 9234 316046 9290 316102
rect 9358 316046 9414 316102
rect 9482 316046 9538 316102
rect 9606 316046 9662 316102
rect 9234 315922 9290 315978
rect 9358 315922 9414 315978
rect 9482 315922 9538 315978
rect 9606 315922 9662 315978
rect 27692 385262 27748 385318
rect 9234 298294 9290 298350
rect 9358 298294 9414 298350
rect 9482 298294 9538 298350
rect 9606 298294 9662 298350
rect 9234 298170 9290 298226
rect 9358 298170 9414 298226
rect 9482 298170 9538 298226
rect 9606 298170 9662 298226
rect 9234 298046 9290 298102
rect 9358 298046 9414 298102
rect 9482 298046 9538 298102
rect 9606 298046 9662 298102
rect 9234 297922 9290 297978
rect 9358 297922 9414 297978
rect 9482 297922 9538 297978
rect 9606 297922 9662 297978
rect 9234 280294 9290 280350
rect 9358 280294 9414 280350
rect 9482 280294 9538 280350
rect 9606 280294 9662 280350
rect 9234 280170 9290 280226
rect 9358 280170 9414 280226
rect 9482 280170 9538 280226
rect 9606 280170 9662 280226
rect 9234 280046 9290 280102
rect 9358 280046 9414 280102
rect 9482 280046 9538 280102
rect 9606 280046 9662 280102
rect 9234 279922 9290 279978
rect 9358 279922 9414 279978
rect 9482 279922 9538 279978
rect 9606 279922 9662 279978
rect 9234 262294 9290 262350
rect 9358 262294 9414 262350
rect 9482 262294 9538 262350
rect 9606 262294 9662 262350
rect 9234 262170 9290 262226
rect 9358 262170 9414 262226
rect 9482 262170 9538 262226
rect 9606 262170 9662 262226
rect 9234 262046 9290 262102
rect 9358 262046 9414 262102
rect 9482 262046 9538 262102
rect 9606 262046 9662 262102
rect 9234 261922 9290 261978
rect 9358 261922 9414 261978
rect 9482 261922 9538 261978
rect 9606 261922 9662 261978
rect 9234 244294 9290 244350
rect 9358 244294 9414 244350
rect 9482 244294 9538 244350
rect 9606 244294 9662 244350
rect 9234 244170 9290 244226
rect 9358 244170 9414 244226
rect 9482 244170 9538 244226
rect 9606 244170 9662 244226
rect 9234 244046 9290 244102
rect 9358 244046 9414 244102
rect 9482 244046 9538 244102
rect 9606 244046 9662 244102
rect 9234 243922 9290 243978
rect 9358 243922 9414 243978
rect 9482 243922 9538 243978
rect 9606 243922 9662 243978
rect 9234 226294 9290 226350
rect 9358 226294 9414 226350
rect 9482 226294 9538 226350
rect 9606 226294 9662 226350
rect 9234 226170 9290 226226
rect 9358 226170 9414 226226
rect 9482 226170 9538 226226
rect 9606 226170 9662 226226
rect 9234 226046 9290 226102
rect 9358 226046 9414 226102
rect 9482 226046 9538 226102
rect 9606 226046 9662 226102
rect 9234 225922 9290 225978
rect 9358 225922 9414 225978
rect 9482 225922 9538 225978
rect 9606 225922 9662 225978
rect 9234 208294 9290 208350
rect 9358 208294 9414 208350
rect 9482 208294 9538 208350
rect 9606 208294 9662 208350
rect 9234 208170 9290 208226
rect 9358 208170 9414 208226
rect 9482 208170 9538 208226
rect 9606 208170 9662 208226
rect 9234 208046 9290 208102
rect 9358 208046 9414 208102
rect 9482 208046 9538 208102
rect 9606 208046 9662 208102
rect 9234 207922 9290 207978
rect 9358 207922 9414 207978
rect 9482 207922 9538 207978
rect 9606 207922 9662 207978
rect 9234 190294 9290 190350
rect 9358 190294 9414 190350
rect 9482 190294 9538 190350
rect 9606 190294 9662 190350
rect 9234 190170 9290 190226
rect 9358 190170 9414 190226
rect 9482 190170 9538 190226
rect 9606 190170 9662 190226
rect 9234 190046 9290 190102
rect 9358 190046 9414 190102
rect 9482 190046 9538 190102
rect 9606 190046 9662 190102
rect 9234 189922 9290 189978
rect 9358 189922 9414 189978
rect 9482 189922 9538 189978
rect 9606 189922 9662 189978
rect 9234 172294 9290 172350
rect 9358 172294 9414 172350
rect 9482 172294 9538 172350
rect 9606 172294 9662 172350
rect 9234 172170 9290 172226
rect 9358 172170 9414 172226
rect 9482 172170 9538 172226
rect 9606 172170 9662 172226
rect 9234 172046 9290 172102
rect 9358 172046 9414 172102
rect 9482 172046 9538 172102
rect 9606 172046 9662 172102
rect 9234 171922 9290 171978
rect 9358 171922 9414 171978
rect 9482 171922 9538 171978
rect 9606 171922 9662 171978
rect 9234 154294 9290 154350
rect 9358 154294 9414 154350
rect 9482 154294 9538 154350
rect 9606 154294 9662 154350
rect 9234 154170 9290 154226
rect 9358 154170 9414 154226
rect 9482 154170 9538 154226
rect 9606 154170 9662 154226
rect 9234 154046 9290 154102
rect 9358 154046 9414 154102
rect 9482 154046 9538 154102
rect 9606 154046 9662 154102
rect 9234 153922 9290 153978
rect 9358 153922 9414 153978
rect 9482 153922 9538 153978
rect 9606 153922 9662 153978
rect 5514 148294 5570 148350
rect 5638 148294 5694 148350
rect 5762 148294 5818 148350
rect 5886 148294 5942 148350
rect 5514 148170 5570 148226
rect 5638 148170 5694 148226
rect 5762 148170 5818 148226
rect 5886 148170 5942 148226
rect 5514 148046 5570 148102
rect 5638 148046 5694 148102
rect 5762 148046 5818 148102
rect 5886 148046 5942 148102
rect 5514 147922 5570 147978
rect 5638 147922 5694 147978
rect 5762 147922 5818 147978
rect 5886 147922 5942 147978
rect 5514 130294 5570 130350
rect 5638 130294 5694 130350
rect 5762 130294 5818 130350
rect 5886 130294 5942 130350
rect 5514 130170 5570 130226
rect 5638 130170 5694 130226
rect 5762 130170 5818 130226
rect 5886 130170 5942 130226
rect 5514 130046 5570 130102
rect 5638 130046 5694 130102
rect 5762 130046 5818 130102
rect 5886 130046 5942 130102
rect 5514 129922 5570 129978
rect 5638 129922 5694 129978
rect 5762 129922 5818 129978
rect 5886 129922 5942 129978
rect 5514 112294 5570 112350
rect 5638 112294 5694 112350
rect 5762 112294 5818 112350
rect 5886 112294 5942 112350
rect 5514 112170 5570 112226
rect 5638 112170 5694 112226
rect 5762 112170 5818 112226
rect 5886 112170 5942 112226
rect 5514 112046 5570 112102
rect 5638 112046 5694 112102
rect 5762 112046 5818 112102
rect 5886 112046 5942 112102
rect 5514 111922 5570 111978
rect 5638 111922 5694 111978
rect 5762 111922 5818 111978
rect 5886 111922 5942 111978
rect 5514 94294 5570 94350
rect 5638 94294 5694 94350
rect 5762 94294 5818 94350
rect 5886 94294 5942 94350
rect 5514 94170 5570 94226
rect 5638 94170 5694 94226
rect 5762 94170 5818 94226
rect 5886 94170 5942 94226
rect 5514 94046 5570 94102
rect 5638 94046 5694 94102
rect 5762 94046 5818 94102
rect 5886 94046 5942 94102
rect 5514 93922 5570 93978
rect 5638 93922 5694 93978
rect 5762 93922 5818 93978
rect 5886 93922 5942 93978
rect 5514 76294 5570 76350
rect 5638 76294 5694 76350
rect 5762 76294 5818 76350
rect 5886 76294 5942 76350
rect 5514 76170 5570 76226
rect 5638 76170 5694 76226
rect 5762 76170 5818 76226
rect 5886 76170 5942 76226
rect 5514 76046 5570 76102
rect 5638 76046 5694 76102
rect 5762 76046 5818 76102
rect 5886 76046 5942 76102
rect 5514 75922 5570 75978
rect 5638 75922 5694 75978
rect 5762 75922 5818 75978
rect 5886 75922 5942 75978
rect 5514 58294 5570 58350
rect 5638 58294 5694 58350
rect 5762 58294 5818 58350
rect 5886 58294 5942 58350
rect 5514 58170 5570 58226
rect 5638 58170 5694 58226
rect 5762 58170 5818 58226
rect 5886 58170 5942 58226
rect 5514 58046 5570 58102
rect 5638 58046 5694 58102
rect 5762 58046 5818 58102
rect 5886 58046 5942 58102
rect 5514 57922 5570 57978
rect 5638 57922 5694 57978
rect 5762 57922 5818 57978
rect 5886 57922 5942 57978
rect 5514 40294 5570 40350
rect 5638 40294 5694 40350
rect 5762 40294 5818 40350
rect 5886 40294 5942 40350
rect 5514 40170 5570 40226
rect 5638 40170 5694 40226
rect 5762 40170 5818 40226
rect 5886 40170 5942 40226
rect 5514 40046 5570 40102
rect 5638 40046 5694 40102
rect 5762 40046 5818 40102
rect 5886 40046 5942 40102
rect 5514 39922 5570 39978
rect 5638 39922 5694 39978
rect 5762 39922 5818 39978
rect 5886 39922 5942 39978
rect 5514 22294 5570 22350
rect 5638 22294 5694 22350
rect 5762 22294 5818 22350
rect 5886 22294 5942 22350
rect 5514 22170 5570 22226
rect 5638 22170 5694 22226
rect 5762 22170 5818 22226
rect 5886 22170 5942 22226
rect 5514 22046 5570 22102
rect 5638 22046 5694 22102
rect 5762 22046 5818 22102
rect 5886 22046 5942 22102
rect 5514 21922 5570 21978
rect 5638 21922 5694 21978
rect 5762 21922 5818 21978
rect 5886 21922 5942 21978
rect -860 4294 -804 4350
rect -736 4294 -680 4350
rect -612 4294 -556 4350
rect -488 4294 -432 4350
rect -860 4170 -804 4226
rect -736 4170 -680 4226
rect -612 4170 -556 4226
rect -488 4170 -432 4226
rect -860 4046 -804 4102
rect -736 4046 -680 4102
rect -612 4046 -556 4102
rect -488 4046 -432 4102
rect -860 3922 -804 3978
rect -736 3922 -680 3978
rect -612 3922 -556 3978
rect -488 3922 -432 3978
rect -860 -216 -804 -160
rect -736 -216 -680 -160
rect -612 -216 -556 -160
rect -488 -216 -432 -160
rect -860 -340 -804 -284
rect -736 -340 -680 -284
rect -612 -340 -556 -284
rect -488 -340 -432 -284
rect -860 -464 -804 -408
rect -736 -464 -680 -408
rect -612 -464 -556 -408
rect -488 -464 -432 -408
rect -860 -588 -804 -532
rect -736 -588 -680 -532
rect -612 -588 -556 -532
rect -488 -588 -432 -532
rect 5514 4294 5570 4350
rect 5638 4294 5694 4350
rect 5762 4294 5818 4350
rect 5886 4294 5942 4350
rect 5514 4170 5570 4226
rect 5638 4170 5694 4226
rect 5762 4170 5818 4226
rect 5886 4170 5942 4226
rect 5514 4046 5570 4102
rect 5638 4046 5694 4102
rect 5762 4046 5818 4102
rect 5886 4046 5942 4102
rect 5514 3922 5570 3978
rect 5638 3922 5694 3978
rect 5762 3922 5818 3978
rect 5886 3922 5942 3978
rect 5514 -216 5570 -160
rect 5638 -216 5694 -160
rect 5762 -216 5818 -160
rect 5886 -216 5942 -160
rect 5514 -340 5570 -284
rect 5638 -340 5694 -284
rect 5762 -340 5818 -284
rect 5886 -340 5942 -284
rect 5514 -464 5570 -408
rect 5638 -464 5694 -408
rect 5762 -464 5818 -408
rect 5886 -464 5942 -408
rect 5514 -588 5570 -532
rect 5638 -588 5694 -532
rect 5762 -588 5818 -532
rect 5886 -588 5942 -532
rect -1820 -1176 -1764 -1120
rect -1696 -1176 -1640 -1120
rect -1572 -1176 -1516 -1120
rect -1448 -1176 -1392 -1120
rect -1820 -1300 -1764 -1244
rect -1696 -1300 -1640 -1244
rect -1572 -1300 -1516 -1244
rect -1448 -1300 -1392 -1244
rect -1820 -1424 -1764 -1368
rect -1696 -1424 -1640 -1368
rect -1572 -1424 -1516 -1368
rect -1448 -1424 -1392 -1368
rect -1820 -1548 -1764 -1492
rect -1696 -1548 -1640 -1492
rect -1572 -1548 -1516 -1492
rect -1448 -1548 -1392 -1492
rect 9234 136294 9290 136350
rect 9358 136294 9414 136350
rect 9482 136294 9538 136350
rect 9606 136294 9662 136350
rect 9234 136170 9290 136226
rect 9358 136170 9414 136226
rect 9482 136170 9538 136226
rect 9606 136170 9662 136226
rect 9234 136046 9290 136102
rect 9358 136046 9414 136102
rect 9482 136046 9538 136102
rect 9606 136046 9662 136102
rect 9234 135922 9290 135978
rect 9358 135922 9414 135978
rect 9482 135922 9538 135978
rect 9606 135922 9662 135978
rect 9234 118294 9290 118350
rect 9358 118294 9414 118350
rect 9482 118294 9538 118350
rect 9606 118294 9662 118350
rect 9234 118170 9290 118226
rect 9358 118170 9414 118226
rect 9482 118170 9538 118226
rect 9606 118170 9662 118226
rect 9234 118046 9290 118102
rect 9358 118046 9414 118102
rect 9482 118046 9538 118102
rect 9606 118046 9662 118102
rect 9234 117922 9290 117978
rect 9358 117922 9414 117978
rect 9482 117922 9538 117978
rect 9606 117922 9662 117978
rect 9234 100294 9290 100350
rect 9358 100294 9414 100350
rect 9482 100294 9538 100350
rect 9606 100294 9662 100350
rect 9234 100170 9290 100226
rect 9358 100170 9414 100226
rect 9482 100170 9538 100226
rect 9606 100170 9662 100226
rect 9234 100046 9290 100102
rect 9358 100046 9414 100102
rect 9482 100046 9538 100102
rect 9606 100046 9662 100102
rect 9234 99922 9290 99978
rect 9358 99922 9414 99978
rect 9482 99922 9538 99978
rect 9606 99922 9662 99978
rect 9234 82294 9290 82350
rect 9358 82294 9414 82350
rect 9482 82294 9538 82350
rect 9606 82294 9662 82350
rect 9234 82170 9290 82226
rect 9358 82170 9414 82226
rect 9482 82170 9538 82226
rect 9606 82170 9662 82226
rect 9234 82046 9290 82102
rect 9358 82046 9414 82102
rect 9482 82046 9538 82102
rect 9606 82046 9662 82102
rect 9234 81922 9290 81978
rect 9358 81922 9414 81978
rect 9482 81922 9538 81978
rect 9606 81922 9662 81978
rect 36234 382294 36290 382350
rect 36358 382294 36414 382350
rect 36482 382294 36538 382350
rect 36606 382294 36662 382350
rect 36234 382170 36290 382226
rect 36358 382170 36414 382226
rect 36482 382170 36538 382226
rect 36606 382170 36662 382226
rect 36234 382046 36290 382102
rect 36358 382046 36414 382102
rect 36482 382046 36538 382102
rect 36606 382046 36662 382102
rect 36234 381922 36290 381978
rect 36358 381922 36414 381978
rect 36482 381922 36538 381978
rect 36606 381922 36662 381978
rect 36234 364294 36290 364350
rect 36358 364294 36414 364350
rect 36482 364294 36538 364350
rect 36606 364294 36662 364350
rect 36234 364170 36290 364226
rect 36358 364170 36414 364226
rect 36482 364170 36538 364226
rect 36606 364170 36662 364226
rect 36234 364046 36290 364102
rect 36358 364046 36414 364102
rect 36482 364046 36538 364102
rect 36606 364046 36662 364102
rect 36234 363922 36290 363978
rect 36358 363922 36414 363978
rect 36482 363922 36538 363978
rect 36606 363922 36662 363978
rect 36234 346294 36290 346350
rect 36358 346294 36414 346350
rect 36482 346294 36538 346350
rect 36606 346294 36662 346350
rect 36234 346170 36290 346226
rect 36358 346170 36414 346226
rect 36482 346170 36538 346226
rect 36606 346170 36662 346226
rect 36234 346046 36290 346102
rect 36358 346046 36414 346102
rect 36482 346046 36538 346102
rect 36606 346046 36662 346102
rect 36234 345922 36290 345978
rect 36358 345922 36414 345978
rect 36482 345922 36538 345978
rect 36606 345922 36662 345978
rect 36234 328294 36290 328350
rect 36358 328294 36414 328350
rect 36482 328294 36538 328350
rect 36606 328294 36662 328350
rect 36234 328170 36290 328226
rect 36358 328170 36414 328226
rect 36482 328170 36538 328226
rect 36606 328170 36662 328226
rect 36234 328046 36290 328102
rect 36358 328046 36414 328102
rect 36482 328046 36538 328102
rect 36606 328046 36662 328102
rect 36234 327922 36290 327978
rect 36358 327922 36414 327978
rect 36482 327922 36538 327978
rect 36606 327922 36662 327978
rect 36234 310294 36290 310350
rect 36358 310294 36414 310350
rect 36482 310294 36538 310350
rect 36606 310294 36662 310350
rect 36234 310170 36290 310226
rect 36358 310170 36414 310226
rect 36482 310170 36538 310226
rect 36606 310170 36662 310226
rect 36234 310046 36290 310102
rect 36358 310046 36414 310102
rect 36482 310046 36538 310102
rect 36606 310046 36662 310102
rect 36234 309922 36290 309978
rect 36358 309922 36414 309978
rect 36482 309922 36538 309978
rect 36606 309922 36662 309978
rect 36234 292294 36290 292350
rect 36358 292294 36414 292350
rect 36482 292294 36538 292350
rect 36606 292294 36662 292350
rect 36234 292170 36290 292226
rect 36358 292170 36414 292226
rect 36482 292170 36538 292226
rect 36606 292170 36662 292226
rect 36234 292046 36290 292102
rect 36358 292046 36414 292102
rect 36482 292046 36538 292102
rect 36606 292046 36662 292102
rect 36234 291922 36290 291978
rect 36358 291922 36414 291978
rect 36482 291922 36538 291978
rect 36606 291922 36662 291978
rect 36234 274294 36290 274350
rect 36358 274294 36414 274350
rect 36482 274294 36538 274350
rect 36606 274294 36662 274350
rect 36234 274170 36290 274226
rect 36358 274170 36414 274226
rect 36482 274170 36538 274226
rect 36606 274170 36662 274226
rect 36234 274046 36290 274102
rect 36358 274046 36414 274102
rect 36482 274046 36538 274102
rect 36606 274046 36662 274102
rect 36234 273922 36290 273978
rect 36358 273922 36414 273978
rect 36482 273922 36538 273978
rect 36606 273922 36662 273978
rect 36234 256294 36290 256350
rect 36358 256294 36414 256350
rect 36482 256294 36538 256350
rect 36606 256294 36662 256350
rect 36234 256170 36290 256226
rect 36358 256170 36414 256226
rect 36482 256170 36538 256226
rect 36606 256170 36662 256226
rect 36234 256046 36290 256102
rect 36358 256046 36414 256102
rect 36482 256046 36538 256102
rect 36606 256046 36662 256102
rect 36234 255922 36290 255978
rect 36358 255922 36414 255978
rect 36482 255922 36538 255978
rect 36606 255922 36662 255978
rect 36234 238294 36290 238350
rect 36358 238294 36414 238350
rect 36482 238294 36538 238350
rect 36606 238294 36662 238350
rect 36234 238170 36290 238226
rect 36358 238170 36414 238226
rect 36482 238170 36538 238226
rect 36606 238170 36662 238226
rect 36234 238046 36290 238102
rect 36358 238046 36414 238102
rect 36482 238046 36538 238102
rect 36606 238046 36662 238102
rect 36234 237922 36290 237978
rect 36358 237922 36414 237978
rect 36482 237922 36538 237978
rect 36606 237922 36662 237978
rect 36234 220294 36290 220350
rect 36358 220294 36414 220350
rect 36482 220294 36538 220350
rect 36606 220294 36662 220350
rect 36234 220170 36290 220226
rect 36358 220170 36414 220226
rect 36482 220170 36538 220226
rect 36606 220170 36662 220226
rect 36234 220046 36290 220102
rect 36358 220046 36414 220102
rect 36482 220046 36538 220102
rect 36606 220046 36662 220102
rect 36234 219922 36290 219978
rect 36358 219922 36414 219978
rect 36482 219922 36538 219978
rect 36606 219922 36662 219978
rect 36234 202294 36290 202350
rect 36358 202294 36414 202350
rect 36482 202294 36538 202350
rect 36606 202294 36662 202350
rect 36234 202170 36290 202226
rect 36358 202170 36414 202226
rect 36482 202170 36538 202226
rect 36606 202170 36662 202226
rect 36234 202046 36290 202102
rect 36358 202046 36414 202102
rect 36482 202046 36538 202102
rect 36606 202046 36662 202102
rect 36234 201922 36290 201978
rect 36358 201922 36414 201978
rect 36482 201922 36538 201978
rect 36606 201922 36662 201978
rect 36234 184294 36290 184350
rect 36358 184294 36414 184350
rect 36482 184294 36538 184350
rect 36606 184294 36662 184350
rect 36234 184170 36290 184226
rect 36358 184170 36414 184226
rect 36482 184170 36538 184226
rect 36606 184170 36662 184226
rect 36234 184046 36290 184102
rect 36358 184046 36414 184102
rect 36482 184046 36538 184102
rect 36606 184046 36662 184102
rect 36234 183922 36290 183978
rect 36358 183922 36414 183978
rect 36482 183922 36538 183978
rect 36606 183922 36662 183978
rect 36234 166294 36290 166350
rect 36358 166294 36414 166350
rect 36482 166294 36538 166350
rect 36606 166294 36662 166350
rect 36234 166170 36290 166226
rect 36358 166170 36414 166226
rect 36482 166170 36538 166226
rect 36606 166170 36662 166226
rect 36234 166046 36290 166102
rect 36358 166046 36414 166102
rect 36482 166046 36538 166102
rect 36606 166046 36662 166102
rect 36234 165922 36290 165978
rect 36358 165922 36414 165978
rect 36482 165922 36538 165978
rect 36606 165922 36662 165978
rect 36234 148294 36290 148350
rect 36358 148294 36414 148350
rect 36482 148294 36538 148350
rect 36606 148294 36662 148350
rect 36234 148170 36290 148226
rect 36358 148170 36414 148226
rect 36482 148170 36538 148226
rect 36606 148170 36662 148226
rect 36234 148046 36290 148102
rect 36358 148046 36414 148102
rect 36482 148046 36538 148102
rect 36606 148046 36662 148102
rect 36234 147922 36290 147978
rect 36358 147922 36414 147978
rect 36482 147922 36538 147978
rect 36606 147922 36662 147978
rect 36234 130294 36290 130350
rect 36358 130294 36414 130350
rect 36482 130294 36538 130350
rect 36606 130294 36662 130350
rect 36234 130170 36290 130226
rect 36358 130170 36414 130226
rect 36482 130170 36538 130226
rect 36606 130170 36662 130226
rect 36234 130046 36290 130102
rect 36358 130046 36414 130102
rect 36482 130046 36538 130102
rect 36606 130046 36662 130102
rect 36234 129922 36290 129978
rect 36358 129922 36414 129978
rect 36482 129922 36538 129978
rect 36606 129922 36662 129978
rect 36234 112294 36290 112350
rect 36358 112294 36414 112350
rect 36482 112294 36538 112350
rect 36606 112294 36662 112350
rect 36234 112170 36290 112226
rect 36358 112170 36414 112226
rect 36482 112170 36538 112226
rect 36606 112170 36662 112226
rect 36234 112046 36290 112102
rect 36358 112046 36414 112102
rect 36482 112046 36538 112102
rect 36606 112046 36662 112102
rect 36234 111922 36290 111978
rect 36358 111922 36414 111978
rect 36482 111922 36538 111978
rect 36606 111922 36662 111978
rect 36234 94294 36290 94350
rect 36358 94294 36414 94350
rect 36482 94294 36538 94350
rect 36606 94294 36662 94350
rect 36234 94170 36290 94226
rect 36358 94170 36414 94226
rect 36482 94170 36538 94226
rect 36606 94170 36662 94226
rect 36234 94046 36290 94102
rect 36358 94046 36414 94102
rect 36482 94046 36538 94102
rect 36606 94046 36662 94102
rect 36234 93922 36290 93978
rect 36358 93922 36414 93978
rect 36482 93922 36538 93978
rect 36606 93922 36662 93978
rect 36234 76294 36290 76350
rect 36358 76294 36414 76350
rect 36482 76294 36538 76350
rect 36606 76294 36662 76350
rect 36234 76170 36290 76226
rect 36358 76170 36414 76226
rect 36482 76170 36538 76226
rect 36606 76170 36662 76226
rect 36234 76046 36290 76102
rect 36358 76046 36414 76102
rect 36482 76046 36538 76102
rect 36606 76046 36662 76102
rect 36234 75922 36290 75978
rect 36358 75922 36414 75978
rect 36482 75922 36538 75978
rect 36606 75922 36662 75978
rect 9234 64294 9290 64350
rect 9358 64294 9414 64350
rect 9482 64294 9538 64350
rect 9606 64294 9662 64350
rect 9234 64170 9290 64226
rect 9358 64170 9414 64226
rect 9482 64170 9538 64226
rect 9606 64170 9662 64226
rect 9234 64046 9290 64102
rect 9358 64046 9414 64102
rect 9482 64046 9538 64102
rect 9606 64046 9662 64102
rect 9234 63922 9290 63978
rect 9358 63922 9414 63978
rect 9482 63922 9538 63978
rect 9606 63922 9662 63978
rect 9234 46294 9290 46350
rect 9358 46294 9414 46350
rect 9482 46294 9538 46350
rect 9606 46294 9662 46350
rect 9234 46170 9290 46226
rect 9358 46170 9414 46226
rect 9482 46170 9538 46226
rect 9606 46170 9662 46226
rect 9234 46046 9290 46102
rect 9358 46046 9414 46102
rect 9482 46046 9538 46102
rect 9606 46046 9662 46102
rect 9234 45922 9290 45978
rect 9358 45922 9414 45978
rect 9482 45922 9538 45978
rect 9606 45922 9662 45978
rect 9234 28294 9290 28350
rect 9358 28294 9414 28350
rect 9482 28294 9538 28350
rect 9606 28294 9662 28350
rect 9234 28170 9290 28226
rect 9358 28170 9414 28226
rect 9482 28170 9538 28226
rect 9606 28170 9662 28226
rect 9234 28046 9290 28102
rect 9358 28046 9414 28102
rect 9482 28046 9538 28102
rect 9606 28046 9662 28102
rect 9234 27922 9290 27978
rect 9358 27922 9414 27978
rect 9482 27922 9538 27978
rect 9606 27922 9662 27978
rect 9234 10294 9290 10350
rect 9358 10294 9414 10350
rect 9482 10294 9538 10350
rect 9606 10294 9662 10350
rect 9234 10170 9290 10226
rect 9358 10170 9414 10226
rect 9482 10170 9538 10226
rect 9606 10170 9662 10226
rect 9234 10046 9290 10102
rect 9358 10046 9414 10102
rect 9482 10046 9538 10102
rect 9606 10046 9662 10102
rect 9234 9922 9290 9978
rect 9358 9922 9414 9978
rect 9482 9922 9538 9978
rect 9606 9922 9662 9978
rect 9234 -1176 9290 -1120
rect 9358 -1176 9414 -1120
rect 9482 -1176 9538 -1120
rect 9606 -1176 9662 -1120
rect 9234 -1300 9290 -1244
rect 9358 -1300 9414 -1244
rect 9482 -1300 9538 -1244
rect 9606 -1300 9662 -1244
rect 9234 -1424 9290 -1368
rect 9358 -1424 9414 -1368
rect 9482 -1424 9538 -1368
rect 9606 -1424 9662 -1368
rect 9234 -1548 9290 -1492
rect 9358 -1548 9414 -1492
rect 9482 -1548 9538 -1492
rect 9606 -1548 9662 -1492
rect 36234 58294 36290 58350
rect 36358 58294 36414 58350
rect 36482 58294 36538 58350
rect 36606 58294 36662 58350
rect 36234 58170 36290 58226
rect 36358 58170 36414 58226
rect 36482 58170 36538 58226
rect 36606 58170 36662 58226
rect 36234 58046 36290 58102
rect 36358 58046 36414 58102
rect 36482 58046 36538 58102
rect 36606 58046 36662 58102
rect 36234 57922 36290 57978
rect 36358 57922 36414 57978
rect 36482 57922 36538 57978
rect 36606 57922 36662 57978
rect 36234 40294 36290 40350
rect 36358 40294 36414 40350
rect 36482 40294 36538 40350
rect 36606 40294 36662 40350
rect 36234 40170 36290 40226
rect 36358 40170 36414 40226
rect 36482 40170 36538 40226
rect 36606 40170 36662 40226
rect 36234 40046 36290 40102
rect 36358 40046 36414 40102
rect 36482 40046 36538 40102
rect 36606 40046 36662 40102
rect 36234 39922 36290 39978
rect 36358 39922 36414 39978
rect 36482 39922 36538 39978
rect 36606 39922 36662 39978
rect 36234 22294 36290 22350
rect 36358 22294 36414 22350
rect 36482 22294 36538 22350
rect 36606 22294 36662 22350
rect 36234 22170 36290 22226
rect 36358 22170 36414 22226
rect 36482 22170 36538 22226
rect 36606 22170 36662 22226
rect 36234 22046 36290 22102
rect 36358 22046 36414 22102
rect 36482 22046 36538 22102
rect 36606 22046 36662 22102
rect 36234 21922 36290 21978
rect 36358 21922 36414 21978
rect 36482 21922 36538 21978
rect 36606 21922 36662 21978
rect 36234 4294 36290 4350
rect 36358 4294 36414 4350
rect 36482 4294 36538 4350
rect 36606 4294 36662 4350
rect 36234 4170 36290 4226
rect 36358 4170 36414 4226
rect 36482 4170 36538 4226
rect 36606 4170 36662 4226
rect 36234 4046 36290 4102
rect 36358 4046 36414 4102
rect 36482 4046 36538 4102
rect 36606 4046 36662 4102
rect 36234 3922 36290 3978
rect 36358 3922 36414 3978
rect 36482 3922 36538 3978
rect 36606 3922 36662 3978
rect 36234 -216 36290 -160
rect 36358 -216 36414 -160
rect 36482 -216 36538 -160
rect 36606 -216 36662 -160
rect 36234 -340 36290 -284
rect 36358 -340 36414 -284
rect 36482 -340 36538 -284
rect 36606 -340 36662 -284
rect 36234 -464 36290 -408
rect 36358 -464 36414 -408
rect 36482 -464 36538 -408
rect 36606 -464 36662 -408
rect 36234 -588 36290 -532
rect 36358 -588 36414 -532
rect 36482 -588 36538 -532
rect 36606 -588 36662 -532
rect 39954 598116 40010 598172
rect 40078 598116 40134 598172
rect 40202 598116 40258 598172
rect 40326 598116 40382 598172
rect 39954 597992 40010 598048
rect 40078 597992 40134 598048
rect 40202 597992 40258 598048
rect 40326 597992 40382 598048
rect 39954 597868 40010 597924
rect 40078 597868 40134 597924
rect 40202 597868 40258 597924
rect 40326 597868 40382 597924
rect 39954 597744 40010 597800
rect 40078 597744 40134 597800
rect 40202 597744 40258 597800
rect 40326 597744 40382 597800
rect 39954 586294 40010 586350
rect 40078 586294 40134 586350
rect 40202 586294 40258 586350
rect 40326 586294 40382 586350
rect 39954 586170 40010 586226
rect 40078 586170 40134 586226
rect 40202 586170 40258 586226
rect 40326 586170 40382 586226
rect 39954 586046 40010 586102
rect 40078 586046 40134 586102
rect 40202 586046 40258 586102
rect 40326 586046 40382 586102
rect 39954 585922 40010 585978
rect 40078 585922 40134 585978
rect 40202 585922 40258 585978
rect 40326 585922 40382 585978
rect 39954 568294 40010 568350
rect 40078 568294 40134 568350
rect 40202 568294 40258 568350
rect 40326 568294 40382 568350
rect 39954 568170 40010 568226
rect 40078 568170 40134 568226
rect 40202 568170 40258 568226
rect 40326 568170 40382 568226
rect 39954 568046 40010 568102
rect 40078 568046 40134 568102
rect 40202 568046 40258 568102
rect 40326 568046 40382 568102
rect 39954 567922 40010 567978
rect 40078 567922 40134 567978
rect 40202 567922 40258 567978
rect 40326 567922 40382 567978
rect 39954 550294 40010 550350
rect 40078 550294 40134 550350
rect 40202 550294 40258 550350
rect 40326 550294 40382 550350
rect 39954 550170 40010 550226
rect 40078 550170 40134 550226
rect 40202 550170 40258 550226
rect 40326 550170 40382 550226
rect 39954 550046 40010 550102
rect 40078 550046 40134 550102
rect 40202 550046 40258 550102
rect 40326 550046 40382 550102
rect 39954 549922 40010 549978
rect 40078 549922 40134 549978
rect 40202 549922 40258 549978
rect 40326 549922 40382 549978
rect 66954 597156 67010 597212
rect 67078 597156 67134 597212
rect 67202 597156 67258 597212
rect 67326 597156 67382 597212
rect 66954 597032 67010 597088
rect 67078 597032 67134 597088
rect 67202 597032 67258 597088
rect 67326 597032 67382 597088
rect 66954 596908 67010 596964
rect 67078 596908 67134 596964
rect 67202 596908 67258 596964
rect 67326 596908 67382 596964
rect 66954 596784 67010 596840
rect 67078 596784 67134 596840
rect 67202 596784 67258 596840
rect 67326 596784 67382 596840
rect 66954 580294 67010 580350
rect 67078 580294 67134 580350
rect 67202 580294 67258 580350
rect 67326 580294 67382 580350
rect 66954 580170 67010 580226
rect 67078 580170 67134 580226
rect 67202 580170 67258 580226
rect 67326 580170 67382 580226
rect 66954 580046 67010 580102
rect 67078 580046 67134 580102
rect 67202 580046 67258 580102
rect 67326 580046 67382 580102
rect 66954 579922 67010 579978
rect 67078 579922 67134 579978
rect 67202 579922 67258 579978
rect 67326 579922 67382 579978
rect 66954 562294 67010 562350
rect 67078 562294 67134 562350
rect 67202 562294 67258 562350
rect 67326 562294 67382 562350
rect 66954 562170 67010 562226
rect 67078 562170 67134 562226
rect 67202 562170 67258 562226
rect 67326 562170 67382 562226
rect 66954 562046 67010 562102
rect 67078 562046 67134 562102
rect 67202 562046 67258 562102
rect 67326 562046 67382 562102
rect 66954 561922 67010 561978
rect 67078 561922 67134 561978
rect 67202 561922 67258 561978
rect 67326 561922 67382 561978
rect 66954 544294 67010 544350
rect 67078 544294 67134 544350
rect 67202 544294 67258 544350
rect 67326 544294 67382 544350
rect 66954 544170 67010 544226
rect 67078 544170 67134 544226
rect 67202 544170 67258 544226
rect 67326 544170 67382 544226
rect 66954 544046 67010 544102
rect 67078 544046 67134 544102
rect 67202 544046 67258 544102
rect 67326 544046 67382 544102
rect 66954 543922 67010 543978
rect 67078 543922 67134 543978
rect 67202 543922 67258 543978
rect 67326 543922 67382 543978
rect 70674 598116 70730 598172
rect 70798 598116 70854 598172
rect 70922 598116 70978 598172
rect 71046 598116 71102 598172
rect 70674 597992 70730 598048
rect 70798 597992 70854 598048
rect 70922 597992 70978 598048
rect 71046 597992 71102 598048
rect 70674 597868 70730 597924
rect 70798 597868 70854 597924
rect 70922 597868 70978 597924
rect 71046 597868 71102 597924
rect 70674 597744 70730 597800
rect 70798 597744 70854 597800
rect 70922 597744 70978 597800
rect 71046 597744 71102 597800
rect 70674 586294 70730 586350
rect 70798 586294 70854 586350
rect 70922 586294 70978 586350
rect 71046 586294 71102 586350
rect 70674 586170 70730 586226
rect 70798 586170 70854 586226
rect 70922 586170 70978 586226
rect 71046 586170 71102 586226
rect 70674 586046 70730 586102
rect 70798 586046 70854 586102
rect 70922 586046 70978 586102
rect 71046 586046 71102 586102
rect 70674 585922 70730 585978
rect 70798 585922 70854 585978
rect 70922 585922 70978 585978
rect 71046 585922 71102 585978
rect 70674 568294 70730 568350
rect 70798 568294 70854 568350
rect 70922 568294 70978 568350
rect 71046 568294 71102 568350
rect 70674 568170 70730 568226
rect 70798 568170 70854 568226
rect 70922 568170 70978 568226
rect 71046 568170 71102 568226
rect 70674 568046 70730 568102
rect 70798 568046 70854 568102
rect 70922 568046 70978 568102
rect 71046 568046 71102 568102
rect 70674 567922 70730 567978
rect 70798 567922 70854 567978
rect 70922 567922 70978 567978
rect 71046 567922 71102 567978
rect 70674 550294 70730 550350
rect 70798 550294 70854 550350
rect 70922 550294 70978 550350
rect 71046 550294 71102 550350
rect 70674 550170 70730 550226
rect 70798 550170 70854 550226
rect 70922 550170 70978 550226
rect 71046 550170 71102 550226
rect 70674 550046 70730 550102
rect 70798 550046 70854 550102
rect 70922 550046 70978 550102
rect 71046 550046 71102 550102
rect 70674 549922 70730 549978
rect 70798 549922 70854 549978
rect 70922 549922 70978 549978
rect 71046 549922 71102 549978
rect 97674 597156 97730 597212
rect 97798 597156 97854 597212
rect 97922 597156 97978 597212
rect 98046 597156 98102 597212
rect 97674 597032 97730 597088
rect 97798 597032 97854 597088
rect 97922 597032 97978 597088
rect 98046 597032 98102 597088
rect 97674 596908 97730 596964
rect 97798 596908 97854 596964
rect 97922 596908 97978 596964
rect 98046 596908 98102 596964
rect 97674 596784 97730 596840
rect 97798 596784 97854 596840
rect 97922 596784 97978 596840
rect 98046 596784 98102 596840
rect 97674 580294 97730 580350
rect 97798 580294 97854 580350
rect 97922 580294 97978 580350
rect 98046 580294 98102 580350
rect 97674 580170 97730 580226
rect 97798 580170 97854 580226
rect 97922 580170 97978 580226
rect 98046 580170 98102 580226
rect 97674 580046 97730 580102
rect 97798 580046 97854 580102
rect 97922 580046 97978 580102
rect 98046 580046 98102 580102
rect 97674 579922 97730 579978
rect 97798 579922 97854 579978
rect 97922 579922 97978 579978
rect 98046 579922 98102 579978
rect 97674 562294 97730 562350
rect 97798 562294 97854 562350
rect 97922 562294 97978 562350
rect 98046 562294 98102 562350
rect 97674 562170 97730 562226
rect 97798 562170 97854 562226
rect 97922 562170 97978 562226
rect 98046 562170 98102 562226
rect 97674 562046 97730 562102
rect 97798 562046 97854 562102
rect 97922 562046 97978 562102
rect 98046 562046 98102 562102
rect 97674 561922 97730 561978
rect 97798 561922 97854 561978
rect 97922 561922 97978 561978
rect 98046 561922 98102 561978
rect 101394 598116 101450 598172
rect 101518 598116 101574 598172
rect 101642 598116 101698 598172
rect 101766 598116 101822 598172
rect 101394 597992 101450 598048
rect 101518 597992 101574 598048
rect 101642 597992 101698 598048
rect 101766 597992 101822 598048
rect 101394 597868 101450 597924
rect 101518 597868 101574 597924
rect 101642 597868 101698 597924
rect 101766 597868 101822 597924
rect 101394 597744 101450 597800
rect 101518 597744 101574 597800
rect 101642 597744 101698 597800
rect 101766 597744 101822 597800
rect 101394 586294 101450 586350
rect 101518 586294 101574 586350
rect 101642 586294 101698 586350
rect 101766 586294 101822 586350
rect 101394 586170 101450 586226
rect 101518 586170 101574 586226
rect 101642 586170 101698 586226
rect 101766 586170 101822 586226
rect 101394 586046 101450 586102
rect 101518 586046 101574 586102
rect 101642 586046 101698 586102
rect 101766 586046 101822 586102
rect 101394 585922 101450 585978
rect 101518 585922 101574 585978
rect 101642 585922 101698 585978
rect 101766 585922 101822 585978
rect 101394 568294 101450 568350
rect 101518 568294 101574 568350
rect 101642 568294 101698 568350
rect 101766 568294 101822 568350
rect 101394 568170 101450 568226
rect 101518 568170 101574 568226
rect 101642 568170 101698 568226
rect 101766 568170 101822 568226
rect 101394 568046 101450 568102
rect 101518 568046 101574 568102
rect 101642 568046 101698 568102
rect 101766 568046 101822 568102
rect 101394 567922 101450 567978
rect 101518 567922 101574 567978
rect 101642 567922 101698 567978
rect 101766 567922 101822 567978
rect 128394 597156 128450 597212
rect 128518 597156 128574 597212
rect 128642 597156 128698 597212
rect 128766 597156 128822 597212
rect 128394 597032 128450 597088
rect 128518 597032 128574 597088
rect 128642 597032 128698 597088
rect 128766 597032 128822 597088
rect 128394 596908 128450 596964
rect 128518 596908 128574 596964
rect 128642 596908 128698 596964
rect 128766 596908 128822 596964
rect 128394 596784 128450 596840
rect 128518 596784 128574 596840
rect 128642 596784 128698 596840
rect 128766 596784 128822 596840
rect 128394 580294 128450 580350
rect 128518 580294 128574 580350
rect 128642 580294 128698 580350
rect 128766 580294 128822 580350
rect 128394 580170 128450 580226
rect 128518 580170 128574 580226
rect 128642 580170 128698 580226
rect 128766 580170 128822 580226
rect 128394 580046 128450 580102
rect 128518 580046 128574 580102
rect 128642 580046 128698 580102
rect 128766 580046 128822 580102
rect 128394 579922 128450 579978
rect 128518 579922 128574 579978
rect 128642 579922 128698 579978
rect 128766 579922 128822 579978
rect 128394 562294 128450 562350
rect 128518 562294 128574 562350
rect 128642 562294 128698 562350
rect 128766 562294 128822 562350
rect 128394 562170 128450 562226
rect 128518 562170 128574 562226
rect 128642 562170 128698 562226
rect 128766 562170 128822 562226
rect 114035 561947 114091 562003
rect 114159 561947 114215 562003
rect 114283 561947 114339 562003
rect 114407 561947 114463 562003
rect 114531 561947 114587 562003
rect 114655 561947 114711 562003
rect 114779 561947 114835 562003
rect 114903 561947 114959 562003
rect 115027 561947 115083 562003
rect 115151 561947 115207 562003
rect 115275 561947 115331 562003
rect 115399 561947 115455 562003
rect 115523 561947 115579 562003
rect 115647 561947 115703 562003
rect 115771 561947 115827 562003
rect 115895 561947 115951 562003
rect 116019 561947 116075 562003
rect 116143 561947 116199 562003
rect 116267 561947 116323 562003
rect 116391 561947 116447 562003
rect 116515 561947 116571 562003
rect 116639 561947 116695 562003
rect 116763 561947 116819 562003
rect 116887 561947 116943 562003
rect 117011 561947 117067 562003
rect 117135 561947 117191 562003
rect 117259 561947 117315 562003
rect 117383 561947 117439 562003
rect 117507 561947 117563 562003
rect 117631 561947 117687 562003
rect 117755 561947 117811 562003
rect 117879 561947 117935 562003
rect 118003 561947 118059 562003
rect 118127 561947 118183 562003
rect 118251 561947 118307 562003
rect 118375 561947 118431 562003
rect 118499 561947 118555 562003
rect 118623 561947 118679 562003
rect 118747 561947 118803 562003
rect 118871 561947 118927 562003
rect 118995 561947 119051 562003
rect 119119 561947 119175 562003
rect 119243 561947 119299 562003
rect 119367 561947 119423 562003
rect 119491 561947 119547 562003
rect 119615 561947 119671 562003
rect 119739 561947 119795 562003
rect 119863 561947 119919 562003
rect 119987 561947 120043 562003
rect 120111 561947 120167 562003
rect 120235 561947 120291 562003
rect 120359 561947 120415 562003
rect 128394 562046 128450 562102
rect 128518 562046 128574 562102
rect 128642 562046 128698 562102
rect 128766 562046 128822 562102
rect 128394 561922 128450 561978
rect 128518 561922 128574 561978
rect 128642 561922 128698 561978
rect 128766 561922 128822 561978
rect 101394 550294 101450 550350
rect 101518 550294 101574 550350
rect 101642 550294 101698 550350
rect 101766 550294 101822 550350
rect 101394 550170 101450 550226
rect 101518 550170 101574 550226
rect 101642 550170 101698 550226
rect 101766 550170 101822 550226
rect 101394 550046 101450 550102
rect 101518 550046 101574 550102
rect 101642 550046 101698 550102
rect 101766 550046 101822 550102
rect 101394 549922 101450 549978
rect 101518 549922 101574 549978
rect 101642 549922 101698 549978
rect 101766 549922 101822 549978
rect 132114 598116 132170 598172
rect 132238 598116 132294 598172
rect 132362 598116 132418 598172
rect 132486 598116 132542 598172
rect 132114 597992 132170 598048
rect 132238 597992 132294 598048
rect 132362 597992 132418 598048
rect 132486 597992 132542 598048
rect 132114 597868 132170 597924
rect 132238 597868 132294 597924
rect 132362 597868 132418 597924
rect 132486 597868 132542 597924
rect 132114 597744 132170 597800
rect 132238 597744 132294 597800
rect 132362 597744 132418 597800
rect 132486 597744 132542 597800
rect 132114 586294 132170 586350
rect 132238 586294 132294 586350
rect 132362 586294 132418 586350
rect 132486 586294 132542 586350
rect 132114 586170 132170 586226
rect 132238 586170 132294 586226
rect 132362 586170 132418 586226
rect 132486 586170 132542 586226
rect 132114 586046 132170 586102
rect 132238 586046 132294 586102
rect 132362 586046 132418 586102
rect 132486 586046 132542 586102
rect 132114 585922 132170 585978
rect 132238 585922 132294 585978
rect 132362 585922 132418 585978
rect 132486 585922 132542 585978
rect 132114 568294 132170 568350
rect 132238 568294 132294 568350
rect 132362 568294 132418 568350
rect 132486 568294 132542 568350
rect 132114 568170 132170 568226
rect 132238 568170 132294 568226
rect 132362 568170 132418 568226
rect 132486 568170 132542 568226
rect 132114 568046 132170 568102
rect 132238 568046 132294 568102
rect 132362 568046 132418 568102
rect 132486 568046 132542 568102
rect 132114 567922 132170 567978
rect 132238 567922 132294 567978
rect 132362 567922 132418 567978
rect 132486 567922 132542 567978
rect 132114 550294 132170 550350
rect 132238 550294 132294 550350
rect 132362 550294 132418 550350
rect 132486 550294 132542 550350
rect 132114 550170 132170 550226
rect 132238 550170 132294 550226
rect 132362 550170 132418 550226
rect 132486 550170 132542 550226
rect 132114 550046 132170 550102
rect 132238 550046 132294 550102
rect 132362 550046 132418 550102
rect 132486 550046 132542 550102
rect 132114 549922 132170 549978
rect 132238 549922 132294 549978
rect 132362 549922 132418 549978
rect 132486 549922 132542 549978
rect 159114 597156 159170 597212
rect 159238 597156 159294 597212
rect 159362 597156 159418 597212
rect 159486 597156 159542 597212
rect 159114 597032 159170 597088
rect 159238 597032 159294 597088
rect 159362 597032 159418 597088
rect 159486 597032 159542 597088
rect 159114 596908 159170 596964
rect 159238 596908 159294 596964
rect 159362 596908 159418 596964
rect 159486 596908 159542 596964
rect 159114 596784 159170 596840
rect 159238 596784 159294 596840
rect 159362 596784 159418 596840
rect 159486 596784 159542 596840
rect 159114 580294 159170 580350
rect 159238 580294 159294 580350
rect 159362 580294 159418 580350
rect 159486 580294 159542 580350
rect 159114 580170 159170 580226
rect 159238 580170 159294 580226
rect 159362 580170 159418 580226
rect 159486 580170 159542 580226
rect 159114 580046 159170 580102
rect 159238 580046 159294 580102
rect 159362 580046 159418 580102
rect 159486 580046 159542 580102
rect 159114 579922 159170 579978
rect 159238 579922 159294 579978
rect 159362 579922 159418 579978
rect 159486 579922 159542 579978
rect 159114 562294 159170 562350
rect 159238 562294 159294 562350
rect 159362 562294 159418 562350
rect 159486 562294 159542 562350
rect 159114 562170 159170 562226
rect 159238 562170 159294 562226
rect 159362 562170 159418 562226
rect 159486 562170 159542 562226
rect 159114 562046 159170 562102
rect 159238 562046 159294 562102
rect 159362 562046 159418 562102
rect 159486 562046 159542 562102
rect 159114 561922 159170 561978
rect 159238 561922 159294 561978
rect 159362 561922 159418 561978
rect 159486 561922 159542 561978
rect 97674 544294 97730 544350
rect 97798 544294 97854 544350
rect 97922 544294 97978 544350
rect 98046 544294 98102 544350
rect 97674 544170 97730 544226
rect 97798 544170 97854 544226
rect 97922 544170 97978 544226
rect 98046 544170 98102 544226
rect 97674 544046 97730 544102
rect 97798 544046 97854 544102
rect 97922 544046 97978 544102
rect 98046 544046 98102 544102
rect 100965 544234 101021 544290
rect 100965 544110 101021 544166
rect 101089 544234 101145 544290
rect 101213 544234 101269 544290
rect 101337 544234 101393 544290
rect 101461 544234 101517 544290
rect 101089 544110 101145 544166
rect 101213 544110 101269 544166
rect 101337 544110 101393 544166
rect 101461 544110 101517 544166
rect 101585 544234 101641 544290
rect 101709 544234 101765 544290
rect 101833 544234 101889 544290
rect 101957 544234 102013 544290
rect 101585 544110 101641 544166
rect 101709 544110 101765 544166
rect 101833 544110 101889 544166
rect 101957 544110 102013 544166
rect 102081 544234 102137 544290
rect 102205 544234 102261 544290
rect 102329 544234 102385 544290
rect 102453 544234 102509 544290
rect 102081 544110 102137 544166
rect 102205 544110 102261 544166
rect 102329 544110 102385 544166
rect 102453 544110 102509 544166
rect 102577 544234 102633 544290
rect 102701 544234 102757 544290
rect 102825 544234 102881 544290
rect 102949 544234 103005 544290
rect 102577 544110 102633 544166
rect 102701 544110 102757 544166
rect 102825 544110 102881 544166
rect 102949 544110 103005 544166
rect 103073 544234 103129 544290
rect 103197 544234 103253 544290
rect 103321 544234 103377 544290
rect 103445 544234 103501 544290
rect 103073 544110 103129 544166
rect 103197 544110 103253 544166
rect 103321 544110 103377 544166
rect 103445 544110 103501 544166
rect 103569 544234 103625 544290
rect 103693 544234 103749 544290
rect 103817 544234 103873 544290
rect 103941 544234 103997 544290
rect 103569 544110 103625 544166
rect 103693 544110 103749 544166
rect 103817 544110 103873 544166
rect 103941 544110 103997 544166
rect 104065 544234 104121 544290
rect 104189 544234 104245 544290
rect 104313 544234 104369 544290
rect 104437 544234 104493 544290
rect 104065 544110 104121 544166
rect 104189 544110 104245 544166
rect 104313 544110 104369 544166
rect 104437 544110 104493 544166
rect 104561 544234 104617 544290
rect 104685 544234 104741 544290
rect 104809 544234 104865 544290
rect 104933 544234 104989 544290
rect 104561 544110 104617 544166
rect 104685 544110 104741 544166
rect 104809 544110 104865 544166
rect 104933 544110 104989 544166
rect 105057 544234 105113 544290
rect 105181 544234 105237 544290
rect 105305 544234 105361 544290
rect 105429 544234 105485 544290
rect 105057 544110 105113 544166
rect 105181 544110 105237 544166
rect 105305 544110 105361 544166
rect 105429 544110 105485 544166
rect 105553 544234 105609 544290
rect 105677 544234 105733 544290
rect 105801 544234 105857 544290
rect 105925 544234 105981 544290
rect 105553 544110 105609 544166
rect 105677 544110 105733 544166
rect 105801 544110 105857 544166
rect 105925 544110 105981 544166
rect 106049 544234 106105 544290
rect 106173 544234 106229 544290
rect 106297 544234 106353 544290
rect 106421 544234 106477 544290
rect 106049 544110 106105 544166
rect 106173 544110 106229 544166
rect 106297 544110 106353 544166
rect 106421 544110 106477 544166
rect 106545 544234 106601 544290
rect 106669 544234 106725 544290
rect 106793 544234 106849 544290
rect 106917 544234 106973 544290
rect 106545 544110 106601 544166
rect 106669 544110 106725 544166
rect 106793 544110 106849 544166
rect 106917 544110 106973 544166
rect 107041 544234 107097 544290
rect 107165 544234 107221 544290
rect 107289 544234 107345 544290
rect 107413 544234 107469 544290
rect 107041 544110 107097 544166
rect 107165 544110 107221 544166
rect 107289 544110 107345 544166
rect 107413 544110 107469 544166
rect 107537 544234 107593 544290
rect 107661 544234 107717 544290
rect 107785 544234 107841 544290
rect 107909 544234 107965 544290
rect 107537 544110 107593 544166
rect 107661 544110 107717 544166
rect 107785 544110 107841 544166
rect 107909 544110 107965 544166
rect 108033 544234 108089 544290
rect 108157 544234 108213 544290
rect 108281 544234 108337 544290
rect 108405 544234 108461 544290
rect 108033 544110 108089 544166
rect 108157 544110 108213 544166
rect 108281 544110 108337 544166
rect 108405 544110 108461 544166
rect 108529 544234 108585 544290
rect 108653 544234 108709 544290
rect 108777 544234 108833 544290
rect 108901 544234 108957 544290
rect 108529 544110 108585 544166
rect 108653 544110 108709 544166
rect 108777 544110 108833 544166
rect 108901 544110 108957 544166
rect 109025 544234 109081 544290
rect 109149 544234 109205 544290
rect 109273 544234 109329 544290
rect 109397 544234 109453 544290
rect 109025 544110 109081 544166
rect 109149 544110 109205 544166
rect 109273 544110 109329 544166
rect 109397 544110 109453 544166
rect 109521 544234 109577 544290
rect 109645 544234 109701 544290
rect 109769 544234 109825 544290
rect 109893 544234 109949 544290
rect 109521 544110 109577 544166
rect 109645 544110 109701 544166
rect 109769 544110 109825 544166
rect 109893 544110 109949 544166
rect 110017 544234 110073 544290
rect 110141 544234 110197 544290
rect 110265 544234 110321 544290
rect 110389 544234 110445 544290
rect 110017 544110 110073 544166
rect 110141 544110 110197 544166
rect 110265 544110 110321 544166
rect 110389 544110 110445 544166
rect 110513 544234 110569 544290
rect 110637 544234 110693 544290
rect 110761 544234 110817 544290
rect 110885 544234 110941 544290
rect 110513 544110 110569 544166
rect 110637 544110 110693 544166
rect 110761 544110 110817 544166
rect 110885 544110 110941 544166
rect 111009 544234 111065 544290
rect 111133 544234 111189 544290
rect 111257 544234 111313 544290
rect 111381 544234 111437 544290
rect 111009 544110 111065 544166
rect 111133 544110 111189 544166
rect 111257 544110 111313 544166
rect 111381 544110 111437 544166
rect 111505 544234 111561 544290
rect 111629 544234 111685 544290
rect 111753 544234 111809 544290
rect 111877 544234 111933 544290
rect 111505 544110 111561 544166
rect 111629 544110 111685 544166
rect 111753 544110 111809 544166
rect 111877 544110 111933 544166
rect 112001 544234 112057 544290
rect 112125 544234 112181 544290
rect 112249 544234 112305 544290
rect 112373 544234 112429 544290
rect 112001 544110 112057 544166
rect 112125 544110 112181 544166
rect 112249 544110 112305 544166
rect 112373 544110 112429 544166
rect 112497 544234 112553 544290
rect 112621 544234 112677 544290
rect 112745 544234 112801 544290
rect 112869 544234 112925 544290
rect 112497 544110 112553 544166
rect 112621 544110 112677 544166
rect 112745 544110 112801 544166
rect 112869 544110 112925 544166
rect 112993 544234 113049 544290
rect 113117 544234 113173 544290
rect 113241 544234 113297 544290
rect 113365 544234 113421 544290
rect 112993 544110 113049 544166
rect 113117 544110 113173 544166
rect 113241 544110 113297 544166
rect 113365 544110 113421 544166
rect 113489 544234 113545 544290
rect 113613 544234 113669 544290
rect 113737 544234 113793 544290
rect 113861 544234 113917 544290
rect 113489 544110 113545 544166
rect 113613 544110 113669 544166
rect 113737 544110 113793 544166
rect 113861 544110 113917 544166
rect 113985 544234 114041 544290
rect 114109 544234 114165 544290
rect 114233 544234 114289 544290
rect 114357 544234 114413 544290
rect 113985 544110 114041 544166
rect 114109 544110 114165 544166
rect 114233 544110 114289 544166
rect 114357 544110 114413 544166
rect 114481 544234 114537 544290
rect 114605 544234 114661 544290
rect 114729 544234 114785 544290
rect 114853 544234 114909 544290
rect 114481 544110 114537 544166
rect 114605 544110 114661 544166
rect 114729 544110 114785 544166
rect 114853 544110 114909 544166
rect 114977 544234 115033 544290
rect 115101 544234 115157 544290
rect 115225 544234 115281 544290
rect 115349 544234 115405 544290
rect 114977 544110 115033 544166
rect 115101 544110 115157 544166
rect 115225 544110 115281 544166
rect 115349 544110 115405 544166
rect 115473 544234 115529 544290
rect 115597 544234 115653 544290
rect 115721 544234 115777 544290
rect 115845 544234 115901 544290
rect 115473 544110 115529 544166
rect 115597 544110 115653 544166
rect 115721 544110 115777 544166
rect 115845 544110 115901 544166
rect 115969 544234 116025 544290
rect 116093 544234 116149 544290
rect 116217 544234 116273 544290
rect 116341 544234 116397 544290
rect 115969 544110 116025 544166
rect 116093 544110 116149 544166
rect 116217 544110 116273 544166
rect 116341 544110 116397 544166
rect 116465 544234 116521 544290
rect 116589 544234 116645 544290
rect 116713 544234 116769 544290
rect 116837 544234 116893 544290
rect 116465 544110 116521 544166
rect 116589 544110 116645 544166
rect 116713 544110 116769 544166
rect 116837 544110 116893 544166
rect 116961 544234 117017 544290
rect 117085 544234 117141 544290
rect 117209 544234 117265 544290
rect 117333 544234 117389 544290
rect 116961 544110 117017 544166
rect 117085 544110 117141 544166
rect 117209 544110 117265 544166
rect 117333 544110 117389 544166
rect 117457 544234 117513 544290
rect 117581 544234 117637 544290
rect 117705 544234 117761 544290
rect 117829 544234 117885 544290
rect 117457 544110 117513 544166
rect 117581 544110 117637 544166
rect 117705 544110 117761 544166
rect 117829 544110 117885 544166
rect 128394 544294 128450 544350
rect 128518 544294 128574 544350
rect 128642 544294 128698 544350
rect 128766 544294 128822 544350
rect 128394 544170 128450 544226
rect 128518 544170 128574 544226
rect 128642 544170 128698 544226
rect 128766 544170 128822 544226
rect 97674 543922 97730 543978
rect 97798 543922 97854 543978
rect 97922 543922 97978 543978
rect 98046 543922 98102 543978
rect 128394 544046 128450 544102
rect 128518 544046 128574 544102
rect 128642 544046 128698 544102
rect 128766 544046 128822 544102
rect 128394 543922 128450 543978
rect 128518 543922 128574 543978
rect 128642 543922 128698 543978
rect 128766 543922 128822 543978
rect 100823 543835 100879 543891
rect 100927 543835 100983 543891
rect 101031 543835 101087 543891
rect 101135 543835 101191 543891
rect 101239 543835 101295 543891
rect 101343 543835 101399 543891
rect 101447 543835 101503 543891
rect 101551 543835 101607 543891
rect 101655 543835 101711 543891
rect 101759 543835 101815 543891
rect 101863 543835 101919 543891
rect 101967 543835 102023 543891
rect 102071 543835 102127 543891
rect 102175 543835 102231 543891
rect 102279 543835 102335 543891
rect 102383 543835 102439 543891
rect 102487 543835 102543 543891
rect 102591 543835 102647 543891
rect 102695 543835 102751 543891
rect 102799 543835 102855 543891
rect 102903 543835 102959 543891
rect 103007 543835 103063 543891
rect 103111 543835 103167 543891
rect 103215 543835 103271 543891
rect 103319 543835 103375 543891
rect 103423 543835 103479 543891
rect 103527 543835 103583 543891
rect 103631 543835 103687 543891
rect 103735 543835 103791 543891
rect 103839 543835 103895 543891
rect 103943 543835 103999 543891
rect 104047 543835 104103 543891
rect 104151 543835 104207 543891
rect 104255 543835 104311 543891
rect 104359 543835 104415 543891
rect 104463 543835 104519 543891
rect 104567 543835 104623 543891
rect 104671 543835 104727 543891
rect 104775 543835 104831 543891
rect 104879 543835 104935 543891
rect 104983 543835 105039 543891
rect 105087 543835 105143 543891
rect 105191 543835 105247 543891
rect 105295 543835 105351 543891
rect 105399 543835 105455 543891
rect 105503 543835 105559 543891
rect 105607 543835 105663 543891
rect 105711 543835 105767 543891
rect 105815 543835 105871 543891
rect 105919 543835 105975 543891
rect 106023 543835 106079 543891
rect 106127 543835 106183 543891
rect 106231 543835 106287 543891
rect 106335 543835 106391 543891
rect 106439 543835 106495 543891
rect 106543 543835 106599 543891
rect 106647 543835 106703 543891
rect 106751 543835 106807 543891
rect 106855 543835 106911 543891
rect 106959 543835 107015 543891
rect 107063 543835 107119 543891
rect 107167 543835 107223 543891
rect 107271 543835 107327 543891
rect 107375 543835 107431 543891
rect 107479 543835 107535 543891
rect 107583 543835 107639 543891
rect 107687 543835 107743 543891
rect 107791 543835 107847 543891
rect 107895 543835 107951 543891
rect 107999 543835 108055 543891
rect 108103 543835 108159 543891
rect 108207 543835 108263 543891
rect 108311 543835 108367 543891
rect 108415 543835 108471 543891
rect 108519 543835 108575 543891
rect 108623 543835 108679 543891
rect 108727 543835 108783 543891
rect 108831 543835 108887 543891
rect 108935 543835 108991 543891
rect 109039 543835 109095 543891
rect 109143 543835 109199 543891
rect 109247 543835 109303 543891
rect 109351 543835 109407 543891
rect 109455 543835 109511 543891
rect 109559 543835 109615 543891
rect 109663 543835 109719 543891
rect 109767 543835 109823 543891
rect 109871 543835 109927 543891
rect 109975 543835 110031 543891
rect 110079 543835 110135 543891
rect 110183 543835 110239 543891
rect 110287 543835 110343 543891
rect 110391 543835 110447 543891
rect 110495 543835 110551 543891
rect 110599 543835 110655 543891
rect 110703 543835 110759 543891
rect 110807 543835 110863 543891
rect 110911 543835 110967 543891
rect 111015 543835 111071 543891
rect 111119 543835 111175 543891
rect 111223 543835 111279 543891
rect 111327 543835 111383 543891
rect 111431 543835 111487 543891
rect 111535 543835 111591 543891
rect 111639 543835 111695 543891
rect 111743 543835 111799 543891
rect 111847 543835 111903 543891
rect 111951 543835 112007 543891
rect 112055 543835 112111 543891
rect 112159 543835 112215 543891
rect 112263 543835 112319 543891
rect 112367 543835 112423 543891
rect 112471 543835 112527 543891
rect 112575 543835 112631 543891
rect 112679 543835 112735 543891
rect 112783 543835 112839 543891
rect 112887 543835 112943 543891
rect 112991 543835 113047 543891
rect 113095 543835 113151 543891
rect 113199 543835 113255 543891
rect 113303 543835 113359 543891
rect 113407 543835 113463 543891
rect 113511 543835 113567 543891
rect 113615 543835 113671 543891
rect 113719 543835 113775 543891
rect 113823 543835 113879 543891
rect 113927 543835 113983 543891
rect 114031 543835 114087 543891
rect 114135 543835 114191 543891
rect 114239 543835 114295 543891
rect 114343 543835 114399 543891
rect 114447 543835 114503 543891
rect 114551 543835 114607 543891
rect 114655 543835 114711 543891
rect 114759 543835 114815 543891
rect 114863 543835 114919 543891
rect 114967 543835 115023 543891
rect 115071 543835 115127 543891
rect 115175 543835 115231 543891
rect 115279 543835 115335 543891
rect 115383 543835 115439 543891
rect 115487 543835 115543 543891
rect 115591 543835 115647 543891
rect 115695 543835 115751 543891
rect 115799 543835 115855 543891
rect 115903 543835 115959 543891
rect 116007 543835 116063 543891
rect 116111 543835 116167 543891
rect 116215 543835 116271 543891
rect 116319 543835 116375 543891
rect 116423 543835 116479 543891
rect 116527 543835 116583 543891
rect 116631 543835 116687 543891
rect 116735 543835 116791 543891
rect 116839 543835 116895 543891
rect 116943 543835 116999 543891
rect 117047 543835 117103 543891
rect 117151 543835 117207 543891
rect 117255 543835 117311 543891
rect 117359 543835 117415 543891
rect 117463 543835 117519 543891
rect 117567 543835 117623 543891
rect 117671 543835 117727 543891
rect 159114 544294 159170 544350
rect 159238 544294 159294 544350
rect 159362 544294 159418 544350
rect 159486 544294 159542 544350
rect 159114 544170 159170 544226
rect 159238 544170 159294 544226
rect 159362 544170 159418 544226
rect 159486 544170 159542 544226
rect 159114 544046 159170 544102
rect 159238 544046 159294 544102
rect 159362 544046 159418 544102
rect 159486 544046 159542 544102
rect 159114 543922 159170 543978
rect 159238 543922 159294 543978
rect 159362 543922 159418 543978
rect 159486 543922 159542 543978
rect 39954 532294 40010 532350
rect 40078 532294 40134 532350
rect 40202 532294 40258 532350
rect 40326 532294 40382 532350
rect 39954 532170 40010 532226
rect 40078 532170 40134 532226
rect 40202 532170 40258 532226
rect 40326 532170 40382 532226
rect 69507 532247 69563 532303
rect 69631 532247 69687 532303
rect 69755 532247 69811 532303
rect 69879 532247 69935 532303
rect 70003 532247 70059 532303
rect 70127 532247 70183 532303
rect 70251 532247 70307 532303
rect 70375 532247 70431 532303
rect 70499 532247 70555 532303
rect 70623 532247 70679 532303
rect 70747 532247 70803 532303
rect 70871 532247 70927 532303
rect 70995 532247 71051 532303
rect 71119 532247 71175 532303
rect 71243 532247 71299 532303
rect 71367 532247 71423 532303
rect 71491 532247 71547 532303
rect 71615 532247 71671 532303
rect 71739 532247 71795 532303
rect 71863 532247 71919 532303
rect 71987 532247 72043 532303
rect 72111 532247 72167 532303
rect 72235 532247 72291 532303
rect 72359 532247 72415 532303
rect 72483 532247 72539 532303
rect 72607 532247 72663 532303
rect 72731 532247 72787 532303
rect 72855 532247 72911 532303
rect 72979 532247 73035 532303
rect 73103 532247 73159 532303
rect 73227 532247 73283 532303
rect 73351 532247 73407 532303
rect 73475 532247 73531 532303
rect 73599 532247 73655 532303
rect 73723 532247 73779 532303
rect 73847 532247 73903 532303
rect 73971 532247 74027 532303
rect 74095 532247 74151 532303
rect 74219 532247 74275 532303
rect 74343 532247 74399 532303
rect 74467 532247 74523 532303
rect 74591 532247 74647 532303
rect 74715 532247 74771 532303
rect 74839 532247 74895 532303
rect 74963 532247 75019 532303
rect 75087 532247 75143 532303
rect 75211 532247 75267 532303
rect 75335 532247 75391 532303
rect 75459 532247 75515 532303
rect 75583 532247 75639 532303
rect 75707 532247 75763 532303
rect 75831 532247 75887 532303
rect 75955 532247 76011 532303
rect 76079 532247 76135 532303
rect 76203 532247 76259 532303
rect 76327 532247 76383 532303
rect 76451 532247 76507 532303
rect 76575 532247 76631 532303
rect 76699 532247 76755 532303
rect 76823 532247 76879 532303
rect 76947 532247 77003 532303
rect 77071 532247 77127 532303
rect 77195 532247 77251 532303
rect 77319 532247 77375 532303
rect 77443 532247 77499 532303
rect 77567 532247 77623 532303
rect 77691 532247 77747 532303
rect 77815 532247 77871 532303
rect 77939 532247 77995 532303
rect 78063 532247 78119 532303
rect 78187 532247 78243 532303
rect 39954 532046 40010 532102
rect 40078 532046 40134 532102
rect 40202 532046 40258 532102
rect 40326 532046 40382 532102
rect 39954 531922 40010 531978
rect 40078 531922 40134 531978
rect 40202 531922 40258 531978
rect 40326 531922 40382 531978
rect 69181 531947 69237 532003
rect 69305 531947 69361 532003
rect 69429 531947 69485 532003
rect 69553 531947 69609 532003
rect 69677 531947 69733 532003
rect 69801 531947 69857 532003
rect 69925 531947 69981 532003
rect 70049 531947 70105 532003
rect 70173 531947 70229 532003
rect 70297 531947 70353 532003
rect 70421 531947 70477 532003
rect 70545 531947 70601 532003
rect 70669 531947 70725 532003
rect 70793 531947 70849 532003
rect 70917 531947 70973 532003
rect 71041 531947 71097 532003
rect 71165 531947 71221 532003
rect 71289 531947 71345 532003
rect 71413 531947 71469 532003
rect 71537 531947 71593 532003
rect 71661 531947 71717 532003
rect 71785 531947 71841 532003
rect 71909 531947 71965 532003
rect 72033 531947 72089 532003
rect 72157 531947 72213 532003
rect 72281 531947 72337 532003
rect 72405 531947 72461 532003
rect 72529 531947 72585 532003
rect 72653 531947 72709 532003
rect 72777 531947 72833 532003
rect 72901 531947 72957 532003
rect 73025 531947 73081 532003
rect 73149 531947 73205 532003
rect 73273 531947 73329 532003
rect 73397 531947 73453 532003
rect 73521 531947 73577 532003
rect 73645 531947 73701 532003
rect 73769 531947 73825 532003
rect 73893 531947 73949 532003
rect 74017 531947 74073 532003
rect 74141 531947 74197 532003
rect 74265 531947 74321 532003
rect 74389 531947 74445 532003
rect 74513 531947 74569 532003
rect 74637 531947 74693 532003
rect 74761 531947 74817 532003
rect 74885 531947 74941 532003
rect 75009 531947 75065 532003
rect 75133 531947 75189 532003
rect 75257 531947 75313 532003
rect 75381 531947 75437 532003
rect 75505 531947 75561 532003
rect 75629 531947 75685 532003
rect 75753 531947 75809 532003
rect 75877 531947 75933 532003
rect 76001 531947 76057 532003
rect 76125 531947 76181 532003
rect 76249 531947 76305 532003
rect 76373 531947 76429 532003
rect 76497 531947 76553 532003
rect 76621 531947 76677 532003
rect 76745 531947 76801 532003
rect 76869 531947 76925 532003
rect 76993 531947 77049 532003
rect 77117 531947 77173 532003
rect 77241 531947 77297 532003
rect 77365 531947 77421 532003
rect 77489 531947 77545 532003
rect 77613 531947 77669 532003
rect 159114 526294 159170 526350
rect 159238 526294 159294 526350
rect 159362 526294 159418 526350
rect 159486 526294 159542 526350
rect 91381 526097 91437 526153
rect 91505 526097 91561 526153
rect 91629 526097 91685 526153
rect 91753 526097 91809 526153
rect 91877 526097 91933 526153
rect 92001 526097 92057 526153
rect 92125 526097 92181 526153
rect 92249 526097 92305 526153
rect 92373 526097 92429 526153
rect 92497 526097 92553 526153
rect 92621 526097 92677 526153
rect 92745 526097 92801 526153
rect 92869 526097 92925 526153
rect 92993 526097 93049 526153
rect 93117 526097 93173 526153
rect 93241 526097 93297 526153
rect 93365 526097 93421 526153
rect 93489 526097 93545 526153
rect 93613 526097 93669 526153
rect 93737 526097 93793 526153
rect 93861 526097 93917 526153
rect 93985 526097 94041 526153
rect 94109 526097 94165 526153
rect 94233 526097 94289 526153
rect 94357 526097 94413 526153
rect 94481 526097 94537 526153
rect 94605 526097 94661 526153
rect 94729 526097 94785 526153
rect 94853 526097 94909 526153
rect 94977 526097 95033 526153
rect 95101 526097 95157 526153
rect 95225 526097 95281 526153
rect 95349 526097 95405 526153
rect 95473 526097 95529 526153
rect 95597 526097 95653 526153
rect 95721 526097 95777 526153
rect 95845 526097 95901 526153
rect 95969 526097 96025 526153
rect 96093 526097 96149 526153
rect 96217 526097 96273 526153
rect 96341 526097 96397 526153
rect 96465 526097 96521 526153
rect 96589 526097 96645 526153
rect 96713 526097 96769 526153
rect 96837 526097 96893 526153
rect 96961 526097 97017 526153
rect 97085 526097 97141 526153
rect 97209 526097 97265 526153
rect 97333 526097 97389 526153
rect 97457 526097 97513 526153
rect 97581 526097 97637 526153
rect 97705 526097 97761 526153
rect 97829 526097 97885 526153
rect 97953 526097 98009 526153
rect 98077 526097 98133 526153
rect 98201 526097 98257 526153
rect 98325 526097 98381 526153
rect 98449 526097 98505 526153
rect 98573 526097 98629 526153
rect 98697 526097 98753 526153
rect 98821 526097 98877 526153
rect 98945 526097 99001 526153
rect 99069 526097 99125 526153
rect 99193 526097 99249 526153
rect 99317 526097 99373 526153
rect 99441 526097 99497 526153
rect 99565 526097 99621 526153
rect 99689 526097 99745 526153
rect 99813 526097 99869 526153
rect 99937 526097 99993 526153
rect 100061 526097 100117 526153
rect 100185 526097 100241 526153
rect 100309 526097 100365 526153
rect 100433 526097 100489 526153
rect 100557 526097 100613 526153
rect 100681 526097 100737 526153
rect 100805 526097 100861 526153
rect 100929 526097 100985 526153
rect 101053 526097 101109 526153
rect 101177 526097 101233 526153
rect 101301 526097 101357 526153
rect 101425 526097 101481 526153
rect 101549 526097 101605 526153
rect 101673 526097 101729 526153
rect 101797 526097 101853 526153
rect 101921 526097 101977 526153
rect 102045 526097 102101 526153
rect 102169 526097 102225 526153
rect 102293 526097 102349 526153
rect 102417 526097 102473 526153
rect 102541 526097 102597 526153
rect 102665 526097 102721 526153
rect 102789 526097 102845 526153
rect 102913 526097 102969 526153
rect 103037 526097 103093 526153
rect 103161 526097 103217 526153
rect 103285 526097 103341 526153
rect 103409 526097 103465 526153
rect 103533 526097 103589 526153
rect 103657 526097 103713 526153
rect 103781 526097 103837 526153
rect 103905 526097 103961 526153
rect 104029 526097 104085 526153
rect 104153 526097 104209 526153
rect 104277 526097 104333 526153
rect 104401 526097 104457 526153
rect 104525 526097 104581 526153
rect 104649 526097 104705 526153
rect 104773 526097 104829 526153
rect 104897 526097 104953 526153
rect 105021 526097 105077 526153
rect 105145 526097 105201 526153
rect 105269 526097 105325 526153
rect 105393 526097 105449 526153
rect 105517 526097 105573 526153
rect 105641 526097 105697 526153
rect 105765 526097 105821 526153
rect 105889 526097 105945 526153
rect 106013 526097 106069 526153
rect 106137 526097 106193 526153
rect 106261 526097 106317 526153
rect 106385 526097 106441 526153
rect 106509 526097 106565 526153
rect 106633 526097 106689 526153
rect 106757 526097 106813 526153
rect 106881 526097 106937 526153
rect 107005 526097 107061 526153
rect 107129 526097 107185 526153
rect 107253 526097 107309 526153
rect 107377 526097 107433 526153
rect 107501 526097 107557 526153
rect 107625 526097 107681 526153
rect 107749 526097 107805 526153
rect 107873 526097 107929 526153
rect 107997 526097 108053 526153
rect 108121 526097 108177 526153
rect 108245 526097 108301 526153
rect 108369 526097 108425 526153
rect 108493 526097 108549 526153
rect 108617 526097 108673 526153
rect 108741 526097 108797 526153
rect 108865 526097 108921 526153
rect 108989 526097 109045 526153
rect 109113 526097 109169 526153
rect 159114 526170 159170 526226
rect 159238 526170 159294 526226
rect 159362 526170 159418 526226
rect 159486 526170 159542 526226
rect 159114 526046 159170 526102
rect 159238 526046 159294 526102
rect 159362 526046 159418 526102
rect 159486 526046 159542 526102
rect 159114 525922 159170 525978
rect 159238 525922 159294 525978
rect 159362 525922 159418 525978
rect 159486 525922 159542 525978
rect 91234 525835 91290 525891
rect 91338 525835 91394 525891
rect 91442 525835 91498 525891
rect 91546 525835 91602 525891
rect 91650 525835 91706 525891
rect 91754 525835 91810 525891
rect 91858 525835 91914 525891
rect 91962 525835 92018 525891
rect 92066 525835 92122 525891
rect 92170 525835 92226 525891
rect 92274 525835 92330 525891
rect 92378 525835 92434 525891
rect 92482 525835 92538 525891
rect 92586 525835 92642 525891
rect 92690 525835 92746 525891
rect 92794 525835 92850 525891
rect 92898 525835 92954 525891
rect 93002 525835 93058 525891
rect 93106 525835 93162 525891
rect 93210 525835 93266 525891
rect 93314 525835 93370 525891
rect 93418 525835 93474 525891
rect 93522 525835 93578 525891
rect 93626 525835 93682 525891
rect 93730 525835 93786 525891
rect 93834 525835 93890 525891
rect 93938 525835 93994 525891
rect 94042 525835 94098 525891
rect 94146 525835 94202 525891
rect 94250 525835 94306 525891
rect 94354 525835 94410 525891
rect 94458 525835 94514 525891
rect 94562 525835 94618 525891
rect 94666 525835 94722 525891
rect 94770 525835 94826 525891
rect 94874 525835 94930 525891
rect 94978 525835 95034 525891
rect 95082 525835 95138 525891
rect 95186 525835 95242 525891
rect 95290 525835 95346 525891
rect 95394 525835 95450 525891
rect 95498 525835 95554 525891
rect 95602 525835 95658 525891
rect 95706 525835 95762 525891
rect 95810 525835 95866 525891
rect 95914 525835 95970 525891
rect 96018 525835 96074 525891
rect 96122 525835 96178 525891
rect 96226 525835 96282 525891
rect 96330 525835 96386 525891
rect 96434 525835 96490 525891
rect 96538 525835 96594 525891
rect 96642 525835 96698 525891
rect 96746 525835 96802 525891
rect 96850 525835 96906 525891
rect 96954 525835 97010 525891
rect 97058 525835 97114 525891
rect 97162 525835 97218 525891
rect 97266 525835 97322 525891
rect 97370 525835 97426 525891
rect 97474 525835 97530 525891
rect 97578 525835 97634 525891
rect 97682 525835 97738 525891
rect 97786 525835 97842 525891
rect 97890 525835 97946 525891
rect 97994 525835 98050 525891
rect 98098 525835 98154 525891
rect 98202 525835 98258 525891
rect 98306 525835 98362 525891
rect 98410 525835 98466 525891
rect 98514 525835 98570 525891
rect 98618 525835 98674 525891
rect 98722 525835 98778 525891
rect 98826 525835 98882 525891
rect 98930 525835 98986 525891
rect 99034 525835 99090 525891
rect 99138 525835 99194 525891
rect 99242 525835 99298 525891
rect 99346 525835 99402 525891
rect 99450 525835 99506 525891
rect 99554 525835 99610 525891
rect 99658 525835 99714 525891
rect 99762 525835 99818 525891
rect 99866 525835 99922 525891
rect 99970 525835 100026 525891
rect 100074 525835 100130 525891
rect 100178 525835 100234 525891
rect 100282 525835 100338 525891
rect 100386 525835 100442 525891
rect 100490 525835 100546 525891
rect 100594 525835 100650 525891
rect 100698 525835 100754 525891
rect 100802 525835 100858 525891
rect 100906 525835 100962 525891
rect 101010 525835 101066 525891
rect 101114 525835 101170 525891
rect 101218 525835 101274 525891
rect 101322 525835 101378 525891
rect 101426 525835 101482 525891
rect 101530 525835 101586 525891
rect 101634 525835 101690 525891
rect 101738 525835 101794 525891
rect 101842 525835 101898 525891
rect 101946 525835 102002 525891
rect 102050 525835 102106 525891
rect 102154 525835 102210 525891
rect 102258 525835 102314 525891
rect 102362 525835 102418 525891
rect 102466 525835 102522 525891
rect 102570 525835 102626 525891
rect 102674 525835 102730 525891
rect 102778 525835 102834 525891
rect 102882 525835 102938 525891
rect 102986 525835 103042 525891
rect 103090 525835 103146 525891
rect 103194 525835 103250 525891
rect 103298 525835 103354 525891
rect 103402 525835 103458 525891
rect 103506 525835 103562 525891
rect 103610 525835 103666 525891
rect 103714 525835 103770 525891
rect 103818 525835 103874 525891
rect 103922 525835 103978 525891
rect 104026 525835 104082 525891
rect 104130 525835 104186 525891
rect 104234 525835 104290 525891
rect 104338 525835 104394 525891
rect 104442 525835 104498 525891
rect 104546 525835 104602 525891
rect 104650 525835 104706 525891
rect 104754 525835 104810 525891
rect 104858 525835 104914 525891
rect 104962 525835 105018 525891
rect 105066 525835 105122 525891
rect 105170 525835 105226 525891
rect 105274 525835 105330 525891
rect 105378 525835 105434 525891
rect 105482 525835 105538 525891
rect 105586 525835 105642 525891
rect 105690 525835 105746 525891
rect 105794 525835 105850 525891
rect 105898 525835 105954 525891
rect 106002 525835 106058 525891
rect 106106 525835 106162 525891
rect 106210 525835 106266 525891
rect 106314 525835 106370 525891
rect 106418 525835 106474 525891
rect 106522 525835 106578 525891
rect 106626 525835 106682 525891
rect 106730 525835 106786 525891
rect 106834 525835 106890 525891
rect 106938 525835 106994 525891
rect 107042 525835 107098 525891
rect 107146 525835 107202 525891
rect 107250 525835 107306 525891
rect 107354 525835 107410 525891
rect 107458 525835 107514 525891
rect 107562 525835 107618 525891
rect 107666 525835 107722 525891
rect 107770 525835 107826 525891
rect 107874 525835 107930 525891
rect 107978 525835 108034 525891
rect 108082 525835 108138 525891
rect 108186 525835 108242 525891
rect 108290 525835 108346 525891
rect 108394 525835 108450 525891
rect 108498 525835 108554 525891
rect 108602 525835 108658 525891
rect 108706 525835 108762 525891
rect 108810 525835 108866 525891
rect 39954 514294 40010 514350
rect 40078 514294 40134 514350
rect 40202 514294 40258 514350
rect 40326 514294 40382 514350
rect 39954 514170 40010 514226
rect 40078 514170 40134 514226
rect 40202 514170 40258 514226
rect 40326 514170 40382 514226
rect 39954 514046 40010 514102
rect 40078 514046 40134 514102
rect 40202 514046 40258 514102
rect 40326 514046 40382 514102
rect 39954 513922 40010 513978
rect 40078 513922 40134 513978
rect 40202 513922 40258 513978
rect 40326 513922 40382 513978
rect 60355 514356 60411 514412
rect 60479 514356 60535 514412
rect 60603 514356 60659 514412
rect 60727 514356 60783 514412
rect 60851 514356 60907 514412
rect 60975 514356 61031 514412
rect 61099 514356 61155 514412
rect 61223 514356 61279 514412
rect 61347 514356 61403 514412
rect 61471 514356 61527 514412
rect 61595 514356 61651 514412
rect 61719 514356 61775 514412
rect 61843 514356 61899 514412
rect 61967 514356 62023 514412
rect 62091 514356 62147 514412
rect 62215 514356 62271 514412
rect 62339 514356 62395 514412
rect 62463 514356 62519 514412
rect 62587 514356 62643 514412
rect 62711 514356 62767 514412
rect 62835 514356 62891 514412
rect 62959 514356 63015 514412
rect 63083 514356 63139 514412
rect 63207 514356 63263 514412
rect 63331 514356 63387 514412
rect 63455 514356 63511 514412
rect 63579 514356 63635 514412
rect 63703 514356 63759 514412
rect 63827 514356 63883 514412
rect 63951 514356 64007 514412
rect 64075 514356 64131 514412
rect 64199 514356 64255 514412
rect 64323 514356 64379 514412
rect 64447 514356 64503 514412
rect 64571 514356 64627 514412
rect 64695 514356 64751 514412
rect 64819 514356 64875 514412
rect 64943 514356 64999 514412
rect 65067 514356 65123 514412
rect 65191 514356 65247 514412
rect 65315 514356 65371 514412
rect 65439 514356 65495 514412
rect 60355 514232 60411 514288
rect 60479 514232 60535 514288
rect 60603 514232 60659 514288
rect 60727 514232 60783 514288
rect 60851 514232 60907 514288
rect 60975 514232 61031 514288
rect 61099 514232 61155 514288
rect 61223 514232 61279 514288
rect 61347 514232 61403 514288
rect 61471 514232 61527 514288
rect 61595 514232 61651 514288
rect 61719 514232 61775 514288
rect 61843 514232 61899 514288
rect 61967 514232 62023 514288
rect 62091 514232 62147 514288
rect 62215 514232 62271 514288
rect 62339 514232 62395 514288
rect 62463 514232 62519 514288
rect 62587 514232 62643 514288
rect 62711 514232 62767 514288
rect 62835 514232 62891 514288
rect 62959 514232 63015 514288
rect 63083 514232 63139 514288
rect 63207 514232 63263 514288
rect 63331 514232 63387 514288
rect 63455 514232 63511 514288
rect 63579 514232 63635 514288
rect 63703 514232 63759 514288
rect 63827 514232 63883 514288
rect 63951 514232 64007 514288
rect 64075 514232 64131 514288
rect 64199 514232 64255 514288
rect 64323 514232 64379 514288
rect 64447 514232 64503 514288
rect 64571 514232 64627 514288
rect 64695 514232 64751 514288
rect 64819 514232 64875 514288
rect 64943 514232 64999 514288
rect 65067 514232 65123 514288
rect 65191 514232 65247 514288
rect 65315 514232 65371 514288
rect 65439 514232 65495 514288
rect 60355 514108 60411 514164
rect 60479 514108 60535 514164
rect 60603 514108 60659 514164
rect 60727 514108 60783 514164
rect 60851 514108 60907 514164
rect 60975 514108 61031 514164
rect 61099 514108 61155 514164
rect 61223 514108 61279 514164
rect 61347 514108 61403 514164
rect 61471 514108 61527 514164
rect 61595 514108 61651 514164
rect 61719 514108 61775 514164
rect 61843 514108 61899 514164
rect 61967 514108 62023 514164
rect 62091 514108 62147 514164
rect 62215 514108 62271 514164
rect 62339 514108 62395 514164
rect 62463 514108 62519 514164
rect 62587 514108 62643 514164
rect 62711 514108 62767 514164
rect 62835 514108 62891 514164
rect 62959 514108 63015 514164
rect 63083 514108 63139 514164
rect 63207 514108 63263 514164
rect 63331 514108 63387 514164
rect 63455 514108 63511 514164
rect 63579 514108 63635 514164
rect 63703 514108 63759 514164
rect 63827 514108 63883 514164
rect 63951 514108 64007 514164
rect 64075 514108 64131 514164
rect 64199 514108 64255 514164
rect 64323 514108 64379 514164
rect 64447 514108 64503 514164
rect 64571 514108 64627 514164
rect 64695 514108 64751 514164
rect 64819 514108 64875 514164
rect 64943 514108 64999 514164
rect 65067 514108 65123 514164
rect 65191 514108 65247 514164
rect 65315 514108 65371 514164
rect 65439 514108 65495 514164
rect 60355 513984 60411 514040
rect 60479 513984 60535 514040
rect 60603 513984 60659 514040
rect 60727 513984 60783 514040
rect 60851 513984 60907 514040
rect 60975 513984 61031 514040
rect 61099 513984 61155 514040
rect 61223 513984 61279 514040
rect 61347 513984 61403 514040
rect 61471 513984 61527 514040
rect 61595 513984 61651 514040
rect 61719 513984 61775 514040
rect 61843 513984 61899 514040
rect 61967 513984 62023 514040
rect 62091 513984 62147 514040
rect 62215 513984 62271 514040
rect 62339 513984 62395 514040
rect 62463 513984 62519 514040
rect 62587 513984 62643 514040
rect 62711 513984 62767 514040
rect 62835 513984 62891 514040
rect 62959 513984 63015 514040
rect 63083 513984 63139 514040
rect 63207 513984 63263 514040
rect 63331 513984 63387 514040
rect 63455 513984 63511 514040
rect 63579 513984 63635 514040
rect 63703 513984 63759 514040
rect 63827 513984 63883 514040
rect 63951 513984 64007 514040
rect 64075 513984 64131 514040
rect 64199 513984 64255 514040
rect 64323 513984 64379 514040
rect 64447 513984 64503 514040
rect 64571 513984 64627 514040
rect 64695 513984 64751 514040
rect 64819 513984 64875 514040
rect 64943 513984 64999 514040
rect 65067 513984 65123 514040
rect 65191 513984 65247 514040
rect 65315 513984 65371 514040
rect 65439 513984 65495 514040
rect 60355 513860 60411 513916
rect 60479 513860 60535 513916
rect 60603 513860 60659 513916
rect 60727 513860 60783 513916
rect 60851 513860 60907 513916
rect 60975 513860 61031 513916
rect 61099 513860 61155 513916
rect 61223 513860 61279 513916
rect 61347 513860 61403 513916
rect 61471 513860 61527 513916
rect 61595 513860 61651 513916
rect 61719 513860 61775 513916
rect 61843 513860 61899 513916
rect 61967 513860 62023 513916
rect 62091 513860 62147 513916
rect 62215 513860 62271 513916
rect 62339 513860 62395 513916
rect 62463 513860 62519 513916
rect 62587 513860 62643 513916
rect 62711 513860 62767 513916
rect 62835 513860 62891 513916
rect 62959 513860 63015 513916
rect 63083 513860 63139 513916
rect 63207 513860 63263 513916
rect 63331 513860 63387 513916
rect 63455 513860 63511 513916
rect 63579 513860 63635 513916
rect 63703 513860 63759 513916
rect 63827 513860 63883 513916
rect 63951 513860 64007 513916
rect 64075 513860 64131 513916
rect 64199 513860 64255 513916
rect 64323 513860 64379 513916
rect 64447 513860 64503 513916
rect 64571 513860 64627 513916
rect 64695 513860 64751 513916
rect 64819 513860 64875 513916
rect 64943 513860 64999 513916
rect 65067 513860 65123 513916
rect 65191 513860 65247 513916
rect 65315 513860 65371 513916
rect 65439 513860 65495 513916
rect 85231 508234 85287 508290
rect 85231 508110 85287 508166
rect 85355 508234 85411 508290
rect 85479 508234 85535 508290
rect 85603 508234 85659 508290
rect 85727 508234 85783 508290
rect 85355 508110 85411 508166
rect 85479 508110 85535 508166
rect 85603 508110 85659 508166
rect 85727 508110 85783 508166
rect 85851 508234 85907 508290
rect 85975 508234 86031 508290
rect 86099 508234 86155 508290
rect 86223 508234 86279 508290
rect 85851 508110 85907 508166
rect 85975 508110 86031 508166
rect 86099 508110 86155 508166
rect 86223 508110 86279 508166
rect 86347 508234 86403 508290
rect 86471 508234 86527 508290
rect 86595 508234 86651 508290
rect 86719 508234 86775 508290
rect 86347 508110 86403 508166
rect 86471 508110 86527 508166
rect 86595 508110 86651 508166
rect 86719 508110 86775 508166
rect 86843 508234 86899 508290
rect 86967 508234 87023 508290
rect 87091 508234 87147 508290
rect 87215 508234 87271 508290
rect 86843 508110 86899 508166
rect 86967 508110 87023 508166
rect 87091 508110 87147 508166
rect 87215 508110 87271 508166
rect 87339 508234 87395 508290
rect 87463 508234 87519 508290
rect 87587 508234 87643 508290
rect 87711 508234 87767 508290
rect 87339 508110 87395 508166
rect 87463 508110 87519 508166
rect 87587 508110 87643 508166
rect 87711 508110 87767 508166
rect 87835 508234 87891 508290
rect 87959 508234 88015 508290
rect 88083 508234 88139 508290
rect 88207 508234 88263 508290
rect 87835 508110 87891 508166
rect 87959 508110 88015 508166
rect 88083 508110 88139 508166
rect 88207 508110 88263 508166
rect 88331 508234 88387 508290
rect 88455 508234 88511 508290
rect 88579 508234 88635 508290
rect 88703 508234 88759 508290
rect 88331 508110 88387 508166
rect 88455 508110 88511 508166
rect 88579 508110 88635 508166
rect 88703 508110 88759 508166
rect 88827 508234 88883 508290
rect 88951 508234 89007 508290
rect 89075 508234 89131 508290
rect 89199 508234 89255 508290
rect 88827 508110 88883 508166
rect 88951 508110 89007 508166
rect 89075 508110 89131 508166
rect 89199 508110 89255 508166
rect 89323 508234 89379 508290
rect 89447 508234 89503 508290
rect 89571 508234 89627 508290
rect 89695 508234 89751 508290
rect 89323 508110 89379 508166
rect 89447 508110 89503 508166
rect 89571 508110 89627 508166
rect 89695 508110 89751 508166
rect 89819 508234 89875 508290
rect 89943 508234 89999 508290
rect 90067 508234 90123 508290
rect 90191 508234 90247 508290
rect 89819 508110 89875 508166
rect 89943 508110 89999 508166
rect 90067 508110 90123 508166
rect 90191 508110 90247 508166
rect 90315 508234 90371 508290
rect 90439 508234 90495 508290
rect 90563 508234 90619 508290
rect 90687 508234 90743 508290
rect 90315 508110 90371 508166
rect 90439 508110 90495 508166
rect 90563 508110 90619 508166
rect 90687 508110 90743 508166
rect 90811 508234 90867 508290
rect 90935 508234 90991 508290
rect 91059 508234 91115 508290
rect 91183 508234 91239 508290
rect 90811 508110 90867 508166
rect 90935 508110 90991 508166
rect 91059 508110 91115 508166
rect 91183 508110 91239 508166
rect 91307 508234 91363 508290
rect 91431 508234 91487 508290
rect 91555 508234 91611 508290
rect 91679 508234 91735 508290
rect 91307 508110 91363 508166
rect 91431 508110 91487 508166
rect 91555 508110 91611 508166
rect 91679 508110 91735 508166
rect 91803 508234 91859 508290
rect 91927 508234 91983 508290
rect 92051 508234 92107 508290
rect 92175 508234 92231 508290
rect 91803 508110 91859 508166
rect 91927 508110 91983 508166
rect 92051 508110 92107 508166
rect 92175 508110 92231 508166
rect 92299 508234 92355 508290
rect 92423 508234 92479 508290
rect 92547 508234 92603 508290
rect 92671 508234 92727 508290
rect 92299 508110 92355 508166
rect 92423 508110 92479 508166
rect 92547 508110 92603 508166
rect 92671 508110 92727 508166
rect 92795 508234 92851 508290
rect 92919 508234 92975 508290
rect 93043 508234 93099 508290
rect 93167 508234 93223 508290
rect 92795 508110 92851 508166
rect 92919 508110 92975 508166
rect 93043 508110 93099 508166
rect 93167 508110 93223 508166
rect 93291 508234 93347 508290
rect 93415 508234 93471 508290
rect 93539 508234 93595 508290
rect 93663 508234 93719 508290
rect 93291 508110 93347 508166
rect 93415 508110 93471 508166
rect 93539 508110 93595 508166
rect 93663 508110 93719 508166
rect 159114 508294 159170 508350
rect 159238 508294 159294 508350
rect 159362 508294 159418 508350
rect 159486 508294 159542 508350
rect 159114 508170 159170 508226
rect 159238 508170 159294 508226
rect 159362 508170 159418 508226
rect 159486 508170 159542 508226
rect 159114 508046 159170 508102
rect 159238 508046 159294 508102
rect 159362 508046 159418 508102
rect 159486 508046 159542 508102
rect 159114 507922 159170 507978
rect 159238 507922 159294 507978
rect 159362 507922 159418 507978
rect 159486 507922 159542 507978
rect 85062 507835 85118 507891
rect 85166 507835 85222 507891
rect 85270 507835 85326 507891
rect 85374 507835 85430 507891
rect 85478 507835 85534 507891
rect 85582 507835 85638 507891
rect 85686 507835 85742 507891
rect 85790 507835 85846 507891
rect 85894 507835 85950 507891
rect 85998 507835 86054 507891
rect 86102 507835 86158 507891
rect 86206 507835 86262 507891
rect 86310 507835 86366 507891
rect 86414 507835 86470 507891
rect 86518 507835 86574 507891
rect 86622 507835 86678 507891
rect 86726 507835 86782 507891
rect 86830 507835 86886 507891
rect 86934 507835 86990 507891
rect 87038 507835 87094 507891
rect 87142 507835 87198 507891
rect 87246 507835 87302 507891
rect 87350 507835 87406 507891
rect 87454 507835 87510 507891
rect 87558 507835 87614 507891
rect 87662 507835 87718 507891
rect 87766 507835 87822 507891
rect 87870 507835 87926 507891
rect 87974 507835 88030 507891
rect 88078 507835 88134 507891
rect 88182 507835 88238 507891
rect 88286 507835 88342 507891
rect 88390 507835 88446 507891
rect 88494 507835 88550 507891
rect 88598 507835 88654 507891
rect 88702 507835 88758 507891
rect 88806 507835 88862 507891
rect 88910 507835 88966 507891
rect 89014 507835 89070 507891
rect 89118 507835 89174 507891
rect 89222 507835 89278 507891
rect 89326 507835 89382 507891
rect 89430 507835 89486 507891
rect 89534 507835 89590 507891
rect 89638 507835 89694 507891
rect 89742 507835 89798 507891
rect 89846 507835 89902 507891
rect 89950 507835 90006 507891
rect 90054 507835 90110 507891
rect 90158 507835 90214 507891
rect 90262 507835 90318 507891
rect 90366 507835 90422 507891
rect 90470 507835 90526 507891
rect 90574 507835 90630 507891
rect 90678 507835 90734 507891
rect 90782 507835 90838 507891
rect 90886 507835 90942 507891
rect 90990 507835 91046 507891
rect 91094 507835 91150 507891
rect 91198 507835 91254 507891
rect 91302 507835 91358 507891
rect 91406 507835 91462 507891
rect 91510 507835 91566 507891
rect 91614 507835 91670 507891
rect 91718 507835 91774 507891
rect 91822 507835 91878 507891
rect 91926 507835 91982 507891
rect 92030 507835 92086 507891
rect 92134 507835 92190 507891
rect 92238 507835 92294 507891
rect 92342 507835 92398 507891
rect 92446 507835 92502 507891
rect 92550 507835 92606 507891
rect 92654 507835 92710 507891
rect 92758 507835 92814 507891
rect 92862 507835 92918 507891
rect 92966 507835 93022 507891
rect 93070 507835 93126 507891
rect 93174 507835 93230 507891
rect 93278 507835 93334 507891
rect 93382 507835 93438 507891
rect 39954 496294 40010 496350
rect 40078 496294 40134 496350
rect 40202 496294 40258 496350
rect 40326 496294 40382 496350
rect 39954 496170 40010 496226
rect 40078 496170 40134 496226
rect 40202 496170 40258 496226
rect 40326 496170 40382 496226
rect 39954 496046 40010 496102
rect 40078 496046 40134 496102
rect 40202 496046 40258 496102
rect 40326 496046 40382 496102
rect 39954 495922 40010 495978
rect 40078 495922 40134 495978
rect 40202 495922 40258 495978
rect 40326 495922 40382 495978
rect 39954 478294 40010 478350
rect 40078 478294 40134 478350
rect 40202 478294 40258 478350
rect 40326 478294 40382 478350
rect 39954 478170 40010 478226
rect 40078 478170 40134 478226
rect 40202 478170 40258 478226
rect 40326 478170 40382 478226
rect 39954 478046 40010 478102
rect 40078 478046 40134 478102
rect 40202 478046 40258 478102
rect 40326 478046 40382 478102
rect 39954 477922 40010 477978
rect 40078 477922 40134 477978
rect 40202 477922 40258 477978
rect 40326 477922 40382 477978
rect 39954 460294 40010 460350
rect 40078 460294 40134 460350
rect 40202 460294 40258 460350
rect 40326 460294 40382 460350
rect 39954 460170 40010 460226
rect 40078 460170 40134 460226
rect 40202 460170 40258 460226
rect 40326 460170 40382 460226
rect 39954 460046 40010 460102
rect 40078 460046 40134 460102
rect 40202 460046 40258 460102
rect 40326 460046 40382 460102
rect 39954 459922 40010 459978
rect 40078 459922 40134 459978
rect 40202 459922 40258 459978
rect 40326 459922 40382 459978
rect 39954 442294 40010 442350
rect 40078 442294 40134 442350
rect 40202 442294 40258 442350
rect 40326 442294 40382 442350
rect 39954 442170 40010 442226
rect 40078 442170 40134 442226
rect 40202 442170 40258 442226
rect 40326 442170 40382 442226
rect 39954 442046 40010 442102
rect 40078 442046 40134 442102
rect 40202 442046 40258 442102
rect 40326 442046 40382 442102
rect 39954 441922 40010 441978
rect 40078 441922 40134 441978
rect 40202 441922 40258 441978
rect 40326 441922 40382 441978
rect 39954 424294 40010 424350
rect 40078 424294 40134 424350
rect 40202 424294 40258 424350
rect 40326 424294 40382 424350
rect 39954 424170 40010 424226
rect 40078 424170 40134 424226
rect 40202 424170 40258 424226
rect 40326 424170 40382 424226
rect 39954 424046 40010 424102
rect 40078 424046 40134 424102
rect 40202 424046 40258 424102
rect 40326 424046 40382 424102
rect 39954 423922 40010 423978
rect 40078 423922 40134 423978
rect 40202 423922 40258 423978
rect 40326 423922 40382 423978
rect 63508 496357 63564 496413
rect 63632 496357 63688 496413
rect 63756 496357 63812 496413
rect 63880 496357 63936 496413
rect 64004 496357 64060 496413
rect 64128 496357 64184 496413
rect 64252 496357 64308 496413
rect 64376 496357 64432 496413
rect 64500 496357 64556 496413
rect 64624 496357 64680 496413
rect 64748 496357 64804 496413
rect 64872 496357 64928 496413
rect 64996 496357 65052 496413
rect 65120 496357 65176 496413
rect 65244 496357 65300 496413
rect 65368 496357 65424 496413
rect 65492 496357 65548 496413
rect 65616 496357 65672 496413
rect 65740 496357 65796 496413
rect 65864 496357 65920 496413
rect 65988 496357 66044 496413
rect 66112 496357 66168 496413
rect 66236 496357 66292 496413
rect 66360 496357 66416 496413
rect 66484 496357 66540 496413
rect 66608 496357 66664 496413
rect 66732 496357 66788 496413
rect 66856 496357 66912 496413
rect 66980 496357 67036 496413
rect 67104 496357 67160 496413
rect 67228 496357 67284 496413
rect 67352 496357 67408 496413
rect 67476 496357 67532 496413
rect 67600 496357 67656 496413
rect 67724 496357 67780 496413
rect 67848 496357 67904 496413
rect 67972 496357 68028 496413
rect 68096 496357 68152 496413
rect 68220 496357 68276 496413
rect 68344 496357 68400 496413
rect 68468 496357 68524 496413
rect 68592 496357 68648 496413
rect 68716 496357 68772 496413
rect 68840 496357 68896 496413
rect 68964 496357 69020 496413
rect 69088 496357 69144 496413
rect 69212 496357 69268 496413
rect 69336 496357 69392 496413
rect 63508 496233 63564 496289
rect 63632 496233 63688 496289
rect 63756 496233 63812 496289
rect 63880 496233 63936 496289
rect 64004 496233 64060 496289
rect 64128 496233 64184 496289
rect 64252 496233 64308 496289
rect 64376 496233 64432 496289
rect 64500 496233 64556 496289
rect 64624 496233 64680 496289
rect 64748 496233 64804 496289
rect 64872 496233 64928 496289
rect 64996 496233 65052 496289
rect 65120 496233 65176 496289
rect 65244 496233 65300 496289
rect 65368 496233 65424 496289
rect 65492 496233 65548 496289
rect 65616 496233 65672 496289
rect 65740 496233 65796 496289
rect 65864 496233 65920 496289
rect 65988 496233 66044 496289
rect 66112 496233 66168 496289
rect 66236 496233 66292 496289
rect 66360 496233 66416 496289
rect 66484 496233 66540 496289
rect 66608 496233 66664 496289
rect 66732 496233 66788 496289
rect 66856 496233 66912 496289
rect 66980 496233 67036 496289
rect 67104 496233 67160 496289
rect 67228 496233 67284 496289
rect 67352 496233 67408 496289
rect 67476 496233 67532 496289
rect 67600 496233 67656 496289
rect 67724 496233 67780 496289
rect 67848 496233 67904 496289
rect 67972 496233 68028 496289
rect 68096 496233 68152 496289
rect 68220 496233 68276 496289
rect 68344 496233 68400 496289
rect 68468 496233 68524 496289
rect 68592 496233 68648 496289
rect 68716 496233 68772 496289
rect 68840 496233 68896 496289
rect 68964 496233 69020 496289
rect 69088 496233 69144 496289
rect 69212 496233 69268 496289
rect 69336 496233 69392 496289
rect 63671 495947 63727 496003
rect 63795 495947 63851 496003
rect 63919 495947 63975 496003
rect 64043 495947 64099 496003
rect 64167 495947 64223 496003
rect 64291 495947 64347 496003
rect 64415 495947 64471 496003
rect 64539 495947 64595 496003
rect 64663 495947 64719 496003
rect 64787 495947 64843 496003
rect 64911 495947 64967 496003
rect 65035 495947 65091 496003
rect 65159 495947 65215 496003
rect 65283 495947 65339 496003
rect 65407 495947 65463 496003
rect 65531 495947 65587 496003
rect 65655 495947 65711 496003
rect 65779 495947 65835 496003
rect 65903 495947 65959 496003
rect 66027 495947 66083 496003
rect 66151 495947 66207 496003
rect 66275 495947 66331 496003
rect 66399 495947 66455 496003
rect 66523 495947 66579 496003
rect 66647 495947 66703 496003
rect 66771 495947 66827 496003
rect 66895 495947 66951 496003
rect 67019 495947 67075 496003
rect 67143 495947 67199 496003
rect 67267 495947 67323 496003
rect 67391 495947 67447 496003
rect 67515 495947 67571 496003
rect 67639 495947 67695 496003
rect 67763 495947 67819 496003
rect 67887 495947 67943 496003
rect 68011 495947 68067 496003
rect 68135 495947 68191 496003
rect 68259 495947 68315 496003
rect 68383 495947 68439 496003
rect 68507 495947 68563 496003
rect 68631 495947 68687 496003
rect 68755 495947 68811 496003
rect 68879 495947 68935 496003
rect 69003 495947 69059 496003
rect 69127 495947 69183 496003
rect 69251 495947 69307 496003
rect 69375 495947 69431 496003
rect 69499 495947 69555 496003
rect 69623 495947 69679 496003
rect 80593 490234 80649 490290
rect 80717 490234 80773 490290
rect 80841 490234 80897 490290
rect 80965 490234 81021 490290
rect 81089 490234 81145 490290
rect 81213 490234 81269 490290
rect 81337 490234 81393 490290
rect 81461 490234 81517 490290
rect 81585 490234 81641 490290
rect 81709 490234 81765 490290
rect 81833 490234 81889 490290
rect 81957 490234 82013 490290
rect 82081 490234 82137 490290
rect 82205 490234 82261 490290
rect 82329 490234 82385 490290
rect 82453 490234 82509 490290
rect 82577 490234 82633 490290
rect 82701 490234 82757 490290
rect 80593 490110 80649 490166
rect 80717 490110 80773 490166
rect 80841 490110 80897 490166
rect 80965 490110 81021 490166
rect 81089 490110 81145 490166
rect 81213 490110 81269 490166
rect 81337 490110 81393 490166
rect 81461 490110 81517 490166
rect 81585 490110 81641 490166
rect 81709 490110 81765 490166
rect 81833 490110 81889 490166
rect 81957 490110 82013 490166
rect 82081 490110 82137 490166
rect 82205 490110 82261 490166
rect 82329 490110 82385 490166
rect 82453 490110 82509 490166
rect 82577 490110 82633 490166
rect 82701 490110 82757 490166
rect 128394 490294 128450 490350
rect 128518 490294 128574 490350
rect 128642 490294 128698 490350
rect 128766 490294 128822 490350
rect 128394 490170 128450 490226
rect 128518 490170 128574 490226
rect 128642 490170 128698 490226
rect 128766 490170 128822 490226
rect 128394 490046 128450 490102
rect 128518 490046 128574 490102
rect 128642 490046 128698 490102
rect 128766 490046 128822 490102
rect 128394 489922 128450 489978
rect 128518 489922 128574 489978
rect 128642 489922 128698 489978
rect 128766 489922 128822 489978
rect 80457 489835 80513 489891
rect 80561 489835 80617 489891
rect 80665 489835 80721 489891
rect 80769 489835 80825 489891
rect 80873 489835 80929 489891
rect 80977 489835 81033 489891
rect 81081 489835 81137 489891
rect 81185 489835 81241 489891
rect 81289 489835 81345 489891
rect 81393 489835 81449 489891
rect 81497 489835 81553 489891
rect 81601 489835 81657 489891
rect 81705 489835 81761 489891
rect 81809 489835 81865 489891
rect 81913 489835 81969 489891
rect 82017 489835 82073 489891
rect 82121 489835 82177 489891
rect 82225 489835 82281 489891
rect 82329 489835 82385 489891
rect 82433 489835 82489 489891
rect 82537 489835 82593 489891
rect 57932 409202 57988 409258
rect 66954 472294 67010 472350
rect 67078 472294 67134 472350
rect 67202 472294 67258 472350
rect 67326 472294 67382 472350
rect 66954 472170 67010 472226
rect 67078 472170 67134 472226
rect 67202 472170 67258 472226
rect 67326 472170 67382 472226
rect 66954 472046 67010 472102
rect 67078 472046 67134 472102
rect 67202 472046 67258 472102
rect 67326 472046 67382 472102
rect 66954 471922 67010 471978
rect 67078 471922 67134 471978
rect 67202 471922 67258 471978
rect 67326 471922 67382 471978
rect 66954 454294 67010 454350
rect 67078 454294 67134 454350
rect 67202 454294 67258 454350
rect 67326 454294 67382 454350
rect 66954 454170 67010 454226
rect 67078 454170 67134 454226
rect 67202 454170 67258 454226
rect 67326 454170 67382 454226
rect 66954 454046 67010 454102
rect 67078 454046 67134 454102
rect 67202 454046 67258 454102
rect 67326 454046 67382 454102
rect 66954 453922 67010 453978
rect 67078 453922 67134 453978
rect 67202 453922 67258 453978
rect 67326 453922 67382 453978
rect 66954 436294 67010 436350
rect 67078 436294 67134 436350
rect 67202 436294 67258 436350
rect 67326 436294 67382 436350
rect 66954 436170 67010 436226
rect 67078 436170 67134 436226
rect 67202 436170 67258 436226
rect 67326 436170 67382 436226
rect 66954 436046 67010 436102
rect 67078 436046 67134 436102
rect 67202 436046 67258 436102
rect 67326 436046 67382 436102
rect 66954 435922 67010 435978
rect 67078 435922 67134 435978
rect 67202 435922 67258 435978
rect 67326 435922 67382 435978
rect 66954 418294 67010 418350
rect 67078 418294 67134 418350
rect 67202 418294 67258 418350
rect 67326 418294 67382 418350
rect 66954 418170 67010 418226
rect 67078 418170 67134 418226
rect 67202 418170 67258 418226
rect 67326 418170 67382 418226
rect 66954 418046 67010 418102
rect 67078 418046 67134 418102
rect 67202 418046 67258 418102
rect 67326 418046 67382 418102
rect 66954 417922 67010 417978
rect 67078 417922 67134 417978
rect 67202 417922 67258 417978
rect 67326 417922 67382 417978
rect 39954 406294 40010 406350
rect 40078 406294 40134 406350
rect 40202 406294 40258 406350
rect 40326 406294 40382 406350
rect 39954 406170 40010 406226
rect 40078 406170 40134 406226
rect 40202 406170 40258 406226
rect 40326 406170 40382 406226
rect 39954 406046 40010 406102
rect 40078 406046 40134 406102
rect 40202 406046 40258 406102
rect 40326 406046 40382 406102
rect 39954 405922 40010 405978
rect 40078 405922 40134 405978
rect 40202 405922 40258 405978
rect 40326 405922 40382 405978
rect 39954 388294 40010 388350
rect 40078 388294 40134 388350
rect 40202 388294 40258 388350
rect 40326 388294 40382 388350
rect 39954 388170 40010 388226
rect 40078 388170 40134 388226
rect 40202 388170 40258 388226
rect 40326 388170 40382 388226
rect 39954 388046 40010 388102
rect 40078 388046 40134 388102
rect 40202 388046 40258 388102
rect 40326 388046 40382 388102
rect 39954 387922 40010 387978
rect 40078 387922 40134 387978
rect 40202 387922 40258 387978
rect 40326 387922 40382 387978
rect 39954 370294 40010 370350
rect 40078 370294 40134 370350
rect 40202 370294 40258 370350
rect 40326 370294 40382 370350
rect 39954 370170 40010 370226
rect 40078 370170 40134 370226
rect 40202 370170 40258 370226
rect 40326 370170 40382 370226
rect 39954 370046 40010 370102
rect 40078 370046 40134 370102
rect 40202 370046 40258 370102
rect 40326 370046 40382 370102
rect 39954 369922 40010 369978
rect 40078 369922 40134 369978
rect 40202 369922 40258 369978
rect 40326 369922 40382 369978
rect 39954 352294 40010 352350
rect 40078 352294 40134 352350
rect 40202 352294 40258 352350
rect 40326 352294 40382 352350
rect 39954 352170 40010 352226
rect 40078 352170 40134 352226
rect 40202 352170 40258 352226
rect 40326 352170 40382 352226
rect 39954 352046 40010 352102
rect 40078 352046 40134 352102
rect 40202 352046 40258 352102
rect 40326 352046 40382 352102
rect 39954 351922 40010 351978
rect 40078 351922 40134 351978
rect 40202 351922 40258 351978
rect 40326 351922 40382 351978
rect 39954 334294 40010 334350
rect 40078 334294 40134 334350
rect 40202 334294 40258 334350
rect 40326 334294 40382 334350
rect 39954 334170 40010 334226
rect 40078 334170 40134 334226
rect 40202 334170 40258 334226
rect 40326 334170 40382 334226
rect 39954 334046 40010 334102
rect 40078 334046 40134 334102
rect 40202 334046 40258 334102
rect 40326 334046 40382 334102
rect 39954 333922 40010 333978
rect 40078 333922 40134 333978
rect 40202 333922 40258 333978
rect 40326 333922 40382 333978
rect 39954 316294 40010 316350
rect 40078 316294 40134 316350
rect 40202 316294 40258 316350
rect 40326 316294 40382 316350
rect 39954 316170 40010 316226
rect 40078 316170 40134 316226
rect 40202 316170 40258 316226
rect 40326 316170 40382 316226
rect 39954 316046 40010 316102
rect 40078 316046 40134 316102
rect 40202 316046 40258 316102
rect 40326 316046 40382 316102
rect 39954 315922 40010 315978
rect 40078 315922 40134 315978
rect 40202 315922 40258 315978
rect 40326 315922 40382 315978
rect 66954 400294 67010 400350
rect 67078 400294 67134 400350
rect 67202 400294 67258 400350
rect 67326 400294 67382 400350
rect 66954 400170 67010 400226
rect 67078 400170 67134 400226
rect 67202 400170 67258 400226
rect 67326 400170 67382 400226
rect 66954 400046 67010 400102
rect 67078 400046 67134 400102
rect 67202 400046 67258 400102
rect 67326 400046 67382 400102
rect 66954 399922 67010 399978
rect 67078 399922 67134 399978
rect 67202 399922 67258 399978
rect 67326 399922 67382 399978
rect 66954 382294 67010 382350
rect 67078 382294 67134 382350
rect 67202 382294 67258 382350
rect 67326 382294 67382 382350
rect 66954 382170 67010 382226
rect 67078 382170 67134 382226
rect 67202 382170 67258 382226
rect 67326 382170 67382 382226
rect 66954 382046 67010 382102
rect 67078 382046 67134 382102
rect 67202 382046 67258 382102
rect 67326 382046 67382 382102
rect 66954 381922 67010 381978
rect 67078 381922 67134 381978
rect 67202 381922 67258 381978
rect 67326 381922 67382 381978
rect 66954 364294 67010 364350
rect 67078 364294 67134 364350
rect 67202 364294 67258 364350
rect 67326 364294 67382 364350
rect 66954 364170 67010 364226
rect 67078 364170 67134 364226
rect 67202 364170 67258 364226
rect 67326 364170 67382 364226
rect 66954 364046 67010 364102
rect 67078 364046 67134 364102
rect 67202 364046 67258 364102
rect 67326 364046 67382 364102
rect 66954 363922 67010 363978
rect 67078 363922 67134 363978
rect 67202 363922 67258 363978
rect 67326 363922 67382 363978
rect 66954 346294 67010 346350
rect 67078 346294 67134 346350
rect 67202 346294 67258 346350
rect 67326 346294 67382 346350
rect 66954 346170 67010 346226
rect 67078 346170 67134 346226
rect 67202 346170 67258 346226
rect 67326 346170 67382 346226
rect 66954 346046 67010 346102
rect 67078 346046 67134 346102
rect 67202 346046 67258 346102
rect 67326 346046 67382 346102
rect 66954 345922 67010 345978
rect 67078 345922 67134 345978
rect 67202 345922 67258 345978
rect 67326 345922 67382 345978
rect 66954 328294 67010 328350
rect 67078 328294 67134 328350
rect 67202 328294 67258 328350
rect 67326 328294 67382 328350
rect 66954 328170 67010 328226
rect 67078 328170 67134 328226
rect 67202 328170 67258 328226
rect 67326 328170 67382 328226
rect 66954 328046 67010 328102
rect 67078 328046 67134 328102
rect 67202 328046 67258 328102
rect 67326 328046 67382 328102
rect 66954 327922 67010 327978
rect 67078 327922 67134 327978
rect 67202 327922 67258 327978
rect 67326 327922 67382 327978
rect 66954 310294 67010 310350
rect 67078 310294 67134 310350
rect 67202 310294 67258 310350
rect 67326 310294 67382 310350
rect 66954 310170 67010 310226
rect 67078 310170 67134 310226
rect 67202 310170 67258 310226
rect 67326 310170 67382 310226
rect 66954 310046 67010 310102
rect 67078 310046 67134 310102
rect 67202 310046 67258 310102
rect 67326 310046 67382 310102
rect 66954 309922 67010 309978
rect 67078 309922 67134 309978
rect 67202 309922 67258 309978
rect 67326 309922 67382 309978
rect 39954 298294 40010 298350
rect 40078 298294 40134 298350
rect 40202 298294 40258 298350
rect 40326 298294 40382 298350
rect 39954 298170 40010 298226
rect 40078 298170 40134 298226
rect 40202 298170 40258 298226
rect 40326 298170 40382 298226
rect 39954 298046 40010 298102
rect 40078 298046 40134 298102
rect 40202 298046 40258 298102
rect 40326 298046 40382 298102
rect 39954 297922 40010 297978
rect 40078 297922 40134 297978
rect 40202 297922 40258 297978
rect 40326 297922 40382 297978
rect 70674 478294 70730 478350
rect 70798 478294 70854 478350
rect 70922 478294 70978 478350
rect 71046 478294 71102 478350
rect 70674 478170 70730 478226
rect 70798 478170 70854 478226
rect 70922 478170 70978 478226
rect 71046 478170 71102 478226
rect 70674 478046 70730 478102
rect 70798 478046 70854 478102
rect 70922 478046 70978 478102
rect 71046 478046 71102 478102
rect 70674 477922 70730 477978
rect 70798 477922 70854 477978
rect 70922 477922 70978 477978
rect 71046 477922 71102 477978
rect 70674 460294 70730 460350
rect 70798 460294 70854 460350
rect 70922 460294 70978 460350
rect 71046 460294 71102 460350
rect 70674 460170 70730 460226
rect 70798 460170 70854 460226
rect 70922 460170 70978 460226
rect 71046 460170 71102 460226
rect 70674 460046 70730 460102
rect 70798 460046 70854 460102
rect 70922 460046 70978 460102
rect 71046 460046 71102 460102
rect 70674 459922 70730 459978
rect 70798 459922 70854 459978
rect 70922 459922 70978 459978
rect 71046 459922 71102 459978
rect 70674 442294 70730 442350
rect 70798 442294 70854 442350
rect 70922 442294 70978 442350
rect 71046 442294 71102 442350
rect 70674 442170 70730 442226
rect 70798 442170 70854 442226
rect 70922 442170 70978 442226
rect 71046 442170 71102 442226
rect 70674 442046 70730 442102
rect 70798 442046 70854 442102
rect 70922 442046 70978 442102
rect 71046 442046 71102 442102
rect 70674 441922 70730 441978
rect 70798 441922 70854 441978
rect 70922 441922 70978 441978
rect 71046 441922 71102 441978
rect 70674 424294 70730 424350
rect 70798 424294 70854 424350
rect 70922 424294 70978 424350
rect 71046 424294 71102 424350
rect 70674 424170 70730 424226
rect 70798 424170 70854 424226
rect 70922 424170 70978 424226
rect 71046 424170 71102 424226
rect 70674 424046 70730 424102
rect 70798 424046 70854 424102
rect 70922 424046 70978 424102
rect 71046 424046 71102 424102
rect 70674 423922 70730 423978
rect 70798 423922 70854 423978
rect 70922 423922 70978 423978
rect 71046 423922 71102 423978
rect 70674 406294 70730 406350
rect 70798 406294 70854 406350
rect 70922 406294 70978 406350
rect 71046 406294 71102 406350
rect 70674 406170 70730 406226
rect 70798 406170 70854 406226
rect 70922 406170 70978 406226
rect 71046 406170 71102 406226
rect 70674 406046 70730 406102
rect 70798 406046 70854 406102
rect 70922 406046 70978 406102
rect 71046 406046 71102 406102
rect 70674 405922 70730 405978
rect 70798 405922 70854 405978
rect 70922 405922 70978 405978
rect 71046 405922 71102 405978
rect 70674 388294 70730 388350
rect 70798 388294 70854 388350
rect 70922 388294 70978 388350
rect 71046 388294 71102 388350
rect 70674 388170 70730 388226
rect 70798 388170 70854 388226
rect 70922 388170 70978 388226
rect 71046 388170 71102 388226
rect 70674 388046 70730 388102
rect 70798 388046 70854 388102
rect 70922 388046 70978 388102
rect 71046 388046 71102 388102
rect 70674 387922 70730 387978
rect 70798 387922 70854 387978
rect 70922 387922 70978 387978
rect 71046 387922 71102 387978
rect 70674 370294 70730 370350
rect 70798 370294 70854 370350
rect 70922 370294 70978 370350
rect 71046 370294 71102 370350
rect 70674 370170 70730 370226
rect 70798 370170 70854 370226
rect 70922 370170 70978 370226
rect 71046 370170 71102 370226
rect 70674 370046 70730 370102
rect 70798 370046 70854 370102
rect 70922 370046 70978 370102
rect 71046 370046 71102 370102
rect 70674 369922 70730 369978
rect 70798 369922 70854 369978
rect 70922 369922 70978 369978
rect 71046 369922 71102 369978
rect 70674 352294 70730 352350
rect 70798 352294 70854 352350
rect 70922 352294 70978 352350
rect 71046 352294 71102 352350
rect 70674 352170 70730 352226
rect 70798 352170 70854 352226
rect 70922 352170 70978 352226
rect 71046 352170 71102 352226
rect 70674 352046 70730 352102
rect 70798 352046 70854 352102
rect 70922 352046 70978 352102
rect 71046 352046 71102 352102
rect 70674 351922 70730 351978
rect 70798 351922 70854 351978
rect 70922 351922 70978 351978
rect 71046 351922 71102 351978
rect 70674 334294 70730 334350
rect 70798 334294 70854 334350
rect 70922 334294 70978 334350
rect 71046 334294 71102 334350
rect 70674 334170 70730 334226
rect 70798 334170 70854 334226
rect 70922 334170 70978 334226
rect 71046 334170 71102 334226
rect 70674 334046 70730 334102
rect 70798 334046 70854 334102
rect 70922 334046 70978 334102
rect 71046 334046 71102 334102
rect 70674 333922 70730 333978
rect 70798 333922 70854 333978
rect 70922 333922 70978 333978
rect 71046 333922 71102 333978
rect 70674 316294 70730 316350
rect 70798 316294 70854 316350
rect 70922 316294 70978 316350
rect 71046 316294 71102 316350
rect 70674 316170 70730 316226
rect 70798 316170 70854 316226
rect 70922 316170 70978 316226
rect 71046 316170 71102 316226
rect 70674 316046 70730 316102
rect 70798 316046 70854 316102
rect 70922 316046 70978 316102
rect 71046 316046 71102 316102
rect 70674 315922 70730 315978
rect 70798 315922 70854 315978
rect 70922 315922 70978 315978
rect 71046 315922 71102 315978
rect 70674 298366 70730 298422
rect 70798 298366 70854 298422
rect 70922 298366 70978 298422
rect 71046 298366 71102 298422
rect 70674 298242 70730 298298
rect 70798 298242 70854 298298
rect 70922 298242 70978 298298
rect 71046 298242 71102 298298
rect 70674 298118 70730 298174
rect 70798 298118 70854 298174
rect 70922 298118 70978 298174
rect 71046 298118 71102 298174
rect 97674 472294 97730 472350
rect 97798 472294 97854 472350
rect 97922 472294 97978 472350
rect 98046 472294 98102 472350
rect 97674 472170 97730 472226
rect 97798 472170 97854 472226
rect 97922 472170 97978 472226
rect 98046 472170 98102 472226
rect 97674 472046 97730 472102
rect 97798 472046 97854 472102
rect 97922 472046 97978 472102
rect 98046 472046 98102 472102
rect 97674 471922 97730 471978
rect 97798 471922 97854 471978
rect 97922 471922 97978 471978
rect 98046 471922 98102 471978
rect 97674 454294 97730 454350
rect 97798 454294 97854 454350
rect 97922 454294 97978 454350
rect 98046 454294 98102 454350
rect 97674 454170 97730 454226
rect 97798 454170 97854 454226
rect 97922 454170 97978 454226
rect 98046 454170 98102 454226
rect 97674 454046 97730 454102
rect 97798 454046 97854 454102
rect 97922 454046 97978 454102
rect 98046 454046 98102 454102
rect 97674 453922 97730 453978
rect 97798 453922 97854 453978
rect 97922 453922 97978 453978
rect 98046 453922 98102 453978
rect 97674 436294 97730 436350
rect 97798 436294 97854 436350
rect 97922 436294 97978 436350
rect 98046 436294 98102 436350
rect 97674 436170 97730 436226
rect 97798 436170 97854 436226
rect 97922 436170 97978 436226
rect 98046 436170 98102 436226
rect 97674 436046 97730 436102
rect 97798 436046 97854 436102
rect 97922 436046 97978 436102
rect 98046 436046 98102 436102
rect 97674 435922 97730 435978
rect 97798 435922 97854 435978
rect 97922 435922 97978 435978
rect 98046 435922 98102 435978
rect 97674 418294 97730 418350
rect 97798 418294 97854 418350
rect 97922 418294 97978 418350
rect 98046 418294 98102 418350
rect 97674 418170 97730 418226
rect 97798 418170 97854 418226
rect 97922 418170 97978 418226
rect 98046 418170 98102 418226
rect 97674 418046 97730 418102
rect 97798 418046 97854 418102
rect 97922 418046 97978 418102
rect 98046 418046 98102 418102
rect 97674 417922 97730 417978
rect 97798 417922 97854 417978
rect 97922 417922 97978 417978
rect 98046 417922 98102 417978
rect 97674 400294 97730 400350
rect 97798 400294 97854 400350
rect 97922 400294 97978 400350
rect 98046 400294 98102 400350
rect 97674 400170 97730 400226
rect 97798 400170 97854 400226
rect 97922 400170 97978 400226
rect 98046 400170 98102 400226
rect 97674 400046 97730 400102
rect 97798 400046 97854 400102
rect 97922 400046 97978 400102
rect 98046 400046 98102 400102
rect 97674 399922 97730 399978
rect 97798 399922 97854 399978
rect 97922 399922 97978 399978
rect 98046 399922 98102 399978
rect 101394 478294 101450 478350
rect 101518 478294 101574 478350
rect 101642 478294 101698 478350
rect 101766 478294 101822 478350
rect 101394 478170 101450 478226
rect 101518 478170 101574 478226
rect 101642 478170 101698 478226
rect 101766 478170 101822 478226
rect 101394 478046 101450 478102
rect 101518 478046 101574 478102
rect 101642 478046 101698 478102
rect 101766 478046 101822 478102
rect 101394 477922 101450 477978
rect 101518 477922 101574 477978
rect 101642 477922 101698 477978
rect 101766 477922 101822 477978
rect 101394 460294 101450 460350
rect 101518 460294 101574 460350
rect 101642 460294 101698 460350
rect 101766 460294 101822 460350
rect 101394 460170 101450 460226
rect 101518 460170 101574 460226
rect 101642 460170 101698 460226
rect 101766 460170 101822 460226
rect 101394 460046 101450 460102
rect 101518 460046 101574 460102
rect 101642 460046 101698 460102
rect 101766 460046 101822 460102
rect 101394 459922 101450 459978
rect 101518 459922 101574 459978
rect 101642 459922 101698 459978
rect 101766 459922 101822 459978
rect 101394 442294 101450 442350
rect 101518 442294 101574 442350
rect 101642 442294 101698 442350
rect 101766 442294 101822 442350
rect 101394 442170 101450 442226
rect 101518 442170 101574 442226
rect 101642 442170 101698 442226
rect 101766 442170 101822 442226
rect 101394 442046 101450 442102
rect 101518 442046 101574 442102
rect 101642 442046 101698 442102
rect 101766 442046 101822 442102
rect 101394 441922 101450 441978
rect 101518 441922 101574 441978
rect 101642 441922 101698 441978
rect 101766 441922 101822 441978
rect 101394 424294 101450 424350
rect 101518 424294 101574 424350
rect 101642 424294 101698 424350
rect 101766 424294 101822 424350
rect 101394 424170 101450 424226
rect 101518 424170 101574 424226
rect 101642 424170 101698 424226
rect 101766 424170 101822 424226
rect 101394 424046 101450 424102
rect 101518 424046 101574 424102
rect 101642 424046 101698 424102
rect 101766 424046 101822 424102
rect 101394 423922 101450 423978
rect 101518 423922 101574 423978
rect 101642 423922 101698 423978
rect 101766 423922 101822 423978
rect 101394 406294 101450 406350
rect 101518 406294 101574 406350
rect 101642 406294 101698 406350
rect 101766 406294 101822 406350
rect 101394 406170 101450 406226
rect 101518 406170 101574 406226
rect 101642 406170 101698 406226
rect 101766 406170 101822 406226
rect 101394 406046 101450 406102
rect 101518 406046 101574 406102
rect 101642 406046 101698 406102
rect 101766 406046 101822 406102
rect 101394 405922 101450 405978
rect 101518 405922 101574 405978
rect 101642 405922 101698 405978
rect 101766 405922 101822 405978
rect 128394 472294 128450 472350
rect 128518 472294 128574 472350
rect 128642 472294 128698 472350
rect 128766 472294 128822 472350
rect 128394 472170 128450 472226
rect 128518 472170 128574 472226
rect 128642 472170 128698 472226
rect 128766 472170 128822 472226
rect 128394 472046 128450 472102
rect 128518 472046 128574 472102
rect 128642 472046 128698 472102
rect 128766 472046 128822 472102
rect 128394 471922 128450 471978
rect 128518 471922 128574 471978
rect 128642 471922 128698 471978
rect 128766 471922 128822 471978
rect 128394 454294 128450 454350
rect 128518 454294 128574 454350
rect 128642 454294 128698 454350
rect 128766 454294 128822 454350
rect 128394 454170 128450 454226
rect 128518 454170 128574 454226
rect 128642 454170 128698 454226
rect 128766 454170 128822 454226
rect 128394 454046 128450 454102
rect 128518 454046 128574 454102
rect 128642 454046 128698 454102
rect 128766 454046 128822 454102
rect 128394 453922 128450 453978
rect 128518 453922 128574 453978
rect 128642 453922 128698 453978
rect 128766 453922 128822 453978
rect 128394 436294 128450 436350
rect 128518 436294 128574 436350
rect 128642 436294 128698 436350
rect 128766 436294 128822 436350
rect 128394 436170 128450 436226
rect 128518 436170 128574 436226
rect 128642 436170 128698 436226
rect 128766 436170 128822 436226
rect 128394 436046 128450 436102
rect 128518 436046 128574 436102
rect 128642 436046 128698 436102
rect 128766 436046 128822 436102
rect 128394 435922 128450 435978
rect 128518 435922 128574 435978
rect 128642 435922 128698 435978
rect 128766 435922 128822 435978
rect 128394 418294 128450 418350
rect 128518 418294 128574 418350
rect 128642 418294 128698 418350
rect 128766 418294 128822 418350
rect 128394 418170 128450 418226
rect 128518 418170 128574 418226
rect 128642 418170 128698 418226
rect 128766 418170 128822 418226
rect 128394 418046 128450 418102
rect 128518 418046 128574 418102
rect 128642 418046 128698 418102
rect 128766 418046 128822 418102
rect 128394 417922 128450 417978
rect 128518 417922 128574 417978
rect 128642 417922 128698 417978
rect 128766 417922 128822 417978
rect 128394 400294 128450 400350
rect 128518 400294 128574 400350
rect 128642 400294 128698 400350
rect 128766 400294 128822 400350
rect 128394 400170 128450 400226
rect 128518 400170 128574 400226
rect 128642 400170 128698 400226
rect 128766 400170 128822 400226
rect 128394 400046 128450 400102
rect 128518 400046 128574 400102
rect 128642 400046 128698 400102
rect 128766 400046 128822 400102
rect 128394 399922 128450 399978
rect 128518 399922 128574 399978
rect 128642 399922 128698 399978
rect 128766 399922 128822 399978
rect 101394 388294 101450 388350
rect 101518 388294 101574 388350
rect 101642 388294 101698 388350
rect 101766 388294 101822 388350
rect 101394 388170 101450 388226
rect 101518 388170 101574 388226
rect 101642 388170 101698 388226
rect 101766 388170 101822 388226
rect 101394 388046 101450 388102
rect 101518 388046 101574 388102
rect 101642 388046 101698 388102
rect 101766 388046 101822 388102
rect 101394 387922 101450 387978
rect 101518 387922 101574 387978
rect 101642 387922 101698 387978
rect 101766 387922 101822 387978
rect 97674 382294 97730 382350
rect 97798 382294 97854 382350
rect 97922 382294 97978 382350
rect 98046 382294 98102 382350
rect 97674 382170 97730 382226
rect 97798 382170 97854 382226
rect 97922 382170 97978 382226
rect 98046 382170 98102 382226
rect 97674 382046 97730 382102
rect 97798 382046 97854 382102
rect 97922 382046 97978 382102
rect 98046 382046 98102 382102
rect 97674 381922 97730 381978
rect 97798 381922 97854 381978
rect 97922 381922 97978 381978
rect 98046 381922 98102 381978
rect 97674 364294 97730 364350
rect 97798 364294 97854 364350
rect 97922 364294 97978 364350
rect 98046 364294 98102 364350
rect 97674 364170 97730 364226
rect 97798 364170 97854 364226
rect 97922 364170 97978 364226
rect 98046 364170 98102 364226
rect 97674 364046 97730 364102
rect 97798 364046 97854 364102
rect 97922 364046 97978 364102
rect 98046 364046 98102 364102
rect 97674 363922 97730 363978
rect 97798 363922 97854 363978
rect 97922 363922 97978 363978
rect 98046 363922 98102 363978
rect 97674 346294 97730 346350
rect 97798 346294 97854 346350
rect 97922 346294 97978 346350
rect 98046 346294 98102 346350
rect 97674 346170 97730 346226
rect 97798 346170 97854 346226
rect 97922 346170 97978 346226
rect 98046 346170 98102 346226
rect 97674 346046 97730 346102
rect 97798 346046 97854 346102
rect 97922 346046 97978 346102
rect 98046 346046 98102 346102
rect 97674 345922 97730 345978
rect 97798 345922 97854 345978
rect 97922 345922 97978 345978
rect 98046 345922 98102 345978
rect 97674 328294 97730 328350
rect 97798 328294 97854 328350
rect 97922 328294 97978 328350
rect 98046 328294 98102 328350
rect 97674 328170 97730 328226
rect 97798 328170 97854 328226
rect 97922 328170 97978 328226
rect 98046 328170 98102 328226
rect 97674 328046 97730 328102
rect 97798 328046 97854 328102
rect 97922 328046 97978 328102
rect 98046 328046 98102 328102
rect 97674 327922 97730 327978
rect 97798 327922 97854 327978
rect 97922 327922 97978 327978
rect 98046 327922 98102 327978
rect 97674 310294 97730 310350
rect 97798 310294 97854 310350
rect 97922 310294 97978 310350
rect 98046 310294 98102 310350
rect 97674 310170 97730 310226
rect 97798 310170 97854 310226
rect 97922 310170 97978 310226
rect 98046 310170 98102 310226
rect 97674 310046 97730 310102
rect 97798 310046 97854 310102
rect 97922 310046 97978 310102
rect 98046 310046 98102 310102
rect 97674 309922 97730 309978
rect 97798 309922 97854 309978
rect 97922 309922 97978 309978
rect 98046 309922 98102 309978
rect 44518 292294 44574 292350
rect 44642 292294 44698 292350
rect 44518 292170 44574 292226
rect 44642 292170 44698 292226
rect 44518 292046 44574 292102
rect 44642 292046 44698 292102
rect 44518 291922 44574 291978
rect 44642 291922 44698 291978
rect 39954 280294 40010 280350
rect 40078 280294 40134 280350
rect 40202 280294 40258 280350
rect 40326 280294 40382 280350
rect 39954 280170 40010 280226
rect 40078 280170 40134 280226
rect 40202 280170 40258 280226
rect 40326 280170 40382 280226
rect 39954 280046 40010 280102
rect 40078 280046 40134 280102
rect 40202 280046 40258 280102
rect 40326 280046 40382 280102
rect 39954 279922 40010 279978
rect 40078 279922 40134 279978
rect 40202 279922 40258 279978
rect 40326 279922 40382 279978
rect 44518 274294 44574 274350
rect 44642 274294 44698 274350
rect 44518 274170 44574 274226
rect 44642 274170 44698 274226
rect 44518 274046 44574 274102
rect 44642 274046 44698 274102
rect 44518 273922 44574 273978
rect 44642 273922 44698 273978
rect 39954 262294 40010 262350
rect 40078 262294 40134 262350
rect 40202 262294 40258 262350
rect 40326 262294 40382 262350
rect 39954 262170 40010 262226
rect 40078 262170 40134 262226
rect 40202 262170 40258 262226
rect 40326 262170 40382 262226
rect 39954 262046 40010 262102
rect 40078 262046 40134 262102
rect 40202 262046 40258 262102
rect 40326 262046 40382 262102
rect 39954 261922 40010 261978
rect 40078 261922 40134 261978
rect 40202 261922 40258 261978
rect 40326 261922 40382 261978
rect 44518 256294 44574 256350
rect 44642 256294 44698 256350
rect 44518 256170 44574 256226
rect 44642 256170 44698 256226
rect 44518 256046 44574 256102
rect 44642 256046 44698 256102
rect 44518 255922 44574 255978
rect 44642 255922 44698 255978
rect 39954 244294 40010 244350
rect 40078 244294 40134 244350
rect 40202 244294 40258 244350
rect 40326 244294 40382 244350
rect 39954 244170 40010 244226
rect 40078 244170 40134 244226
rect 40202 244170 40258 244226
rect 40326 244170 40382 244226
rect 39954 244046 40010 244102
rect 40078 244046 40134 244102
rect 40202 244046 40258 244102
rect 40326 244046 40382 244102
rect 39954 243922 40010 243978
rect 40078 243922 40134 243978
rect 40202 243922 40258 243978
rect 40326 243922 40382 243978
rect 46172 247022 46228 247078
rect 39954 226294 40010 226350
rect 40078 226294 40134 226350
rect 40202 226294 40258 226350
rect 40326 226294 40382 226350
rect 39954 226170 40010 226226
rect 40078 226170 40134 226226
rect 40202 226170 40258 226226
rect 40326 226170 40382 226226
rect 39954 226046 40010 226102
rect 40078 226046 40134 226102
rect 40202 226046 40258 226102
rect 40326 226046 40382 226102
rect 39954 225922 40010 225978
rect 40078 225922 40134 225978
rect 40202 225922 40258 225978
rect 40326 225922 40382 225978
rect 39954 208294 40010 208350
rect 40078 208294 40134 208350
rect 40202 208294 40258 208350
rect 40326 208294 40382 208350
rect 39954 208170 40010 208226
rect 40078 208170 40134 208226
rect 40202 208170 40258 208226
rect 40326 208170 40382 208226
rect 39954 208046 40010 208102
rect 40078 208046 40134 208102
rect 40202 208046 40258 208102
rect 40326 208046 40382 208102
rect 39954 207922 40010 207978
rect 40078 207922 40134 207978
rect 40202 207922 40258 207978
rect 40326 207922 40382 207978
rect 44518 202294 44574 202350
rect 44642 202294 44698 202350
rect 44518 202170 44574 202226
rect 44642 202170 44698 202226
rect 44518 202046 44574 202102
rect 44642 202046 44698 202102
rect 44518 201922 44574 201978
rect 44642 201922 44698 201978
rect 39954 190294 40010 190350
rect 40078 190294 40134 190350
rect 40202 190294 40258 190350
rect 40326 190294 40382 190350
rect 39954 190170 40010 190226
rect 40078 190170 40134 190226
rect 40202 190170 40258 190226
rect 40326 190170 40382 190226
rect 39954 190046 40010 190102
rect 40078 190046 40134 190102
rect 40202 190046 40258 190102
rect 40326 190046 40382 190102
rect 39954 189922 40010 189978
rect 40078 189922 40134 189978
rect 40202 189922 40258 189978
rect 40326 189922 40382 189978
rect 44518 184294 44574 184350
rect 44642 184294 44698 184350
rect 44518 184170 44574 184226
rect 44642 184170 44698 184226
rect 44518 184046 44574 184102
rect 44642 184046 44698 184102
rect 44518 183922 44574 183978
rect 44642 183922 44698 183978
rect 39954 172294 40010 172350
rect 40078 172294 40134 172350
rect 40202 172294 40258 172350
rect 40326 172294 40382 172350
rect 39954 172170 40010 172226
rect 40078 172170 40134 172226
rect 40202 172170 40258 172226
rect 40326 172170 40382 172226
rect 39954 172046 40010 172102
rect 40078 172046 40134 172102
rect 40202 172046 40258 172102
rect 40326 172046 40382 172102
rect 39954 171922 40010 171978
rect 40078 171922 40134 171978
rect 40202 171922 40258 171978
rect 40326 171922 40382 171978
rect 44518 166294 44574 166350
rect 44642 166294 44698 166350
rect 44518 166170 44574 166226
rect 44642 166170 44698 166226
rect 44518 166046 44574 166102
rect 44642 166046 44698 166102
rect 44518 165922 44574 165978
rect 44642 165922 44698 165978
rect 39954 154294 40010 154350
rect 40078 154294 40134 154350
rect 40202 154294 40258 154350
rect 40326 154294 40382 154350
rect 39954 154170 40010 154226
rect 40078 154170 40134 154226
rect 40202 154170 40258 154226
rect 40326 154170 40382 154226
rect 39954 154046 40010 154102
rect 40078 154046 40134 154102
rect 40202 154046 40258 154102
rect 40326 154046 40382 154102
rect 39954 153922 40010 153978
rect 40078 153922 40134 153978
rect 40202 153922 40258 153978
rect 40326 153922 40382 153978
rect 44518 148294 44574 148350
rect 44642 148294 44698 148350
rect 44518 148170 44574 148226
rect 44642 148170 44698 148226
rect 44518 148046 44574 148102
rect 44642 148046 44698 148102
rect 44518 147922 44574 147978
rect 44642 147922 44698 147978
rect 39954 136294 40010 136350
rect 40078 136294 40134 136350
rect 40202 136294 40258 136350
rect 40326 136294 40382 136350
rect 39954 136170 40010 136226
rect 40078 136170 40134 136226
rect 40202 136170 40258 136226
rect 40326 136170 40382 136226
rect 39954 136046 40010 136102
rect 40078 136046 40134 136102
rect 40202 136046 40258 136102
rect 40326 136046 40382 136102
rect 39954 135922 40010 135978
rect 40078 135922 40134 135978
rect 40202 135922 40258 135978
rect 40326 135922 40382 135978
rect 44518 130294 44574 130350
rect 44642 130294 44698 130350
rect 44518 130170 44574 130226
rect 44642 130170 44698 130226
rect 44518 130046 44574 130102
rect 44642 130046 44698 130102
rect 44518 129922 44574 129978
rect 44642 129922 44698 129978
rect 39954 118294 40010 118350
rect 40078 118294 40134 118350
rect 40202 118294 40258 118350
rect 40326 118294 40382 118350
rect 39954 118170 40010 118226
rect 40078 118170 40134 118226
rect 40202 118170 40258 118226
rect 40326 118170 40382 118226
rect 39954 118046 40010 118102
rect 40078 118046 40134 118102
rect 40202 118046 40258 118102
rect 40326 118046 40382 118102
rect 39954 117922 40010 117978
rect 40078 117922 40134 117978
rect 40202 117922 40258 117978
rect 40326 117922 40382 117978
rect 44518 112294 44574 112350
rect 44642 112294 44698 112350
rect 44518 112170 44574 112226
rect 44642 112170 44698 112226
rect 44518 112046 44574 112102
rect 44642 112046 44698 112102
rect 44518 111922 44574 111978
rect 44642 111922 44698 111978
rect 39954 100294 40010 100350
rect 40078 100294 40134 100350
rect 40202 100294 40258 100350
rect 40326 100294 40382 100350
rect 39954 100170 40010 100226
rect 40078 100170 40134 100226
rect 40202 100170 40258 100226
rect 40326 100170 40382 100226
rect 39954 100046 40010 100102
rect 40078 100046 40134 100102
rect 40202 100046 40258 100102
rect 40326 100046 40382 100102
rect 39954 99922 40010 99978
rect 40078 99922 40134 99978
rect 40202 99922 40258 99978
rect 40326 99922 40382 99978
rect 44518 94294 44574 94350
rect 44642 94294 44698 94350
rect 44518 94170 44574 94226
rect 44642 94170 44698 94226
rect 44518 94046 44574 94102
rect 44642 94046 44698 94102
rect 44518 93922 44574 93978
rect 44642 93922 44698 93978
rect 39954 82294 40010 82350
rect 40078 82294 40134 82350
rect 40202 82294 40258 82350
rect 40326 82294 40382 82350
rect 39954 82170 40010 82226
rect 40078 82170 40134 82226
rect 40202 82170 40258 82226
rect 40326 82170 40382 82226
rect 39954 82046 40010 82102
rect 40078 82046 40134 82102
rect 40202 82046 40258 82102
rect 40326 82046 40382 82102
rect 39954 81922 40010 81978
rect 40078 81922 40134 81978
rect 40202 81922 40258 81978
rect 40326 81922 40382 81978
rect 44518 76294 44574 76350
rect 44642 76294 44698 76350
rect 44518 76170 44574 76226
rect 44642 76170 44698 76226
rect 44518 76046 44574 76102
rect 44642 76046 44698 76102
rect 44518 75922 44574 75978
rect 44642 75922 44698 75978
rect 39954 64294 40010 64350
rect 40078 64294 40134 64350
rect 40202 64294 40258 64350
rect 40326 64294 40382 64350
rect 39954 64170 40010 64226
rect 40078 64170 40134 64226
rect 40202 64170 40258 64226
rect 40326 64170 40382 64226
rect 39954 64046 40010 64102
rect 40078 64046 40134 64102
rect 40202 64046 40258 64102
rect 40326 64046 40382 64102
rect 39954 63922 40010 63978
rect 40078 63922 40134 63978
rect 40202 63922 40258 63978
rect 40326 63922 40382 63978
rect 44518 58294 44574 58350
rect 44642 58294 44698 58350
rect 44518 58170 44574 58226
rect 44642 58170 44698 58226
rect 44518 58046 44574 58102
rect 44642 58046 44698 58102
rect 44518 57922 44574 57978
rect 44642 57922 44698 57978
rect 75238 292294 75294 292350
rect 75362 292294 75418 292350
rect 75238 292170 75294 292226
rect 75362 292170 75418 292226
rect 75238 292046 75294 292102
rect 75362 292046 75418 292102
rect 75238 291922 75294 291978
rect 75362 291922 75418 291978
rect 97674 292294 97730 292350
rect 97798 292294 97854 292350
rect 97922 292294 97978 292350
rect 98046 292294 98102 292350
rect 97674 292170 97730 292226
rect 97798 292170 97854 292226
rect 97922 292170 97978 292226
rect 98046 292170 98102 292226
rect 97674 292046 97730 292102
rect 97798 292046 97854 292102
rect 97922 292046 97978 292102
rect 98046 292046 98102 292102
rect 97674 291922 97730 291978
rect 97798 291922 97854 291978
rect 97922 291922 97978 291978
rect 98046 291922 98102 291978
rect 59878 280294 59934 280350
rect 60002 280294 60058 280350
rect 59878 280170 59934 280226
rect 60002 280170 60058 280226
rect 59878 280046 59934 280102
rect 60002 280046 60058 280102
rect 59878 279922 59934 279978
rect 60002 279922 60058 279978
rect 90598 280294 90654 280350
rect 90722 280294 90778 280350
rect 90598 280170 90654 280226
rect 90722 280170 90778 280226
rect 90598 280046 90654 280102
rect 90722 280046 90778 280102
rect 90598 279922 90654 279978
rect 90722 279922 90778 279978
rect 75238 274294 75294 274350
rect 75362 274294 75418 274350
rect 75238 274170 75294 274226
rect 75362 274170 75418 274226
rect 75238 274046 75294 274102
rect 75362 274046 75418 274102
rect 75238 273922 75294 273978
rect 75362 273922 75418 273978
rect 97674 274294 97730 274350
rect 97798 274294 97854 274350
rect 97922 274294 97978 274350
rect 98046 274294 98102 274350
rect 97674 274170 97730 274226
rect 97798 274170 97854 274226
rect 97922 274170 97978 274226
rect 98046 274170 98102 274226
rect 97674 274046 97730 274102
rect 97798 274046 97854 274102
rect 97922 274046 97978 274102
rect 98046 274046 98102 274102
rect 97674 273922 97730 273978
rect 97798 273922 97854 273978
rect 97922 273922 97978 273978
rect 98046 273922 98102 273978
rect 59878 262294 59934 262350
rect 60002 262294 60058 262350
rect 59878 262170 59934 262226
rect 60002 262170 60058 262226
rect 59878 262046 59934 262102
rect 60002 262046 60058 262102
rect 59878 261922 59934 261978
rect 60002 261922 60058 261978
rect 90598 262294 90654 262350
rect 90722 262294 90778 262350
rect 90598 262170 90654 262226
rect 90722 262170 90778 262226
rect 90598 262046 90654 262102
rect 90722 262046 90778 262102
rect 90598 261922 90654 261978
rect 90722 261922 90778 261978
rect 75238 256294 75294 256350
rect 75362 256294 75418 256350
rect 75238 256170 75294 256226
rect 75362 256170 75418 256226
rect 75238 256046 75294 256102
rect 75362 256046 75418 256102
rect 75238 255922 75294 255978
rect 75362 255922 75418 255978
rect 97674 256294 97730 256350
rect 97798 256294 97854 256350
rect 97922 256294 97978 256350
rect 98046 256294 98102 256350
rect 97674 256170 97730 256226
rect 97798 256170 97854 256226
rect 97922 256170 97978 256226
rect 98046 256170 98102 256226
rect 97674 256046 97730 256102
rect 97798 256046 97854 256102
rect 97922 256046 97978 256102
rect 98046 256046 98102 256102
rect 97674 255922 97730 255978
rect 97798 255922 97854 255978
rect 97922 255922 97978 255978
rect 98046 255922 98102 255978
rect 59878 244294 59934 244350
rect 60002 244294 60058 244350
rect 59878 244170 59934 244226
rect 60002 244170 60058 244226
rect 59878 244046 59934 244102
rect 60002 244046 60058 244102
rect 59878 243922 59934 243978
rect 60002 243922 60058 243978
rect 66954 238294 67010 238350
rect 67078 238294 67134 238350
rect 67202 238294 67258 238350
rect 67326 238294 67382 238350
rect 66954 238170 67010 238226
rect 67078 238170 67134 238226
rect 67202 238170 67258 238226
rect 67326 238170 67382 238226
rect 66954 238046 67010 238102
rect 67078 238046 67134 238102
rect 67202 238046 67258 238102
rect 67326 238046 67382 238102
rect 66954 237922 67010 237978
rect 67078 237922 67134 237978
rect 67202 237922 67258 237978
rect 67326 237922 67382 237978
rect 50316 206522 50372 206578
rect 49532 164582 49588 164638
rect 39954 46294 40010 46350
rect 40078 46294 40134 46350
rect 40202 46294 40258 46350
rect 40326 46294 40382 46350
rect 39954 46170 40010 46226
rect 40078 46170 40134 46226
rect 40202 46170 40258 46226
rect 40326 46170 40382 46226
rect 39954 46046 40010 46102
rect 40078 46046 40134 46102
rect 40202 46046 40258 46102
rect 40326 46046 40382 46102
rect 39954 45922 40010 45978
rect 40078 45922 40134 45978
rect 40202 45922 40258 45978
rect 40326 45922 40382 45978
rect 39954 28294 40010 28350
rect 40078 28294 40134 28350
rect 40202 28294 40258 28350
rect 40326 28294 40382 28350
rect 39954 28170 40010 28226
rect 40078 28170 40134 28226
rect 40202 28170 40258 28226
rect 40326 28170 40382 28226
rect 39954 28046 40010 28102
rect 40078 28046 40134 28102
rect 40202 28046 40258 28102
rect 40326 28046 40382 28102
rect 39954 27922 40010 27978
rect 40078 27922 40134 27978
rect 40202 27922 40258 27978
rect 40326 27922 40382 27978
rect 39954 10294 40010 10350
rect 40078 10294 40134 10350
rect 40202 10294 40258 10350
rect 40326 10294 40382 10350
rect 39954 10170 40010 10226
rect 40078 10170 40134 10226
rect 40202 10170 40258 10226
rect 40326 10170 40382 10226
rect 39954 10046 40010 10102
rect 40078 10046 40134 10102
rect 40202 10046 40258 10102
rect 40326 10046 40382 10102
rect 39954 9922 40010 9978
rect 40078 9922 40134 9978
rect 40202 9922 40258 9978
rect 40326 9922 40382 9978
rect 66954 220294 67010 220350
rect 67078 220294 67134 220350
rect 67202 220294 67258 220350
rect 67326 220294 67382 220350
rect 66954 220170 67010 220226
rect 67078 220170 67134 220226
rect 67202 220170 67258 220226
rect 67326 220170 67382 220226
rect 66954 220046 67010 220102
rect 67078 220046 67134 220102
rect 67202 220046 67258 220102
rect 67326 220046 67382 220102
rect 66954 219922 67010 219978
rect 67078 219922 67134 219978
rect 67202 219922 67258 219978
rect 67326 219922 67382 219978
rect 70674 244294 70730 244350
rect 70798 244294 70854 244350
rect 70922 244294 70978 244350
rect 71046 244294 71102 244350
rect 70674 244170 70730 244226
rect 70798 244170 70854 244226
rect 70922 244170 70978 244226
rect 71046 244170 71102 244226
rect 70674 244046 70730 244102
rect 70798 244046 70854 244102
rect 70922 244046 70978 244102
rect 71046 244046 71102 244102
rect 70674 243922 70730 243978
rect 70798 243922 70854 243978
rect 70922 243922 70978 243978
rect 71046 243922 71102 243978
rect 90598 244294 90654 244350
rect 90722 244294 90778 244350
rect 90598 244170 90654 244226
rect 90722 244170 90778 244226
rect 90598 244046 90654 244102
rect 90722 244046 90778 244102
rect 90598 243922 90654 243978
rect 90722 243922 90778 243978
rect 97674 238294 97730 238350
rect 97798 238294 97854 238350
rect 97922 238294 97978 238350
rect 98046 238294 98102 238350
rect 76972 237662 77028 237718
rect 97674 238170 97730 238226
rect 97798 238170 97854 238226
rect 97922 238170 97978 238226
rect 98046 238170 98102 238226
rect 97674 238046 97730 238102
rect 97798 238046 97854 238102
rect 97922 238046 97978 238102
rect 98046 238046 98102 238102
rect 97674 237922 97730 237978
rect 97798 237922 97854 237978
rect 97922 237922 97978 237978
rect 98046 237922 98102 237978
rect 74956 237482 75012 237538
rect 70674 226294 70730 226350
rect 70798 226294 70854 226350
rect 70922 226294 70978 226350
rect 71046 226294 71102 226350
rect 70674 226170 70730 226226
rect 70798 226170 70854 226226
rect 70922 226170 70978 226226
rect 71046 226170 71102 226226
rect 70674 226046 70730 226102
rect 70798 226046 70854 226102
rect 70922 226046 70978 226102
rect 71046 226046 71102 226102
rect 70674 225922 70730 225978
rect 70798 225922 70854 225978
rect 70922 225922 70978 225978
rect 71046 225922 71102 225978
rect 99932 237482 99988 237538
rect 101394 370294 101450 370350
rect 101518 370294 101574 370350
rect 101642 370294 101698 370350
rect 101766 370294 101822 370350
rect 101394 370170 101450 370226
rect 101518 370170 101574 370226
rect 101642 370170 101698 370226
rect 101766 370170 101822 370226
rect 101394 370046 101450 370102
rect 101518 370046 101574 370102
rect 101642 370046 101698 370102
rect 101766 370046 101822 370102
rect 101394 369922 101450 369978
rect 101518 369922 101574 369978
rect 101642 369922 101698 369978
rect 101766 369922 101822 369978
rect 101394 352294 101450 352350
rect 101518 352294 101574 352350
rect 101642 352294 101698 352350
rect 101766 352294 101822 352350
rect 101394 352170 101450 352226
rect 101518 352170 101574 352226
rect 101642 352170 101698 352226
rect 101766 352170 101822 352226
rect 101394 352046 101450 352102
rect 101518 352046 101574 352102
rect 101642 352046 101698 352102
rect 101766 352046 101822 352102
rect 101394 351922 101450 351978
rect 101518 351922 101574 351978
rect 101642 351922 101698 351978
rect 101766 351922 101822 351978
rect 101394 334294 101450 334350
rect 101518 334294 101574 334350
rect 101642 334294 101698 334350
rect 101766 334294 101822 334350
rect 101394 334170 101450 334226
rect 101518 334170 101574 334226
rect 101642 334170 101698 334226
rect 101766 334170 101822 334226
rect 101394 334046 101450 334102
rect 101518 334046 101574 334102
rect 101642 334046 101698 334102
rect 101766 334046 101822 334102
rect 101394 333922 101450 333978
rect 101518 333922 101574 333978
rect 101642 333922 101698 333978
rect 101766 333922 101822 333978
rect 101394 316294 101450 316350
rect 101518 316294 101574 316350
rect 101642 316294 101698 316350
rect 101766 316294 101822 316350
rect 101394 316170 101450 316226
rect 101518 316170 101574 316226
rect 101642 316170 101698 316226
rect 101766 316170 101822 316226
rect 101394 316046 101450 316102
rect 101518 316046 101574 316102
rect 101642 316046 101698 316102
rect 101766 316046 101822 316102
rect 101394 315922 101450 315978
rect 101518 315922 101574 315978
rect 101642 315922 101698 315978
rect 101766 315922 101822 315978
rect 101394 298294 101450 298350
rect 101518 298294 101574 298350
rect 101642 298294 101698 298350
rect 101766 298294 101822 298350
rect 101394 298170 101450 298226
rect 101518 298170 101574 298226
rect 101642 298170 101698 298226
rect 101766 298170 101822 298226
rect 101394 298046 101450 298102
rect 101518 298046 101574 298102
rect 101642 298046 101698 298102
rect 101766 298046 101822 298102
rect 101394 297922 101450 297978
rect 101518 297922 101574 297978
rect 101642 297922 101698 297978
rect 101766 297922 101822 297978
rect 101394 280294 101450 280350
rect 101518 280294 101574 280350
rect 101642 280294 101698 280350
rect 101766 280294 101822 280350
rect 101394 280170 101450 280226
rect 101518 280170 101574 280226
rect 101642 280170 101698 280226
rect 101766 280170 101822 280226
rect 101394 280046 101450 280102
rect 101518 280046 101574 280102
rect 101642 280046 101698 280102
rect 101766 280046 101822 280102
rect 101394 279922 101450 279978
rect 101518 279922 101574 279978
rect 101642 279922 101698 279978
rect 101766 279922 101822 279978
rect 101394 262294 101450 262350
rect 101518 262294 101574 262350
rect 101642 262294 101698 262350
rect 101766 262294 101822 262350
rect 101394 262170 101450 262226
rect 101518 262170 101574 262226
rect 101642 262170 101698 262226
rect 101766 262170 101822 262226
rect 101394 262046 101450 262102
rect 101518 262046 101574 262102
rect 101642 262046 101698 262102
rect 101766 262046 101822 262102
rect 101394 261922 101450 261978
rect 101518 261922 101574 261978
rect 101642 261922 101698 261978
rect 101766 261922 101822 261978
rect 101394 244294 101450 244350
rect 101518 244294 101574 244350
rect 101642 244294 101698 244350
rect 101766 244294 101822 244350
rect 101394 244170 101450 244226
rect 101518 244170 101574 244226
rect 101642 244170 101698 244226
rect 101766 244170 101822 244226
rect 101394 244046 101450 244102
rect 101518 244046 101574 244102
rect 101642 244046 101698 244102
rect 101766 244046 101822 244102
rect 101394 243922 101450 243978
rect 101518 243922 101574 243978
rect 101642 243922 101698 243978
rect 101766 243922 101822 243978
rect 97674 220294 97730 220350
rect 97798 220294 97854 220350
rect 97922 220294 97978 220350
rect 98046 220294 98102 220350
rect 97674 220170 97730 220226
rect 97798 220170 97854 220226
rect 97922 220170 97978 220226
rect 98046 220170 98102 220226
rect 97674 220046 97730 220102
rect 97798 220046 97854 220102
rect 97922 220046 97978 220102
rect 98046 220046 98102 220102
rect 97674 219922 97730 219978
rect 97798 219922 97854 219978
rect 97922 219922 97978 219978
rect 98046 219922 98102 219978
rect 103292 237662 103348 237718
rect 128394 382294 128450 382350
rect 128518 382294 128574 382350
rect 128642 382294 128698 382350
rect 128766 382294 128822 382350
rect 128394 382170 128450 382226
rect 128518 382170 128574 382226
rect 128642 382170 128698 382226
rect 128766 382170 128822 382226
rect 128394 382046 128450 382102
rect 128518 382046 128574 382102
rect 128642 382046 128698 382102
rect 128766 382046 128822 382102
rect 128394 381922 128450 381978
rect 128518 381922 128574 381978
rect 128642 381922 128698 381978
rect 128766 381922 128822 381978
rect 128394 364294 128450 364350
rect 128518 364294 128574 364350
rect 128642 364294 128698 364350
rect 128766 364294 128822 364350
rect 128394 364170 128450 364226
rect 128518 364170 128574 364226
rect 128642 364170 128698 364226
rect 128766 364170 128822 364226
rect 128394 364046 128450 364102
rect 128518 364046 128574 364102
rect 128642 364046 128698 364102
rect 128766 364046 128822 364102
rect 128394 363922 128450 363978
rect 128518 363922 128574 363978
rect 128642 363922 128698 363978
rect 128766 363922 128822 363978
rect 128394 346294 128450 346350
rect 128518 346294 128574 346350
rect 128642 346294 128698 346350
rect 128766 346294 128822 346350
rect 128394 346170 128450 346226
rect 128518 346170 128574 346226
rect 128642 346170 128698 346226
rect 128766 346170 128822 346226
rect 128394 346046 128450 346102
rect 128518 346046 128574 346102
rect 128642 346046 128698 346102
rect 128766 346046 128822 346102
rect 128394 345922 128450 345978
rect 128518 345922 128574 345978
rect 128642 345922 128698 345978
rect 128766 345922 128822 345978
rect 128394 328294 128450 328350
rect 128518 328294 128574 328350
rect 128642 328294 128698 328350
rect 128766 328294 128822 328350
rect 128394 328170 128450 328226
rect 128518 328170 128574 328226
rect 128642 328170 128698 328226
rect 128766 328170 128822 328226
rect 128394 328046 128450 328102
rect 128518 328046 128574 328102
rect 128642 328046 128698 328102
rect 128766 328046 128822 328102
rect 128394 327922 128450 327978
rect 128518 327922 128574 327978
rect 128642 327922 128698 327978
rect 128766 327922 128822 327978
rect 128394 310294 128450 310350
rect 128518 310294 128574 310350
rect 128642 310294 128698 310350
rect 128766 310294 128822 310350
rect 128394 310170 128450 310226
rect 128518 310170 128574 310226
rect 128642 310170 128698 310226
rect 128766 310170 128822 310226
rect 128394 310046 128450 310102
rect 128518 310046 128574 310102
rect 128642 310046 128698 310102
rect 128766 310046 128822 310102
rect 128394 309922 128450 309978
rect 128518 309922 128574 309978
rect 128642 309922 128698 309978
rect 128766 309922 128822 309978
rect 128394 292294 128450 292350
rect 128518 292294 128574 292350
rect 128642 292294 128698 292350
rect 128766 292294 128822 292350
rect 128394 292170 128450 292226
rect 128518 292170 128574 292226
rect 128642 292170 128698 292226
rect 128766 292170 128822 292226
rect 128394 292046 128450 292102
rect 128518 292046 128574 292102
rect 128642 292046 128698 292102
rect 128766 292046 128822 292102
rect 128394 291922 128450 291978
rect 128518 291922 128574 291978
rect 128642 291922 128698 291978
rect 128766 291922 128822 291978
rect 128394 274294 128450 274350
rect 128518 274294 128574 274350
rect 128642 274294 128698 274350
rect 128766 274294 128822 274350
rect 128394 274170 128450 274226
rect 128518 274170 128574 274226
rect 128642 274170 128698 274226
rect 128766 274170 128822 274226
rect 128394 274046 128450 274102
rect 128518 274046 128574 274102
rect 128642 274046 128698 274102
rect 128766 274046 128822 274102
rect 128394 273922 128450 273978
rect 128518 273922 128574 273978
rect 128642 273922 128698 273978
rect 128766 273922 128822 273978
rect 128394 256294 128450 256350
rect 128518 256294 128574 256350
rect 128642 256294 128698 256350
rect 128766 256294 128822 256350
rect 128394 256170 128450 256226
rect 128518 256170 128574 256226
rect 128642 256170 128698 256226
rect 128766 256170 128822 256226
rect 128394 256046 128450 256102
rect 128518 256046 128574 256102
rect 128642 256046 128698 256102
rect 128766 256046 128822 256102
rect 128394 255922 128450 255978
rect 128518 255922 128574 255978
rect 128642 255922 128698 255978
rect 128766 255922 128822 255978
rect 128394 238294 128450 238350
rect 128518 238294 128574 238350
rect 128642 238294 128698 238350
rect 128766 238294 128822 238350
rect 128394 238170 128450 238226
rect 128518 238170 128574 238226
rect 128642 238170 128698 238226
rect 128766 238170 128822 238226
rect 128394 238046 128450 238102
rect 128518 238046 128574 238102
rect 128642 238046 128698 238102
rect 128766 238046 128822 238102
rect 128394 237922 128450 237978
rect 128518 237922 128574 237978
rect 128642 237922 128698 237978
rect 128766 237922 128822 237978
rect 101394 226294 101450 226350
rect 101518 226294 101574 226350
rect 101642 226294 101698 226350
rect 101766 226294 101822 226350
rect 101394 226170 101450 226226
rect 101518 226170 101574 226226
rect 101642 226170 101698 226226
rect 101766 226170 101822 226226
rect 101394 226046 101450 226102
rect 101518 226046 101574 226102
rect 101642 226046 101698 226102
rect 101766 226046 101822 226102
rect 101394 225922 101450 225978
rect 101518 225922 101574 225978
rect 101642 225922 101698 225978
rect 101766 225922 101822 225978
rect 128394 220294 128450 220350
rect 128518 220294 128574 220350
rect 128642 220294 128698 220350
rect 128766 220294 128822 220350
rect 128394 220170 128450 220226
rect 128518 220170 128574 220226
rect 128642 220170 128698 220226
rect 128766 220170 128822 220226
rect 128394 220046 128450 220102
rect 128518 220046 128574 220102
rect 128642 220046 128698 220102
rect 128766 220046 128822 220102
rect 128394 219922 128450 219978
rect 128518 219922 128574 219978
rect 128642 219922 128698 219978
rect 128766 219922 128822 219978
rect 132114 496294 132170 496350
rect 132238 496294 132294 496350
rect 132362 496294 132418 496350
rect 132486 496294 132542 496350
rect 132114 496170 132170 496226
rect 132238 496170 132294 496226
rect 132362 496170 132418 496226
rect 132486 496170 132542 496226
rect 132114 496046 132170 496102
rect 132238 496046 132294 496102
rect 132362 496046 132418 496102
rect 132486 496046 132542 496102
rect 132114 495922 132170 495978
rect 132238 495922 132294 495978
rect 132362 495922 132418 495978
rect 132486 495922 132542 495978
rect 132114 478294 132170 478350
rect 132238 478294 132294 478350
rect 132362 478294 132418 478350
rect 132486 478294 132542 478350
rect 132114 478170 132170 478226
rect 132238 478170 132294 478226
rect 132362 478170 132418 478226
rect 132486 478170 132542 478226
rect 132114 478046 132170 478102
rect 132238 478046 132294 478102
rect 132362 478046 132418 478102
rect 132486 478046 132542 478102
rect 132114 477922 132170 477978
rect 132238 477922 132294 477978
rect 132362 477922 132418 477978
rect 132486 477922 132542 477978
rect 159114 490294 159170 490350
rect 159238 490294 159294 490350
rect 159362 490294 159418 490350
rect 159486 490294 159542 490350
rect 159114 490170 159170 490226
rect 159238 490170 159294 490226
rect 159362 490170 159418 490226
rect 159486 490170 159542 490226
rect 159114 490046 159170 490102
rect 159238 490046 159294 490102
rect 159362 490046 159418 490102
rect 159486 490046 159542 490102
rect 159114 489922 159170 489978
rect 159238 489922 159294 489978
rect 159362 489922 159418 489978
rect 159486 489922 159542 489978
rect 132114 460294 132170 460350
rect 132238 460294 132294 460350
rect 132362 460294 132418 460350
rect 132486 460294 132542 460350
rect 132114 460170 132170 460226
rect 132238 460170 132294 460226
rect 132362 460170 132418 460226
rect 132486 460170 132542 460226
rect 132114 460046 132170 460102
rect 132238 460046 132294 460102
rect 132362 460046 132418 460102
rect 132486 460046 132542 460102
rect 132114 459922 132170 459978
rect 132238 459922 132294 459978
rect 132362 459922 132418 459978
rect 132486 459922 132542 459978
rect 132114 442294 132170 442350
rect 132238 442294 132294 442350
rect 132362 442294 132418 442350
rect 132486 442294 132542 442350
rect 132114 442170 132170 442226
rect 132238 442170 132294 442226
rect 132362 442170 132418 442226
rect 132486 442170 132542 442226
rect 132114 442046 132170 442102
rect 132238 442046 132294 442102
rect 132362 442046 132418 442102
rect 132486 442046 132542 442102
rect 132114 441922 132170 441978
rect 132238 441922 132294 441978
rect 132362 441922 132418 441978
rect 132486 441922 132542 441978
rect 132114 424294 132170 424350
rect 132238 424294 132294 424350
rect 132362 424294 132418 424350
rect 132486 424294 132542 424350
rect 132114 424170 132170 424226
rect 132238 424170 132294 424226
rect 132362 424170 132418 424226
rect 132486 424170 132542 424226
rect 132114 424046 132170 424102
rect 132238 424046 132294 424102
rect 132362 424046 132418 424102
rect 132486 424046 132542 424102
rect 132114 423922 132170 423978
rect 132238 423922 132294 423978
rect 132362 423922 132418 423978
rect 132486 423922 132542 423978
rect 132114 406294 132170 406350
rect 132238 406294 132294 406350
rect 132362 406294 132418 406350
rect 132486 406294 132542 406350
rect 132114 406170 132170 406226
rect 132238 406170 132294 406226
rect 132362 406170 132418 406226
rect 132486 406170 132542 406226
rect 132114 406046 132170 406102
rect 132238 406046 132294 406102
rect 132362 406046 132418 406102
rect 132486 406046 132542 406102
rect 132114 405922 132170 405978
rect 132238 405922 132294 405978
rect 132362 405922 132418 405978
rect 132486 405922 132542 405978
rect 132114 388294 132170 388350
rect 132238 388294 132294 388350
rect 132362 388294 132418 388350
rect 132486 388294 132542 388350
rect 132114 388170 132170 388226
rect 132238 388170 132294 388226
rect 132362 388170 132418 388226
rect 132486 388170 132542 388226
rect 132114 388046 132170 388102
rect 132238 388046 132294 388102
rect 132362 388046 132418 388102
rect 132486 388046 132542 388102
rect 132114 387922 132170 387978
rect 132238 387922 132294 387978
rect 132362 387922 132418 387978
rect 132486 387922 132542 387978
rect 132114 370294 132170 370350
rect 132238 370294 132294 370350
rect 132362 370294 132418 370350
rect 132486 370294 132542 370350
rect 132114 370170 132170 370226
rect 132238 370170 132294 370226
rect 132362 370170 132418 370226
rect 132486 370170 132542 370226
rect 132114 370046 132170 370102
rect 132238 370046 132294 370102
rect 132362 370046 132418 370102
rect 132486 370046 132542 370102
rect 132114 369922 132170 369978
rect 132238 369922 132294 369978
rect 132362 369922 132418 369978
rect 132486 369922 132542 369978
rect 132114 352294 132170 352350
rect 132238 352294 132294 352350
rect 132362 352294 132418 352350
rect 132486 352294 132542 352350
rect 132114 352170 132170 352226
rect 132238 352170 132294 352226
rect 132362 352170 132418 352226
rect 132486 352170 132542 352226
rect 132114 352046 132170 352102
rect 132238 352046 132294 352102
rect 132362 352046 132418 352102
rect 132486 352046 132542 352102
rect 132114 351922 132170 351978
rect 132238 351922 132294 351978
rect 132362 351922 132418 351978
rect 132486 351922 132542 351978
rect 132114 334294 132170 334350
rect 132238 334294 132294 334350
rect 132362 334294 132418 334350
rect 132486 334294 132542 334350
rect 132114 334170 132170 334226
rect 132238 334170 132294 334226
rect 132362 334170 132418 334226
rect 132486 334170 132542 334226
rect 132114 334046 132170 334102
rect 132238 334046 132294 334102
rect 132362 334046 132418 334102
rect 132486 334046 132542 334102
rect 132114 333922 132170 333978
rect 132238 333922 132294 333978
rect 132362 333922 132418 333978
rect 132486 333922 132542 333978
rect 132114 316294 132170 316350
rect 132238 316294 132294 316350
rect 132362 316294 132418 316350
rect 132486 316294 132542 316350
rect 132114 316170 132170 316226
rect 132238 316170 132294 316226
rect 132362 316170 132418 316226
rect 132486 316170 132542 316226
rect 132114 316046 132170 316102
rect 132238 316046 132294 316102
rect 132362 316046 132418 316102
rect 132486 316046 132542 316102
rect 132114 315922 132170 315978
rect 132238 315922 132294 315978
rect 132362 315922 132418 315978
rect 132486 315922 132542 315978
rect 132114 298294 132170 298350
rect 132238 298294 132294 298350
rect 132362 298294 132418 298350
rect 132486 298294 132542 298350
rect 132114 298170 132170 298226
rect 132238 298170 132294 298226
rect 132362 298170 132418 298226
rect 132486 298170 132542 298226
rect 132114 298046 132170 298102
rect 132238 298046 132294 298102
rect 132362 298046 132418 298102
rect 132486 298046 132542 298102
rect 132114 297922 132170 297978
rect 132238 297922 132294 297978
rect 132362 297922 132418 297978
rect 132486 297922 132542 297978
rect 159114 472294 159170 472350
rect 159238 472294 159294 472350
rect 159362 472294 159418 472350
rect 159486 472294 159542 472350
rect 159114 472170 159170 472226
rect 159238 472170 159294 472226
rect 159362 472170 159418 472226
rect 159486 472170 159542 472226
rect 159114 472046 159170 472102
rect 159238 472046 159294 472102
rect 159362 472046 159418 472102
rect 159486 472046 159542 472102
rect 159114 471922 159170 471978
rect 159238 471922 159294 471978
rect 159362 471922 159418 471978
rect 159486 471922 159542 471978
rect 162834 598116 162890 598172
rect 162958 598116 163014 598172
rect 163082 598116 163138 598172
rect 163206 598116 163262 598172
rect 162834 597992 162890 598048
rect 162958 597992 163014 598048
rect 163082 597992 163138 598048
rect 163206 597992 163262 598048
rect 162834 597868 162890 597924
rect 162958 597868 163014 597924
rect 163082 597868 163138 597924
rect 163206 597868 163262 597924
rect 162834 597744 162890 597800
rect 162958 597744 163014 597800
rect 163082 597744 163138 597800
rect 163206 597744 163262 597800
rect 162834 586294 162890 586350
rect 162958 586294 163014 586350
rect 163082 586294 163138 586350
rect 163206 586294 163262 586350
rect 162834 586170 162890 586226
rect 162958 586170 163014 586226
rect 163082 586170 163138 586226
rect 163206 586170 163262 586226
rect 162834 586046 162890 586102
rect 162958 586046 163014 586102
rect 163082 586046 163138 586102
rect 163206 586046 163262 586102
rect 162834 585922 162890 585978
rect 162958 585922 163014 585978
rect 163082 585922 163138 585978
rect 163206 585922 163262 585978
rect 162834 568294 162890 568350
rect 162958 568294 163014 568350
rect 163082 568294 163138 568350
rect 163206 568294 163262 568350
rect 162834 568170 162890 568226
rect 162958 568170 163014 568226
rect 163082 568170 163138 568226
rect 163206 568170 163262 568226
rect 162834 568046 162890 568102
rect 162958 568046 163014 568102
rect 163082 568046 163138 568102
rect 163206 568046 163262 568102
rect 162834 567922 162890 567978
rect 162958 567922 163014 567978
rect 163082 567922 163138 567978
rect 163206 567922 163262 567978
rect 189834 597156 189890 597212
rect 189958 597156 190014 597212
rect 190082 597156 190138 597212
rect 190206 597156 190262 597212
rect 189834 597032 189890 597088
rect 189958 597032 190014 597088
rect 190082 597032 190138 597088
rect 190206 597032 190262 597088
rect 189834 596908 189890 596964
rect 189958 596908 190014 596964
rect 190082 596908 190138 596964
rect 190206 596908 190262 596964
rect 189834 596784 189890 596840
rect 189958 596784 190014 596840
rect 190082 596784 190138 596840
rect 190206 596784 190262 596840
rect 193554 598116 193610 598172
rect 193678 598116 193734 598172
rect 193802 598116 193858 598172
rect 193926 598116 193982 598172
rect 193554 597992 193610 598048
rect 193678 597992 193734 598048
rect 193802 597992 193858 598048
rect 193926 597992 193982 598048
rect 193554 597868 193610 597924
rect 193678 597868 193734 597924
rect 193802 597868 193858 597924
rect 193926 597868 193982 597924
rect 193554 597744 193610 597800
rect 193678 597744 193734 597800
rect 193802 597744 193858 597800
rect 193926 597744 193982 597800
rect 189834 580294 189890 580350
rect 189958 580294 190014 580350
rect 190082 580294 190138 580350
rect 190206 580294 190262 580350
rect 189834 580170 189890 580226
rect 189958 580170 190014 580226
rect 190082 580170 190138 580226
rect 190206 580170 190262 580226
rect 189834 580046 189890 580102
rect 189958 580046 190014 580102
rect 190082 580046 190138 580102
rect 190206 580046 190262 580102
rect 189834 579922 189890 579978
rect 189958 579922 190014 579978
rect 190082 579922 190138 579978
rect 190206 579922 190262 579978
rect 162834 550294 162890 550350
rect 162958 550294 163014 550350
rect 163082 550294 163138 550350
rect 163206 550294 163262 550350
rect 162834 550170 162890 550226
rect 162958 550170 163014 550226
rect 163082 550170 163138 550226
rect 163206 550170 163262 550226
rect 162834 550046 162890 550102
rect 162958 550046 163014 550102
rect 163082 550046 163138 550102
rect 163206 550046 163262 550102
rect 162834 549922 162890 549978
rect 162958 549922 163014 549978
rect 163082 549922 163138 549978
rect 163206 549922 163262 549978
rect 162834 532294 162890 532350
rect 162958 532294 163014 532350
rect 163082 532294 163138 532350
rect 163206 532294 163262 532350
rect 162834 532170 162890 532226
rect 162958 532170 163014 532226
rect 163082 532170 163138 532226
rect 163206 532170 163262 532226
rect 162834 532046 162890 532102
rect 162958 532046 163014 532102
rect 163082 532046 163138 532102
rect 163206 532046 163262 532102
rect 162834 531922 162890 531978
rect 162958 531922 163014 531978
rect 163082 531922 163138 531978
rect 163206 531922 163262 531978
rect 162834 514294 162890 514350
rect 162958 514294 163014 514350
rect 163082 514294 163138 514350
rect 163206 514294 163262 514350
rect 162834 514170 162890 514226
rect 162958 514170 163014 514226
rect 163082 514170 163138 514226
rect 163206 514170 163262 514226
rect 162834 514046 162890 514102
rect 162958 514046 163014 514102
rect 163082 514046 163138 514102
rect 163206 514046 163262 514102
rect 162834 513922 162890 513978
rect 162958 513922 163014 513978
rect 163082 513922 163138 513978
rect 163206 513922 163262 513978
rect 162834 496294 162890 496350
rect 162958 496294 163014 496350
rect 163082 496294 163138 496350
rect 163206 496294 163262 496350
rect 162834 496170 162890 496226
rect 162958 496170 163014 496226
rect 163082 496170 163138 496226
rect 163206 496170 163262 496226
rect 162834 496046 162890 496102
rect 162958 496046 163014 496102
rect 163082 496046 163138 496102
rect 163206 496046 163262 496102
rect 162834 495922 162890 495978
rect 162958 495922 163014 495978
rect 163082 495922 163138 495978
rect 163206 495922 163262 495978
rect 162834 478294 162890 478350
rect 162958 478294 163014 478350
rect 163082 478294 163138 478350
rect 163206 478294 163262 478350
rect 162834 478170 162890 478226
rect 162958 478170 163014 478226
rect 163082 478170 163138 478226
rect 163206 478170 163262 478226
rect 162834 478046 162890 478102
rect 162958 478046 163014 478102
rect 163082 478046 163138 478102
rect 163206 478046 163262 478102
rect 162834 477922 162890 477978
rect 162958 477922 163014 477978
rect 163082 477922 163138 477978
rect 163206 477922 163262 477978
rect 159114 454294 159170 454350
rect 159238 454294 159294 454350
rect 159362 454294 159418 454350
rect 159486 454294 159542 454350
rect 159114 454170 159170 454226
rect 159238 454170 159294 454226
rect 159362 454170 159418 454226
rect 159486 454170 159542 454226
rect 159114 454046 159170 454102
rect 159238 454046 159294 454102
rect 159362 454046 159418 454102
rect 159486 454046 159542 454102
rect 159114 453922 159170 453978
rect 159238 453922 159294 453978
rect 159362 453922 159418 453978
rect 159486 453922 159542 453978
rect 159114 436294 159170 436350
rect 159238 436294 159294 436350
rect 159362 436294 159418 436350
rect 159486 436294 159542 436350
rect 159114 436170 159170 436226
rect 159238 436170 159294 436226
rect 159362 436170 159418 436226
rect 159486 436170 159542 436226
rect 159114 436046 159170 436102
rect 159238 436046 159294 436102
rect 159362 436046 159418 436102
rect 159486 436046 159542 436102
rect 159114 435922 159170 435978
rect 159238 435922 159294 435978
rect 159362 435922 159418 435978
rect 159486 435922 159542 435978
rect 159114 418294 159170 418350
rect 159238 418294 159294 418350
rect 159362 418294 159418 418350
rect 159486 418294 159542 418350
rect 159114 418170 159170 418226
rect 159238 418170 159294 418226
rect 159362 418170 159418 418226
rect 159486 418170 159542 418226
rect 159114 418046 159170 418102
rect 159238 418046 159294 418102
rect 159362 418046 159418 418102
rect 159486 418046 159542 418102
rect 159114 417922 159170 417978
rect 159238 417922 159294 417978
rect 159362 417922 159418 417978
rect 159486 417922 159542 417978
rect 159114 400294 159170 400350
rect 159238 400294 159294 400350
rect 159362 400294 159418 400350
rect 159486 400294 159542 400350
rect 159114 400170 159170 400226
rect 159238 400170 159294 400226
rect 159362 400170 159418 400226
rect 159486 400170 159542 400226
rect 159114 400046 159170 400102
rect 159238 400046 159294 400102
rect 159362 400046 159418 400102
rect 159486 400046 159542 400102
rect 159114 399922 159170 399978
rect 159238 399922 159294 399978
rect 159362 399922 159418 399978
rect 159486 399922 159542 399978
rect 159114 382294 159170 382350
rect 159238 382294 159294 382350
rect 159362 382294 159418 382350
rect 159486 382294 159542 382350
rect 159114 382170 159170 382226
rect 159238 382170 159294 382226
rect 159362 382170 159418 382226
rect 159486 382170 159542 382226
rect 159114 382046 159170 382102
rect 159238 382046 159294 382102
rect 159362 382046 159418 382102
rect 159486 382046 159542 382102
rect 159114 381922 159170 381978
rect 159238 381922 159294 381978
rect 159362 381922 159418 381978
rect 159486 381922 159542 381978
rect 159114 364294 159170 364350
rect 159238 364294 159294 364350
rect 159362 364294 159418 364350
rect 159486 364294 159542 364350
rect 159114 364170 159170 364226
rect 159238 364170 159294 364226
rect 159362 364170 159418 364226
rect 159486 364170 159542 364226
rect 159114 364046 159170 364102
rect 159238 364046 159294 364102
rect 159362 364046 159418 364102
rect 159486 364046 159542 364102
rect 159114 363922 159170 363978
rect 159238 363922 159294 363978
rect 159362 363922 159418 363978
rect 159486 363922 159542 363978
rect 154518 346294 154574 346350
rect 154642 346294 154698 346350
rect 154518 346170 154574 346226
rect 154642 346170 154698 346226
rect 154518 346046 154574 346102
rect 154642 346046 154698 346102
rect 154518 345922 154574 345978
rect 154642 345922 154698 345978
rect 159114 346294 159170 346350
rect 159238 346294 159294 346350
rect 159362 346294 159418 346350
rect 159486 346294 159542 346350
rect 159114 346170 159170 346226
rect 159238 346170 159294 346226
rect 159362 346170 159418 346226
rect 159486 346170 159542 346226
rect 159114 346046 159170 346102
rect 159238 346046 159294 346102
rect 159362 346046 159418 346102
rect 159486 346046 159542 346102
rect 159114 345922 159170 345978
rect 159238 345922 159294 345978
rect 159362 345922 159418 345978
rect 159486 345922 159542 345978
rect 154518 328294 154574 328350
rect 154642 328294 154698 328350
rect 154518 328170 154574 328226
rect 154642 328170 154698 328226
rect 154518 328046 154574 328102
rect 154642 328046 154698 328102
rect 154518 327922 154574 327978
rect 154642 327922 154698 327978
rect 159114 328294 159170 328350
rect 159238 328294 159294 328350
rect 159362 328294 159418 328350
rect 159486 328294 159542 328350
rect 159114 328170 159170 328226
rect 159238 328170 159294 328226
rect 159362 328170 159418 328226
rect 159486 328170 159542 328226
rect 159114 328046 159170 328102
rect 159238 328046 159294 328102
rect 159362 328046 159418 328102
rect 159486 328046 159542 328102
rect 159114 327922 159170 327978
rect 159238 327922 159294 327978
rect 159362 327922 159418 327978
rect 159486 327922 159542 327978
rect 159114 310294 159170 310350
rect 159238 310294 159294 310350
rect 159362 310294 159418 310350
rect 159486 310294 159542 310350
rect 159114 310170 159170 310226
rect 159238 310170 159294 310226
rect 159362 310170 159418 310226
rect 159486 310170 159542 310226
rect 159114 310046 159170 310102
rect 159238 310046 159294 310102
rect 159362 310046 159418 310102
rect 159486 310046 159542 310102
rect 159114 309922 159170 309978
rect 159238 309922 159294 309978
rect 159362 309922 159418 309978
rect 159486 309922 159542 309978
rect 159114 292294 159170 292350
rect 159238 292294 159294 292350
rect 159362 292294 159418 292350
rect 159486 292294 159542 292350
rect 159114 292170 159170 292226
rect 159238 292170 159294 292226
rect 159362 292170 159418 292226
rect 159486 292170 159542 292226
rect 159114 292046 159170 292102
rect 159238 292046 159294 292102
rect 159362 292046 159418 292102
rect 159486 292046 159542 292102
rect 159114 291922 159170 291978
rect 159238 291922 159294 291978
rect 159362 291922 159418 291978
rect 159486 291922 159542 291978
rect 132114 280294 132170 280350
rect 132238 280294 132294 280350
rect 132362 280294 132418 280350
rect 132486 280294 132542 280350
rect 132114 280170 132170 280226
rect 132238 280170 132294 280226
rect 132362 280170 132418 280226
rect 132486 280170 132542 280226
rect 132114 280046 132170 280102
rect 132238 280046 132294 280102
rect 132362 280046 132418 280102
rect 132486 280046 132542 280102
rect 132114 279922 132170 279978
rect 132238 279922 132294 279978
rect 132362 279922 132418 279978
rect 132486 279922 132542 279978
rect 132114 262294 132170 262350
rect 132238 262294 132294 262350
rect 132362 262294 132418 262350
rect 132486 262294 132542 262350
rect 132114 262170 132170 262226
rect 132238 262170 132294 262226
rect 132362 262170 132418 262226
rect 132486 262170 132542 262226
rect 132114 262046 132170 262102
rect 132238 262046 132294 262102
rect 132362 262046 132418 262102
rect 132486 262046 132542 262102
rect 132114 261922 132170 261978
rect 132238 261922 132294 261978
rect 132362 261922 132418 261978
rect 132486 261922 132542 261978
rect 132114 244294 132170 244350
rect 132238 244294 132294 244350
rect 132362 244294 132418 244350
rect 132486 244294 132542 244350
rect 132114 244170 132170 244226
rect 132238 244170 132294 244226
rect 132362 244170 132418 244226
rect 132486 244170 132542 244226
rect 132114 244046 132170 244102
rect 132238 244046 132294 244102
rect 132362 244046 132418 244102
rect 132486 244046 132542 244102
rect 132114 243922 132170 243978
rect 132238 243922 132294 243978
rect 132362 243922 132418 243978
rect 132486 243922 132542 243978
rect 132114 226294 132170 226350
rect 132238 226294 132294 226350
rect 132362 226294 132418 226350
rect 132486 226294 132542 226350
rect 132114 226170 132170 226226
rect 132238 226170 132294 226226
rect 132362 226170 132418 226226
rect 132486 226170 132542 226226
rect 132114 226046 132170 226102
rect 132238 226046 132294 226102
rect 132362 226046 132418 226102
rect 132486 226046 132542 226102
rect 132114 225922 132170 225978
rect 132238 225922 132294 225978
rect 132362 225922 132418 225978
rect 132486 225922 132542 225978
rect 162834 460294 162890 460350
rect 162958 460294 163014 460350
rect 163082 460294 163138 460350
rect 163206 460294 163262 460350
rect 162834 460170 162890 460226
rect 162958 460170 163014 460226
rect 163082 460170 163138 460226
rect 163206 460170 163262 460226
rect 162834 460046 162890 460102
rect 162958 460046 163014 460102
rect 163082 460046 163138 460102
rect 163206 460046 163262 460102
rect 162834 459922 162890 459978
rect 162958 459922 163014 459978
rect 163082 459922 163138 459978
rect 163206 459922 163262 459978
rect 162834 442294 162890 442350
rect 162958 442294 163014 442350
rect 163082 442294 163138 442350
rect 163206 442294 163262 442350
rect 162834 442170 162890 442226
rect 162958 442170 163014 442226
rect 163082 442170 163138 442226
rect 163206 442170 163262 442226
rect 162834 442046 162890 442102
rect 162958 442046 163014 442102
rect 163082 442046 163138 442102
rect 163206 442046 163262 442102
rect 162834 441922 162890 441978
rect 162958 441922 163014 441978
rect 163082 441922 163138 441978
rect 163206 441922 163262 441978
rect 162834 424294 162890 424350
rect 162958 424294 163014 424350
rect 163082 424294 163138 424350
rect 163206 424294 163262 424350
rect 162834 424170 162890 424226
rect 162958 424170 163014 424226
rect 163082 424170 163138 424226
rect 163206 424170 163262 424226
rect 162834 424046 162890 424102
rect 162958 424046 163014 424102
rect 163082 424046 163138 424102
rect 163206 424046 163262 424102
rect 162834 423922 162890 423978
rect 162958 423922 163014 423978
rect 163082 423922 163138 423978
rect 163206 423922 163262 423978
rect 162834 406294 162890 406350
rect 162958 406294 163014 406350
rect 163082 406294 163138 406350
rect 163206 406294 163262 406350
rect 162834 406170 162890 406226
rect 162958 406170 163014 406226
rect 163082 406170 163138 406226
rect 163206 406170 163262 406226
rect 162834 406046 162890 406102
rect 162958 406046 163014 406102
rect 163082 406046 163138 406102
rect 163206 406046 163262 406102
rect 162834 405922 162890 405978
rect 162958 405922 163014 405978
rect 163082 405922 163138 405978
rect 163206 405922 163262 405978
rect 162834 388294 162890 388350
rect 162958 388294 163014 388350
rect 163082 388294 163138 388350
rect 163206 388294 163262 388350
rect 162834 388170 162890 388226
rect 162958 388170 163014 388226
rect 163082 388170 163138 388226
rect 163206 388170 163262 388226
rect 162834 388046 162890 388102
rect 162958 388046 163014 388102
rect 163082 388046 163138 388102
rect 163206 388046 163262 388102
rect 162834 387922 162890 387978
rect 162958 387922 163014 387978
rect 163082 387922 163138 387978
rect 163206 387922 163262 387978
rect 162834 370294 162890 370350
rect 162958 370294 163014 370350
rect 163082 370294 163138 370350
rect 163206 370294 163262 370350
rect 162834 370170 162890 370226
rect 162958 370170 163014 370226
rect 163082 370170 163138 370226
rect 163206 370170 163262 370226
rect 162834 370046 162890 370102
rect 162958 370046 163014 370102
rect 163082 370046 163138 370102
rect 163206 370046 163262 370102
rect 162834 369922 162890 369978
rect 162958 369922 163014 369978
rect 163082 369922 163138 369978
rect 163206 369922 163262 369978
rect 162834 352294 162890 352350
rect 162958 352294 163014 352350
rect 163082 352294 163138 352350
rect 163206 352294 163262 352350
rect 162834 352170 162890 352226
rect 162958 352170 163014 352226
rect 163082 352170 163138 352226
rect 163206 352170 163262 352226
rect 162834 352046 162890 352102
rect 162958 352046 163014 352102
rect 163082 352046 163138 352102
rect 163206 352046 163262 352102
rect 162834 351922 162890 351978
rect 162958 351922 163014 351978
rect 163082 351922 163138 351978
rect 163206 351922 163262 351978
rect 162834 334294 162890 334350
rect 162958 334294 163014 334350
rect 163082 334294 163138 334350
rect 163206 334294 163262 334350
rect 162834 334170 162890 334226
rect 162958 334170 163014 334226
rect 163082 334170 163138 334226
rect 163206 334170 163262 334226
rect 162834 334046 162890 334102
rect 162958 334046 163014 334102
rect 163082 334046 163138 334102
rect 163206 334046 163262 334102
rect 162834 333922 162890 333978
rect 162958 333922 163014 333978
rect 163082 333922 163138 333978
rect 163206 333922 163262 333978
rect 162834 316294 162890 316350
rect 162958 316294 163014 316350
rect 163082 316294 163138 316350
rect 163206 316294 163262 316350
rect 162834 316170 162890 316226
rect 162958 316170 163014 316226
rect 163082 316170 163138 316226
rect 163206 316170 163262 316226
rect 162834 316046 162890 316102
rect 162958 316046 163014 316102
rect 163082 316046 163138 316102
rect 163206 316046 163262 316102
rect 162834 315922 162890 315978
rect 162958 315922 163014 315978
rect 163082 315922 163138 315978
rect 163206 315922 163262 315978
rect 162834 298294 162890 298350
rect 162958 298294 163014 298350
rect 163082 298294 163138 298350
rect 163206 298294 163262 298350
rect 162834 298170 162890 298226
rect 162958 298170 163014 298226
rect 163082 298170 163138 298226
rect 163206 298170 163262 298226
rect 162834 298046 162890 298102
rect 162958 298046 163014 298102
rect 163082 298046 163138 298102
rect 163206 298046 163262 298102
rect 162834 297922 162890 297978
rect 162958 297922 163014 297978
rect 163082 297922 163138 297978
rect 163206 297922 163262 297978
rect 159114 274294 159170 274350
rect 159238 274294 159294 274350
rect 159362 274294 159418 274350
rect 159486 274294 159542 274350
rect 159114 274170 159170 274226
rect 159238 274170 159294 274226
rect 159362 274170 159418 274226
rect 159486 274170 159542 274226
rect 159114 274046 159170 274102
rect 159238 274046 159294 274102
rect 159362 274046 159418 274102
rect 159486 274046 159542 274102
rect 159114 273922 159170 273978
rect 159238 273922 159294 273978
rect 159362 273922 159418 273978
rect 159486 273922 159542 273978
rect 159114 256294 159170 256350
rect 159238 256294 159294 256350
rect 159362 256294 159418 256350
rect 159486 256294 159542 256350
rect 159114 256170 159170 256226
rect 159238 256170 159294 256226
rect 159362 256170 159418 256226
rect 159486 256170 159542 256226
rect 159114 256046 159170 256102
rect 159238 256046 159294 256102
rect 159362 256046 159418 256102
rect 159486 256046 159542 256102
rect 159114 255922 159170 255978
rect 159238 255922 159294 255978
rect 159362 255922 159418 255978
rect 159486 255922 159542 255978
rect 159114 238294 159170 238350
rect 159238 238294 159294 238350
rect 159362 238294 159418 238350
rect 159486 238294 159542 238350
rect 159114 238170 159170 238226
rect 159238 238170 159294 238226
rect 159362 238170 159418 238226
rect 159486 238170 159542 238226
rect 159114 238046 159170 238102
rect 159238 238046 159294 238102
rect 159362 238046 159418 238102
rect 159486 238046 159542 238102
rect 159114 237922 159170 237978
rect 159238 237922 159294 237978
rect 159362 237922 159418 237978
rect 159486 237922 159542 237978
rect 159114 220294 159170 220350
rect 159238 220294 159294 220350
rect 159362 220294 159418 220350
rect 159486 220294 159542 220350
rect 159114 220170 159170 220226
rect 159238 220170 159294 220226
rect 159362 220170 159418 220226
rect 159486 220170 159542 220226
rect 159114 220046 159170 220102
rect 159238 220046 159294 220102
rect 159362 220046 159418 220102
rect 159486 220046 159542 220102
rect 159114 219922 159170 219978
rect 159238 219922 159294 219978
rect 159362 219922 159418 219978
rect 159486 219922 159542 219978
rect 189834 562294 189890 562350
rect 189958 562294 190014 562350
rect 190082 562294 190138 562350
rect 190206 562294 190262 562350
rect 189834 562170 189890 562226
rect 189958 562170 190014 562226
rect 190082 562170 190138 562226
rect 190206 562170 190262 562226
rect 189834 562046 189890 562102
rect 189958 562046 190014 562102
rect 190082 562046 190138 562102
rect 190206 562046 190262 562102
rect 189834 561922 189890 561978
rect 189958 561922 190014 561978
rect 190082 561922 190138 561978
rect 190206 561922 190262 561978
rect 169878 352294 169934 352350
rect 170002 352294 170058 352350
rect 169878 352170 169934 352226
rect 170002 352170 170058 352226
rect 169878 352046 169934 352102
rect 170002 352046 170058 352102
rect 169878 351922 169934 351978
rect 170002 351922 170058 351978
rect 185238 346294 185294 346350
rect 185362 346294 185418 346350
rect 185238 346170 185294 346226
rect 185362 346170 185418 346226
rect 185238 346046 185294 346102
rect 185362 346046 185418 346102
rect 185238 345922 185294 345978
rect 185362 345922 185418 345978
rect 169878 334294 169934 334350
rect 170002 334294 170058 334350
rect 169878 334170 169934 334226
rect 170002 334170 170058 334226
rect 169878 334046 169934 334102
rect 170002 334046 170058 334102
rect 169878 333922 169934 333978
rect 170002 333922 170058 333978
rect 185238 328294 185294 328350
rect 185362 328294 185418 328350
rect 185238 328170 185294 328226
rect 185362 328170 185418 328226
rect 185238 328046 185294 328102
rect 185362 328046 185418 328102
rect 185238 327922 185294 327978
rect 185362 327922 185418 327978
rect 162834 280294 162890 280350
rect 162958 280294 163014 280350
rect 163082 280294 163138 280350
rect 163206 280294 163262 280350
rect 162834 280170 162890 280226
rect 162958 280170 163014 280226
rect 163082 280170 163138 280226
rect 163206 280170 163262 280226
rect 162834 280046 162890 280102
rect 162958 280046 163014 280102
rect 163082 280046 163138 280102
rect 163206 280046 163262 280102
rect 162834 279922 162890 279978
rect 162958 279922 163014 279978
rect 163082 279922 163138 279978
rect 163206 279922 163262 279978
rect 167078 280294 167134 280350
rect 167202 280294 167258 280350
rect 167078 280170 167134 280226
rect 167202 280170 167258 280226
rect 167078 280046 167134 280102
rect 167202 280046 167258 280102
rect 167078 279922 167134 279978
rect 167202 279922 167258 279978
rect 172902 280294 172958 280350
rect 173026 280294 173082 280350
rect 172902 280170 172958 280226
rect 173026 280170 173082 280226
rect 172902 280046 172958 280102
rect 173026 280046 173082 280102
rect 172902 279922 172958 279978
rect 173026 279922 173082 279978
rect 178726 280294 178782 280350
rect 178850 280294 178906 280350
rect 178726 280170 178782 280226
rect 178850 280170 178906 280226
rect 178726 280046 178782 280102
rect 178850 280046 178906 280102
rect 178726 279922 178782 279978
rect 178850 279922 178906 279978
rect 184550 280294 184606 280350
rect 184674 280294 184730 280350
rect 184550 280170 184606 280226
rect 184674 280170 184730 280226
rect 184550 280046 184606 280102
rect 184674 280046 184730 280102
rect 184550 279922 184606 279978
rect 184674 279922 184730 279978
rect 164166 274294 164222 274350
rect 164290 274294 164346 274350
rect 164166 274170 164222 274226
rect 164290 274170 164346 274226
rect 164166 274046 164222 274102
rect 164290 274046 164346 274102
rect 164166 273922 164222 273978
rect 164290 273922 164346 273978
rect 169990 274294 170046 274350
rect 170114 274294 170170 274350
rect 169990 274170 170046 274226
rect 170114 274170 170170 274226
rect 169990 274046 170046 274102
rect 170114 274046 170170 274102
rect 169990 273922 170046 273978
rect 170114 273922 170170 273978
rect 175814 274294 175870 274350
rect 175938 274294 175994 274350
rect 175814 274170 175870 274226
rect 175938 274170 175994 274226
rect 175814 274046 175870 274102
rect 175938 274046 175994 274102
rect 175814 273922 175870 273978
rect 175938 273922 175994 273978
rect 181638 274294 181694 274350
rect 181762 274294 181818 274350
rect 181638 274170 181694 274226
rect 181762 274170 181818 274226
rect 181638 274046 181694 274102
rect 181762 274046 181818 274102
rect 181638 273922 181694 273978
rect 181762 273922 181818 273978
rect 189834 544294 189890 544350
rect 189958 544294 190014 544350
rect 190082 544294 190138 544350
rect 190206 544294 190262 544350
rect 189834 544170 189890 544226
rect 189958 544170 190014 544226
rect 190082 544170 190138 544226
rect 190206 544170 190262 544226
rect 189834 544046 189890 544102
rect 189958 544046 190014 544102
rect 190082 544046 190138 544102
rect 190206 544046 190262 544102
rect 189834 543922 189890 543978
rect 189958 543922 190014 543978
rect 190082 543922 190138 543978
rect 190206 543922 190262 543978
rect 189834 526294 189890 526350
rect 189958 526294 190014 526350
rect 190082 526294 190138 526350
rect 190206 526294 190262 526350
rect 189834 526170 189890 526226
rect 189958 526170 190014 526226
rect 190082 526170 190138 526226
rect 190206 526170 190262 526226
rect 189834 526046 189890 526102
rect 189958 526046 190014 526102
rect 190082 526046 190138 526102
rect 190206 526046 190262 526102
rect 189834 525922 189890 525978
rect 189958 525922 190014 525978
rect 190082 525922 190138 525978
rect 190206 525922 190262 525978
rect 189834 508294 189890 508350
rect 189958 508294 190014 508350
rect 190082 508294 190138 508350
rect 190206 508294 190262 508350
rect 189834 508170 189890 508226
rect 189958 508170 190014 508226
rect 190082 508170 190138 508226
rect 190206 508170 190262 508226
rect 189834 508046 189890 508102
rect 189958 508046 190014 508102
rect 190082 508046 190138 508102
rect 190206 508046 190262 508102
rect 189834 507922 189890 507978
rect 189958 507922 190014 507978
rect 190082 507922 190138 507978
rect 190206 507922 190262 507978
rect 162834 262294 162890 262350
rect 162958 262294 163014 262350
rect 163082 262294 163138 262350
rect 163206 262294 163262 262350
rect 162834 262170 162890 262226
rect 162958 262170 163014 262226
rect 163082 262170 163138 262226
rect 163206 262170 163262 262226
rect 162834 262046 162890 262102
rect 162958 262046 163014 262102
rect 163082 262046 163138 262102
rect 163206 262046 163262 262102
rect 162834 261922 162890 261978
rect 162958 261922 163014 261978
rect 163082 261922 163138 261978
rect 163206 261922 163262 261978
rect 189834 490294 189890 490350
rect 189958 490294 190014 490350
rect 190082 490294 190138 490350
rect 190206 490294 190262 490350
rect 189834 490170 189890 490226
rect 189958 490170 190014 490226
rect 190082 490170 190138 490226
rect 190206 490170 190262 490226
rect 189834 490046 189890 490102
rect 189958 490046 190014 490102
rect 190082 490046 190138 490102
rect 190206 490046 190262 490102
rect 189834 489922 189890 489978
rect 189958 489922 190014 489978
rect 190082 489922 190138 489978
rect 190206 489922 190262 489978
rect 189834 472294 189890 472350
rect 189958 472294 190014 472350
rect 190082 472294 190138 472350
rect 190206 472294 190262 472350
rect 189834 472170 189890 472226
rect 189958 472170 190014 472226
rect 190082 472170 190138 472226
rect 190206 472170 190262 472226
rect 189834 472046 189890 472102
rect 189958 472046 190014 472102
rect 190082 472046 190138 472102
rect 190206 472046 190262 472102
rect 189834 471922 189890 471978
rect 189958 471922 190014 471978
rect 190082 471922 190138 471978
rect 190206 471922 190262 471978
rect 189834 454294 189890 454350
rect 189958 454294 190014 454350
rect 190082 454294 190138 454350
rect 190206 454294 190262 454350
rect 189834 454170 189890 454226
rect 189958 454170 190014 454226
rect 190082 454170 190138 454226
rect 190206 454170 190262 454226
rect 189834 454046 189890 454102
rect 189958 454046 190014 454102
rect 190082 454046 190138 454102
rect 190206 454046 190262 454102
rect 189834 453922 189890 453978
rect 189958 453922 190014 453978
rect 190082 453922 190138 453978
rect 190206 453922 190262 453978
rect 189834 436294 189890 436350
rect 189958 436294 190014 436350
rect 190082 436294 190138 436350
rect 190206 436294 190262 436350
rect 189834 436170 189890 436226
rect 189958 436170 190014 436226
rect 190082 436170 190138 436226
rect 190206 436170 190262 436226
rect 189834 436046 189890 436102
rect 189958 436046 190014 436102
rect 190082 436046 190138 436102
rect 190206 436046 190262 436102
rect 189834 435922 189890 435978
rect 189958 435922 190014 435978
rect 190082 435922 190138 435978
rect 190206 435922 190262 435978
rect 189834 418294 189890 418350
rect 189958 418294 190014 418350
rect 190082 418294 190138 418350
rect 190206 418294 190262 418350
rect 189834 418170 189890 418226
rect 189958 418170 190014 418226
rect 190082 418170 190138 418226
rect 190206 418170 190262 418226
rect 189834 418046 189890 418102
rect 189958 418046 190014 418102
rect 190082 418046 190138 418102
rect 190206 418046 190262 418102
rect 189834 417922 189890 417978
rect 189958 417922 190014 417978
rect 190082 417922 190138 417978
rect 190206 417922 190262 417978
rect 190652 589922 190708 589978
rect 189834 400294 189890 400350
rect 189958 400294 190014 400350
rect 190082 400294 190138 400350
rect 190206 400294 190262 400350
rect 189834 400170 189890 400226
rect 189958 400170 190014 400226
rect 190082 400170 190138 400226
rect 190206 400170 190262 400226
rect 189834 400046 189890 400102
rect 189958 400046 190014 400102
rect 190082 400046 190138 400102
rect 190206 400046 190262 400102
rect 189834 399922 189890 399978
rect 189958 399922 190014 399978
rect 190082 399922 190138 399978
rect 190206 399922 190262 399978
rect 189834 382294 189890 382350
rect 189958 382294 190014 382350
rect 190082 382294 190138 382350
rect 190206 382294 190262 382350
rect 189834 382170 189890 382226
rect 189958 382170 190014 382226
rect 190082 382170 190138 382226
rect 190206 382170 190262 382226
rect 189834 382046 189890 382102
rect 189958 382046 190014 382102
rect 190082 382046 190138 382102
rect 190206 382046 190262 382102
rect 189834 381922 189890 381978
rect 189958 381922 190014 381978
rect 190082 381922 190138 381978
rect 190206 381922 190262 381978
rect 189834 364294 189890 364350
rect 189958 364294 190014 364350
rect 190082 364294 190138 364350
rect 190206 364294 190262 364350
rect 189834 364170 189890 364226
rect 189958 364170 190014 364226
rect 190082 364170 190138 364226
rect 190206 364170 190262 364226
rect 189834 364046 189890 364102
rect 189958 364046 190014 364102
rect 190082 364046 190138 364102
rect 190206 364046 190262 364102
rect 189834 363922 189890 363978
rect 189958 363922 190014 363978
rect 190082 363922 190138 363978
rect 190206 363922 190262 363978
rect 189834 346294 189890 346350
rect 189958 346294 190014 346350
rect 190082 346294 190138 346350
rect 190206 346294 190262 346350
rect 189834 346170 189890 346226
rect 189958 346170 190014 346226
rect 190082 346170 190138 346226
rect 190206 346170 190262 346226
rect 189834 346046 189890 346102
rect 189958 346046 190014 346102
rect 190082 346046 190138 346102
rect 190206 346046 190262 346102
rect 189834 345922 189890 345978
rect 189958 345922 190014 345978
rect 190082 345922 190138 345978
rect 190206 345922 190262 345978
rect 189834 328294 189890 328350
rect 189958 328294 190014 328350
rect 190082 328294 190138 328350
rect 190206 328294 190262 328350
rect 189834 328170 189890 328226
rect 189958 328170 190014 328226
rect 190082 328170 190138 328226
rect 190206 328170 190262 328226
rect 189834 328046 189890 328102
rect 189958 328046 190014 328102
rect 190082 328046 190138 328102
rect 190206 328046 190262 328102
rect 189834 327922 189890 327978
rect 189958 327922 190014 327978
rect 190082 327922 190138 327978
rect 190206 327922 190262 327978
rect 189834 310294 189890 310350
rect 189958 310294 190014 310350
rect 190082 310294 190138 310350
rect 190206 310294 190262 310350
rect 189834 310170 189890 310226
rect 189958 310170 190014 310226
rect 190082 310170 190138 310226
rect 190206 310170 190262 310226
rect 189834 310046 189890 310102
rect 189958 310046 190014 310102
rect 190082 310046 190138 310102
rect 190206 310046 190262 310102
rect 189834 309922 189890 309978
rect 189958 309922 190014 309978
rect 190082 309922 190138 309978
rect 190206 309922 190262 309978
rect 189834 292294 189890 292350
rect 189958 292294 190014 292350
rect 190082 292294 190138 292350
rect 190206 292294 190262 292350
rect 189834 292170 189890 292226
rect 189958 292170 190014 292226
rect 190082 292170 190138 292226
rect 190206 292170 190262 292226
rect 189834 292046 189890 292102
rect 189958 292046 190014 292102
rect 190082 292046 190138 292102
rect 190206 292046 190262 292102
rect 189834 291922 189890 291978
rect 189958 291922 190014 291978
rect 190082 291922 190138 291978
rect 190206 291922 190262 291978
rect 193116 589742 193172 589798
rect 193554 586294 193610 586350
rect 193678 586294 193734 586350
rect 193802 586294 193858 586350
rect 193926 586294 193982 586350
rect 193554 586170 193610 586226
rect 193678 586170 193734 586226
rect 193802 586170 193858 586226
rect 193926 586170 193982 586226
rect 193554 586046 193610 586102
rect 193678 586046 193734 586102
rect 193802 586046 193858 586102
rect 193926 586046 193982 586102
rect 193554 585922 193610 585978
rect 193678 585922 193734 585978
rect 193802 585922 193858 585978
rect 193926 585922 193982 585978
rect 220554 597156 220610 597212
rect 220678 597156 220734 597212
rect 220802 597156 220858 597212
rect 220926 597156 220982 597212
rect 220554 597032 220610 597088
rect 220678 597032 220734 597088
rect 220802 597032 220858 597088
rect 220926 597032 220982 597088
rect 220554 596908 220610 596964
rect 220678 596908 220734 596964
rect 220802 596908 220858 596964
rect 220926 596908 220982 596964
rect 220554 596784 220610 596840
rect 220678 596784 220734 596840
rect 220802 596784 220858 596840
rect 220926 596784 220982 596840
rect 220554 580294 220610 580350
rect 220678 580294 220734 580350
rect 220802 580294 220858 580350
rect 220926 580294 220982 580350
rect 220554 580170 220610 580226
rect 220678 580170 220734 580226
rect 220802 580170 220858 580226
rect 220926 580170 220982 580226
rect 220554 580046 220610 580102
rect 220678 580046 220734 580102
rect 220802 580046 220858 580102
rect 220926 580046 220982 580102
rect 220554 579922 220610 579978
rect 220678 579922 220734 579978
rect 220802 579922 220858 579978
rect 220926 579922 220982 579978
rect 224274 598116 224330 598172
rect 224398 598116 224454 598172
rect 224522 598116 224578 598172
rect 224646 598116 224702 598172
rect 224274 597992 224330 598048
rect 224398 597992 224454 598048
rect 224522 597992 224578 598048
rect 224646 597992 224702 598048
rect 224274 597868 224330 597924
rect 224398 597868 224454 597924
rect 224522 597868 224578 597924
rect 224646 597868 224702 597924
rect 224274 597744 224330 597800
rect 224398 597744 224454 597800
rect 224522 597744 224578 597800
rect 224646 597744 224702 597800
rect 224274 586294 224330 586350
rect 224398 586294 224454 586350
rect 224522 586294 224578 586350
rect 224646 586294 224702 586350
rect 224274 586170 224330 586226
rect 224398 586170 224454 586226
rect 224522 586170 224578 586226
rect 224646 586170 224702 586226
rect 224274 586046 224330 586102
rect 224398 586046 224454 586102
rect 224522 586046 224578 586102
rect 224646 586046 224702 586102
rect 224274 585922 224330 585978
rect 224398 585922 224454 585978
rect 224522 585922 224578 585978
rect 224646 585922 224702 585978
rect 251274 597156 251330 597212
rect 251398 597156 251454 597212
rect 251522 597156 251578 597212
rect 251646 597156 251702 597212
rect 251274 597032 251330 597088
rect 251398 597032 251454 597088
rect 251522 597032 251578 597088
rect 251646 597032 251702 597088
rect 251274 596908 251330 596964
rect 251398 596908 251454 596964
rect 251522 596908 251578 596964
rect 251646 596908 251702 596964
rect 251274 596784 251330 596840
rect 251398 596784 251454 596840
rect 251522 596784 251578 596840
rect 251646 596784 251702 596840
rect 251274 580294 251330 580350
rect 251398 580294 251454 580350
rect 251522 580294 251578 580350
rect 251646 580294 251702 580350
rect 251274 580170 251330 580226
rect 251398 580170 251454 580226
rect 251522 580170 251578 580226
rect 251646 580170 251702 580226
rect 251274 580046 251330 580102
rect 251398 580046 251454 580102
rect 251522 580046 251578 580102
rect 251646 580046 251702 580102
rect 251274 579922 251330 579978
rect 251398 579922 251454 579978
rect 251522 579922 251578 579978
rect 251646 579922 251702 579978
rect 254994 598116 255050 598172
rect 255118 598116 255174 598172
rect 255242 598116 255298 598172
rect 255366 598116 255422 598172
rect 254994 597992 255050 598048
rect 255118 597992 255174 598048
rect 255242 597992 255298 598048
rect 255366 597992 255422 598048
rect 254994 597868 255050 597924
rect 255118 597868 255174 597924
rect 255242 597868 255298 597924
rect 255366 597868 255422 597924
rect 254994 597744 255050 597800
rect 255118 597744 255174 597800
rect 255242 597744 255298 597800
rect 255366 597744 255422 597800
rect 254994 586294 255050 586350
rect 255118 586294 255174 586350
rect 255242 586294 255298 586350
rect 255366 586294 255422 586350
rect 254994 586170 255050 586226
rect 255118 586170 255174 586226
rect 255242 586170 255298 586226
rect 255366 586170 255422 586226
rect 254994 586046 255050 586102
rect 255118 586046 255174 586102
rect 255242 586046 255298 586102
rect 255366 586046 255422 586102
rect 254994 585922 255050 585978
rect 255118 585922 255174 585978
rect 255242 585922 255298 585978
rect 255366 585922 255422 585978
rect 281994 597156 282050 597212
rect 282118 597156 282174 597212
rect 282242 597156 282298 597212
rect 282366 597156 282422 597212
rect 281994 597032 282050 597088
rect 282118 597032 282174 597088
rect 282242 597032 282298 597088
rect 282366 597032 282422 597088
rect 281994 596908 282050 596964
rect 282118 596908 282174 596964
rect 282242 596908 282298 596964
rect 282366 596908 282422 596964
rect 281994 596784 282050 596840
rect 282118 596784 282174 596840
rect 282242 596784 282298 596840
rect 282366 596784 282422 596840
rect 281994 580294 282050 580350
rect 282118 580294 282174 580350
rect 282242 580294 282298 580350
rect 282366 580294 282422 580350
rect 281994 580170 282050 580226
rect 282118 580170 282174 580226
rect 282242 580170 282298 580226
rect 282366 580170 282422 580226
rect 281994 580046 282050 580102
rect 282118 580046 282174 580102
rect 282242 580046 282298 580102
rect 282366 580046 282422 580102
rect 281994 579922 282050 579978
rect 282118 579922 282174 579978
rect 282242 579922 282298 579978
rect 282366 579922 282422 579978
rect 285714 598116 285770 598172
rect 285838 598116 285894 598172
rect 285962 598116 286018 598172
rect 286086 598116 286142 598172
rect 285714 597992 285770 598048
rect 285838 597992 285894 598048
rect 285962 597992 286018 598048
rect 286086 597992 286142 598048
rect 285714 597868 285770 597924
rect 285838 597868 285894 597924
rect 285962 597868 286018 597924
rect 286086 597868 286142 597924
rect 285714 597744 285770 597800
rect 285838 597744 285894 597800
rect 285962 597744 286018 597800
rect 286086 597744 286142 597800
rect 285714 586294 285770 586350
rect 285838 586294 285894 586350
rect 285962 586294 286018 586350
rect 286086 586294 286142 586350
rect 285714 586170 285770 586226
rect 285838 586170 285894 586226
rect 285962 586170 286018 586226
rect 286086 586170 286142 586226
rect 285714 586046 285770 586102
rect 285838 586046 285894 586102
rect 285962 586046 286018 586102
rect 286086 586046 286142 586102
rect 285714 585922 285770 585978
rect 285838 585922 285894 585978
rect 285962 585922 286018 585978
rect 286086 585922 286142 585978
rect 312714 597156 312770 597212
rect 312838 597156 312894 597212
rect 312962 597156 313018 597212
rect 313086 597156 313142 597212
rect 312714 597032 312770 597088
rect 312838 597032 312894 597088
rect 312962 597032 313018 597088
rect 313086 597032 313142 597088
rect 312714 596908 312770 596964
rect 312838 596908 312894 596964
rect 312962 596908 313018 596964
rect 313086 596908 313142 596964
rect 312714 596784 312770 596840
rect 312838 596784 312894 596840
rect 312962 596784 313018 596840
rect 313086 596784 313142 596840
rect 312714 580294 312770 580350
rect 312838 580294 312894 580350
rect 312962 580294 313018 580350
rect 313086 580294 313142 580350
rect 312714 580170 312770 580226
rect 312838 580170 312894 580226
rect 312962 580170 313018 580226
rect 313086 580170 313142 580226
rect 312714 580046 312770 580102
rect 312838 580046 312894 580102
rect 312962 580046 313018 580102
rect 313086 580046 313142 580102
rect 312714 579922 312770 579978
rect 312838 579922 312894 579978
rect 312962 579922 313018 579978
rect 313086 579922 313142 579978
rect 316434 598116 316490 598172
rect 316558 598116 316614 598172
rect 316682 598116 316738 598172
rect 316806 598116 316862 598172
rect 316434 597992 316490 598048
rect 316558 597992 316614 598048
rect 316682 597992 316738 598048
rect 316806 597992 316862 598048
rect 316434 597868 316490 597924
rect 316558 597868 316614 597924
rect 316682 597868 316738 597924
rect 316806 597868 316862 597924
rect 316434 597744 316490 597800
rect 316558 597744 316614 597800
rect 316682 597744 316738 597800
rect 316806 597744 316862 597800
rect 316434 586294 316490 586350
rect 316558 586294 316614 586350
rect 316682 586294 316738 586350
rect 316806 586294 316862 586350
rect 316434 586170 316490 586226
rect 316558 586170 316614 586226
rect 316682 586170 316738 586226
rect 316806 586170 316862 586226
rect 316434 586046 316490 586102
rect 316558 586046 316614 586102
rect 316682 586046 316738 586102
rect 316806 586046 316862 586102
rect 316434 585922 316490 585978
rect 316558 585922 316614 585978
rect 316682 585922 316738 585978
rect 316806 585922 316862 585978
rect 343434 597156 343490 597212
rect 343558 597156 343614 597212
rect 343682 597156 343738 597212
rect 343806 597156 343862 597212
rect 343434 597032 343490 597088
rect 343558 597032 343614 597088
rect 343682 597032 343738 597088
rect 343806 597032 343862 597088
rect 343434 596908 343490 596964
rect 343558 596908 343614 596964
rect 343682 596908 343738 596964
rect 343806 596908 343862 596964
rect 343434 596784 343490 596840
rect 343558 596784 343614 596840
rect 343682 596784 343738 596840
rect 343806 596784 343862 596840
rect 343434 580294 343490 580350
rect 343558 580294 343614 580350
rect 343682 580294 343738 580350
rect 343806 580294 343862 580350
rect 343434 580170 343490 580226
rect 343558 580170 343614 580226
rect 343682 580170 343738 580226
rect 343806 580170 343862 580226
rect 343434 580046 343490 580102
rect 343558 580046 343614 580102
rect 343682 580046 343738 580102
rect 343806 580046 343862 580102
rect 343434 579922 343490 579978
rect 343558 579922 343614 579978
rect 343682 579922 343738 579978
rect 343806 579922 343862 579978
rect 347154 598116 347210 598172
rect 347278 598116 347334 598172
rect 347402 598116 347458 598172
rect 347526 598116 347582 598172
rect 347154 597992 347210 598048
rect 347278 597992 347334 598048
rect 347402 597992 347458 598048
rect 347526 597992 347582 598048
rect 347154 597868 347210 597924
rect 347278 597868 347334 597924
rect 347402 597868 347458 597924
rect 347526 597868 347582 597924
rect 347154 597744 347210 597800
rect 347278 597744 347334 597800
rect 347402 597744 347458 597800
rect 347526 597744 347582 597800
rect 347154 586294 347210 586350
rect 347278 586294 347334 586350
rect 347402 586294 347458 586350
rect 347526 586294 347582 586350
rect 347154 586170 347210 586226
rect 347278 586170 347334 586226
rect 347402 586170 347458 586226
rect 347526 586170 347582 586226
rect 347154 586046 347210 586102
rect 347278 586046 347334 586102
rect 347402 586046 347458 586102
rect 347526 586046 347582 586102
rect 347154 585922 347210 585978
rect 347278 585922 347334 585978
rect 347402 585922 347458 585978
rect 347526 585922 347582 585978
rect 374154 597156 374210 597212
rect 374278 597156 374334 597212
rect 374402 597156 374458 597212
rect 374526 597156 374582 597212
rect 374154 597032 374210 597088
rect 374278 597032 374334 597088
rect 374402 597032 374458 597088
rect 374526 597032 374582 597088
rect 374154 596908 374210 596964
rect 374278 596908 374334 596964
rect 374402 596908 374458 596964
rect 374526 596908 374582 596964
rect 374154 596784 374210 596840
rect 374278 596784 374334 596840
rect 374402 596784 374458 596840
rect 374526 596784 374582 596840
rect 374154 580294 374210 580350
rect 374278 580294 374334 580350
rect 374402 580294 374458 580350
rect 374526 580294 374582 580350
rect 374154 580170 374210 580226
rect 374278 580170 374334 580226
rect 374402 580170 374458 580226
rect 374526 580170 374582 580226
rect 374154 580046 374210 580102
rect 374278 580046 374334 580102
rect 374402 580046 374458 580102
rect 374526 580046 374582 580102
rect 374154 579922 374210 579978
rect 374278 579922 374334 579978
rect 374402 579922 374458 579978
rect 374526 579922 374582 579978
rect 377874 598116 377930 598172
rect 377998 598116 378054 598172
rect 378122 598116 378178 598172
rect 378246 598116 378302 598172
rect 377874 597992 377930 598048
rect 377998 597992 378054 598048
rect 378122 597992 378178 598048
rect 378246 597992 378302 598048
rect 377874 597868 377930 597924
rect 377998 597868 378054 597924
rect 378122 597868 378178 597924
rect 378246 597868 378302 597924
rect 377874 597744 377930 597800
rect 377998 597744 378054 597800
rect 378122 597744 378178 597800
rect 378246 597744 378302 597800
rect 377874 586294 377930 586350
rect 377998 586294 378054 586350
rect 378122 586294 378178 586350
rect 378246 586294 378302 586350
rect 377874 586170 377930 586226
rect 377998 586170 378054 586226
rect 378122 586170 378178 586226
rect 378246 586170 378302 586226
rect 377874 586046 377930 586102
rect 377998 586046 378054 586102
rect 378122 586046 378178 586102
rect 378246 586046 378302 586102
rect 377874 585922 377930 585978
rect 377998 585922 378054 585978
rect 378122 585922 378178 585978
rect 378246 585922 378302 585978
rect 404874 597156 404930 597212
rect 404998 597156 405054 597212
rect 405122 597156 405178 597212
rect 405246 597156 405302 597212
rect 404874 597032 404930 597088
rect 404998 597032 405054 597088
rect 405122 597032 405178 597088
rect 405246 597032 405302 597088
rect 404874 596908 404930 596964
rect 404998 596908 405054 596964
rect 405122 596908 405178 596964
rect 405246 596908 405302 596964
rect 404874 596784 404930 596840
rect 404998 596784 405054 596840
rect 405122 596784 405178 596840
rect 405246 596784 405302 596840
rect 408594 598116 408650 598172
rect 408718 598116 408774 598172
rect 408842 598116 408898 598172
rect 408966 598116 409022 598172
rect 408594 597992 408650 598048
rect 408718 597992 408774 598048
rect 408842 597992 408898 598048
rect 408966 597992 409022 598048
rect 408594 597868 408650 597924
rect 408718 597868 408774 597924
rect 408842 597868 408898 597924
rect 408966 597868 409022 597924
rect 408594 597744 408650 597800
rect 408718 597744 408774 597800
rect 408842 597744 408898 597800
rect 408966 597744 409022 597800
rect 408268 589922 408324 589978
rect 404874 580294 404930 580350
rect 404998 580294 405054 580350
rect 405122 580294 405178 580350
rect 405246 580294 405302 580350
rect 404874 580170 404930 580226
rect 404998 580170 405054 580226
rect 405122 580170 405178 580226
rect 405246 580170 405302 580226
rect 404874 580046 404930 580102
rect 404998 580046 405054 580102
rect 405122 580046 405178 580102
rect 405246 580046 405302 580102
rect 404874 579922 404930 579978
rect 404998 579922 405054 579978
rect 405122 579922 405178 579978
rect 405246 579922 405302 579978
rect 408594 586294 408650 586350
rect 408718 586294 408774 586350
rect 408842 586294 408898 586350
rect 408966 586294 409022 586350
rect 408594 586170 408650 586226
rect 408718 586170 408774 586226
rect 408842 586170 408898 586226
rect 408966 586170 409022 586226
rect 408594 586046 408650 586102
rect 408718 586046 408774 586102
rect 408842 586046 408898 586102
rect 408966 586046 409022 586102
rect 408594 585922 408650 585978
rect 408718 585922 408774 585978
rect 408842 585922 408898 585978
rect 408966 585922 409022 585978
rect 435594 597156 435650 597212
rect 435718 597156 435774 597212
rect 435842 597156 435898 597212
rect 435966 597156 436022 597212
rect 435594 597032 435650 597088
rect 435718 597032 435774 597088
rect 435842 597032 435898 597088
rect 435966 597032 436022 597088
rect 435594 596908 435650 596964
rect 435718 596908 435774 596964
rect 435842 596908 435898 596964
rect 435966 596908 436022 596964
rect 435594 596784 435650 596840
rect 435718 596784 435774 596840
rect 435842 596784 435898 596840
rect 435966 596784 436022 596840
rect 435594 580294 435650 580350
rect 435718 580294 435774 580350
rect 435842 580294 435898 580350
rect 435966 580294 436022 580350
rect 435594 580170 435650 580226
rect 435718 580170 435774 580226
rect 435842 580170 435898 580226
rect 435966 580170 436022 580226
rect 435594 580046 435650 580102
rect 435718 580046 435774 580102
rect 435842 580046 435898 580102
rect 435966 580046 436022 580102
rect 435594 579922 435650 579978
rect 435718 579922 435774 579978
rect 435842 579922 435898 579978
rect 435966 579922 436022 579978
rect 439314 598116 439370 598172
rect 439438 598116 439494 598172
rect 439562 598116 439618 598172
rect 439686 598116 439742 598172
rect 439314 597992 439370 598048
rect 439438 597992 439494 598048
rect 439562 597992 439618 598048
rect 439686 597992 439742 598048
rect 439314 597868 439370 597924
rect 439438 597868 439494 597924
rect 439562 597868 439618 597924
rect 439686 597868 439742 597924
rect 439314 597744 439370 597800
rect 439438 597744 439494 597800
rect 439562 597744 439618 597800
rect 439686 597744 439742 597800
rect 439314 586294 439370 586350
rect 439438 586294 439494 586350
rect 439562 586294 439618 586350
rect 439686 586294 439742 586350
rect 439314 586170 439370 586226
rect 439438 586170 439494 586226
rect 439562 586170 439618 586226
rect 439686 586170 439742 586226
rect 439314 586046 439370 586102
rect 439438 586046 439494 586102
rect 439562 586046 439618 586102
rect 439686 586046 439742 586102
rect 439314 585922 439370 585978
rect 439438 585922 439494 585978
rect 439562 585922 439618 585978
rect 439686 585922 439742 585978
rect 466314 597156 466370 597212
rect 466438 597156 466494 597212
rect 466562 597156 466618 597212
rect 466686 597156 466742 597212
rect 466314 597032 466370 597088
rect 466438 597032 466494 597088
rect 466562 597032 466618 597088
rect 466686 597032 466742 597088
rect 466314 596908 466370 596964
rect 466438 596908 466494 596964
rect 466562 596908 466618 596964
rect 466686 596908 466742 596964
rect 466314 596784 466370 596840
rect 466438 596784 466494 596840
rect 466562 596784 466618 596840
rect 466686 596784 466742 596840
rect 466314 580294 466370 580350
rect 466438 580294 466494 580350
rect 466562 580294 466618 580350
rect 466686 580294 466742 580350
rect 466314 580170 466370 580226
rect 466438 580170 466494 580226
rect 466562 580170 466618 580226
rect 466686 580170 466742 580226
rect 466314 580046 466370 580102
rect 466438 580046 466494 580102
rect 466562 580046 466618 580102
rect 466686 580046 466742 580102
rect 466314 579922 466370 579978
rect 466438 579922 466494 579978
rect 466562 579922 466618 579978
rect 466686 579922 466742 579978
rect 470034 598116 470090 598172
rect 470158 598116 470214 598172
rect 470282 598116 470338 598172
rect 470406 598116 470462 598172
rect 470034 597992 470090 598048
rect 470158 597992 470214 598048
rect 470282 597992 470338 598048
rect 470406 597992 470462 598048
rect 470034 597868 470090 597924
rect 470158 597868 470214 597924
rect 470282 597868 470338 597924
rect 470406 597868 470462 597924
rect 470034 597744 470090 597800
rect 470158 597744 470214 597800
rect 470282 597744 470338 597800
rect 470406 597744 470462 597800
rect 497034 597156 497090 597212
rect 497158 597156 497214 597212
rect 497282 597156 497338 597212
rect 497406 597156 497462 597212
rect 497034 597032 497090 597088
rect 497158 597032 497214 597088
rect 497282 597032 497338 597088
rect 497406 597032 497462 597088
rect 497034 596908 497090 596964
rect 497158 596908 497214 596964
rect 497282 596908 497338 596964
rect 497406 596908 497462 596964
rect 497034 596784 497090 596840
rect 497158 596784 497214 596840
rect 497282 596784 497338 596840
rect 497406 596784 497462 596840
rect 474348 589742 474404 589798
rect 470034 586294 470090 586350
rect 470158 586294 470214 586350
rect 470282 586294 470338 586350
rect 470406 586294 470462 586350
rect 470034 586170 470090 586226
rect 470158 586170 470214 586226
rect 470282 586170 470338 586226
rect 470406 586170 470462 586226
rect 470034 586046 470090 586102
rect 470158 586046 470214 586102
rect 470282 586046 470338 586102
rect 470406 586046 470462 586102
rect 470034 585922 470090 585978
rect 470158 585922 470214 585978
rect 470282 585922 470338 585978
rect 470406 585922 470462 585978
rect 497034 580294 497090 580350
rect 497158 580294 497214 580350
rect 497282 580294 497338 580350
rect 497406 580294 497462 580350
rect 497034 580170 497090 580226
rect 497158 580170 497214 580226
rect 497282 580170 497338 580226
rect 497406 580170 497462 580226
rect 497034 580046 497090 580102
rect 497158 580046 497214 580102
rect 497282 580046 497338 580102
rect 497406 580046 497462 580102
rect 497034 579922 497090 579978
rect 497158 579922 497214 579978
rect 497282 579922 497338 579978
rect 497406 579922 497462 579978
rect 500754 598116 500810 598172
rect 500878 598116 500934 598172
rect 501002 598116 501058 598172
rect 501126 598116 501182 598172
rect 500754 597992 500810 598048
rect 500878 597992 500934 598048
rect 501002 597992 501058 598048
rect 501126 597992 501182 598048
rect 500754 597868 500810 597924
rect 500878 597868 500934 597924
rect 501002 597868 501058 597924
rect 501126 597868 501182 597924
rect 500754 597744 500810 597800
rect 500878 597744 500934 597800
rect 501002 597744 501058 597800
rect 501126 597744 501182 597800
rect 500754 586294 500810 586350
rect 500878 586294 500934 586350
rect 501002 586294 501058 586350
rect 501126 586294 501182 586350
rect 500754 586170 500810 586226
rect 500878 586170 500934 586226
rect 501002 586170 501058 586226
rect 501126 586170 501182 586226
rect 500754 586046 500810 586102
rect 500878 586046 500934 586102
rect 501002 586046 501058 586102
rect 501126 586046 501182 586102
rect 500754 585922 500810 585978
rect 500878 585922 500934 585978
rect 501002 585922 501058 585978
rect 501126 585922 501182 585978
rect 527754 597156 527810 597212
rect 527878 597156 527934 597212
rect 528002 597156 528058 597212
rect 528126 597156 528182 597212
rect 527754 597032 527810 597088
rect 527878 597032 527934 597088
rect 528002 597032 528058 597088
rect 528126 597032 528182 597088
rect 527754 596908 527810 596964
rect 527878 596908 527934 596964
rect 528002 596908 528058 596964
rect 528126 596908 528182 596964
rect 527754 596784 527810 596840
rect 527878 596784 527934 596840
rect 528002 596784 528058 596840
rect 528126 596784 528182 596840
rect 527754 580294 527810 580350
rect 527878 580294 527934 580350
rect 528002 580294 528058 580350
rect 528126 580294 528182 580350
rect 527754 580170 527810 580226
rect 527878 580170 527934 580226
rect 528002 580170 528058 580226
rect 528126 580170 528182 580226
rect 527754 580046 527810 580102
rect 527878 580046 527934 580102
rect 528002 580046 528058 580102
rect 528126 580046 528182 580102
rect 527754 579922 527810 579978
rect 527878 579922 527934 579978
rect 528002 579922 528058 579978
rect 528126 579922 528182 579978
rect 531474 598116 531530 598172
rect 531598 598116 531654 598172
rect 531722 598116 531778 598172
rect 531846 598116 531902 598172
rect 531474 597992 531530 598048
rect 531598 597992 531654 598048
rect 531722 597992 531778 598048
rect 531846 597992 531902 598048
rect 531474 597868 531530 597924
rect 531598 597868 531654 597924
rect 531722 597868 531778 597924
rect 531846 597868 531902 597924
rect 531474 597744 531530 597800
rect 531598 597744 531654 597800
rect 531722 597744 531778 597800
rect 531846 597744 531902 597800
rect 558474 597156 558530 597212
rect 558598 597156 558654 597212
rect 558722 597156 558778 597212
rect 558846 597156 558902 597212
rect 558474 597032 558530 597088
rect 558598 597032 558654 597088
rect 558722 597032 558778 597088
rect 558846 597032 558902 597088
rect 558474 596908 558530 596964
rect 558598 596908 558654 596964
rect 558722 596908 558778 596964
rect 558846 596908 558902 596964
rect 558474 596784 558530 596840
rect 558598 596784 558654 596840
rect 558722 596784 558778 596840
rect 558846 596784 558902 596840
rect 531474 586294 531530 586350
rect 531598 586294 531654 586350
rect 531722 586294 531778 586350
rect 531846 586294 531902 586350
rect 531474 586170 531530 586226
rect 531598 586170 531654 586226
rect 531722 586170 531778 586226
rect 531846 586170 531902 586226
rect 531474 586046 531530 586102
rect 531598 586046 531654 586102
rect 531722 586046 531778 586102
rect 531846 586046 531902 586102
rect 531474 585922 531530 585978
rect 531598 585922 531654 585978
rect 531722 585922 531778 585978
rect 531846 585922 531902 585978
rect 194518 562294 194574 562350
rect 194642 562294 194698 562350
rect 194518 562170 194574 562226
rect 194642 562170 194698 562226
rect 194518 562046 194574 562102
rect 194642 562046 194698 562102
rect 194518 561922 194574 561978
rect 194642 561922 194698 561978
rect 225238 562294 225294 562350
rect 225362 562294 225418 562350
rect 225238 562170 225294 562226
rect 225362 562170 225418 562226
rect 225238 562046 225294 562102
rect 225362 562046 225418 562102
rect 225238 561922 225294 561978
rect 225362 561922 225418 561978
rect 255958 562294 256014 562350
rect 256082 562294 256138 562350
rect 255958 562170 256014 562226
rect 256082 562170 256138 562226
rect 255958 562046 256014 562102
rect 256082 562046 256138 562102
rect 255958 561922 256014 561978
rect 256082 561922 256138 561978
rect 286678 562294 286734 562350
rect 286802 562294 286858 562350
rect 286678 562170 286734 562226
rect 286802 562170 286858 562226
rect 286678 562046 286734 562102
rect 286802 562046 286858 562102
rect 286678 561922 286734 561978
rect 286802 561922 286858 561978
rect 317398 562294 317454 562350
rect 317522 562294 317578 562350
rect 317398 562170 317454 562226
rect 317522 562170 317578 562226
rect 317398 562046 317454 562102
rect 317522 562046 317578 562102
rect 317398 561922 317454 561978
rect 317522 561922 317578 561978
rect 348118 562294 348174 562350
rect 348242 562294 348298 562350
rect 348118 562170 348174 562226
rect 348242 562170 348298 562226
rect 348118 562046 348174 562102
rect 348242 562046 348298 562102
rect 348118 561922 348174 561978
rect 348242 561922 348298 561978
rect 378838 562294 378894 562350
rect 378962 562294 379018 562350
rect 378838 562170 378894 562226
rect 378962 562170 379018 562226
rect 378838 562046 378894 562102
rect 378962 562046 379018 562102
rect 378838 561922 378894 561978
rect 378962 561922 379018 561978
rect 409558 562294 409614 562350
rect 409682 562294 409738 562350
rect 409558 562170 409614 562226
rect 409682 562170 409738 562226
rect 409558 562046 409614 562102
rect 409682 562046 409738 562102
rect 409558 561922 409614 561978
rect 409682 561922 409738 561978
rect 440278 562294 440334 562350
rect 440402 562294 440458 562350
rect 440278 562170 440334 562226
rect 440402 562170 440458 562226
rect 440278 562046 440334 562102
rect 440402 562046 440458 562102
rect 440278 561922 440334 561978
rect 440402 561922 440458 561978
rect 470998 562294 471054 562350
rect 471122 562294 471178 562350
rect 470998 562170 471054 562226
rect 471122 562170 471178 562226
rect 470998 562046 471054 562102
rect 471122 562046 471178 562102
rect 470998 561922 471054 561978
rect 471122 561922 471178 561978
rect 501718 562294 501774 562350
rect 501842 562294 501898 562350
rect 501718 562170 501774 562226
rect 501842 562170 501898 562226
rect 501718 562046 501774 562102
rect 501842 562046 501898 562102
rect 501718 561922 501774 561978
rect 501842 561922 501898 561978
rect 532438 562294 532494 562350
rect 532562 562294 532618 562350
rect 532438 562170 532494 562226
rect 532562 562170 532618 562226
rect 532438 562046 532494 562102
rect 532562 562046 532618 562102
rect 532438 561922 532494 561978
rect 532562 561922 532618 561978
rect 209878 550294 209934 550350
rect 210002 550294 210058 550350
rect 209878 550170 209934 550226
rect 210002 550170 210058 550226
rect 209878 550046 209934 550102
rect 210002 550046 210058 550102
rect 209878 549922 209934 549978
rect 210002 549922 210058 549978
rect 240598 550294 240654 550350
rect 240722 550294 240778 550350
rect 240598 550170 240654 550226
rect 240722 550170 240778 550226
rect 240598 550046 240654 550102
rect 240722 550046 240778 550102
rect 240598 549922 240654 549978
rect 240722 549922 240778 549978
rect 271318 550294 271374 550350
rect 271442 550294 271498 550350
rect 271318 550170 271374 550226
rect 271442 550170 271498 550226
rect 271318 550046 271374 550102
rect 271442 550046 271498 550102
rect 271318 549922 271374 549978
rect 271442 549922 271498 549978
rect 302038 550294 302094 550350
rect 302162 550294 302218 550350
rect 302038 550170 302094 550226
rect 302162 550170 302218 550226
rect 302038 550046 302094 550102
rect 302162 550046 302218 550102
rect 302038 549922 302094 549978
rect 302162 549922 302218 549978
rect 332758 550294 332814 550350
rect 332882 550294 332938 550350
rect 332758 550170 332814 550226
rect 332882 550170 332938 550226
rect 332758 550046 332814 550102
rect 332882 550046 332938 550102
rect 332758 549922 332814 549978
rect 332882 549922 332938 549978
rect 363478 550294 363534 550350
rect 363602 550294 363658 550350
rect 363478 550170 363534 550226
rect 363602 550170 363658 550226
rect 363478 550046 363534 550102
rect 363602 550046 363658 550102
rect 363478 549922 363534 549978
rect 363602 549922 363658 549978
rect 394198 550294 394254 550350
rect 394322 550294 394378 550350
rect 394198 550170 394254 550226
rect 394322 550170 394378 550226
rect 394198 550046 394254 550102
rect 394322 550046 394378 550102
rect 394198 549922 394254 549978
rect 394322 549922 394378 549978
rect 424918 550294 424974 550350
rect 425042 550294 425098 550350
rect 424918 550170 424974 550226
rect 425042 550170 425098 550226
rect 424918 550046 424974 550102
rect 425042 550046 425098 550102
rect 424918 549922 424974 549978
rect 425042 549922 425098 549978
rect 455638 550294 455694 550350
rect 455762 550294 455818 550350
rect 455638 550170 455694 550226
rect 455762 550170 455818 550226
rect 455638 550046 455694 550102
rect 455762 550046 455818 550102
rect 455638 549922 455694 549978
rect 455762 549922 455818 549978
rect 486358 550294 486414 550350
rect 486482 550294 486538 550350
rect 486358 550170 486414 550226
rect 486482 550170 486538 550226
rect 486358 550046 486414 550102
rect 486482 550046 486538 550102
rect 486358 549922 486414 549978
rect 486482 549922 486538 549978
rect 517078 550294 517134 550350
rect 517202 550294 517258 550350
rect 517078 550170 517134 550226
rect 517202 550170 517258 550226
rect 517078 550046 517134 550102
rect 517202 550046 517258 550102
rect 517078 549922 517134 549978
rect 517202 549922 517258 549978
rect 194518 544294 194574 544350
rect 194642 544294 194698 544350
rect 194518 544170 194574 544226
rect 194642 544170 194698 544226
rect 194518 544046 194574 544102
rect 194642 544046 194698 544102
rect 194518 543922 194574 543978
rect 194642 543922 194698 543978
rect 225238 544294 225294 544350
rect 225362 544294 225418 544350
rect 225238 544170 225294 544226
rect 225362 544170 225418 544226
rect 225238 544046 225294 544102
rect 225362 544046 225418 544102
rect 225238 543922 225294 543978
rect 225362 543922 225418 543978
rect 255958 544294 256014 544350
rect 256082 544294 256138 544350
rect 255958 544170 256014 544226
rect 256082 544170 256138 544226
rect 255958 544046 256014 544102
rect 256082 544046 256138 544102
rect 255958 543922 256014 543978
rect 256082 543922 256138 543978
rect 286678 544294 286734 544350
rect 286802 544294 286858 544350
rect 286678 544170 286734 544226
rect 286802 544170 286858 544226
rect 286678 544046 286734 544102
rect 286802 544046 286858 544102
rect 286678 543922 286734 543978
rect 286802 543922 286858 543978
rect 317398 544294 317454 544350
rect 317522 544294 317578 544350
rect 317398 544170 317454 544226
rect 317522 544170 317578 544226
rect 317398 544046 317454 544102
rect 317522 544046 317578 544102
rect 317398 543922 317454 543978
rect 317522 543922 317578 543978
rect 348118 544294 348174 544350
rect 348242 544294 348298 544350
rect 348118 544170 348174 544226
rect 348242 544170 348298 544226
rect 348118 544046 348174 544102
rect 348242 544046 348298 544102
rect 348118 543922 348174 543978
rect 348242 543922 348298 543978
rect 378838 544294 378894 544350
rect 378962 544294 379018 544350
rect 378838 544170 378894 544226
rect 378962 544170 379018 544226
rect 378838 544046 378894 544102
rect 378962 544046 379018 544102
rect 378838 543922 378894 543978
rect 378962 543922 379018 543978
rect 409558 544294 409614 544350
rect 409682 544294 409738 544350
rect 409558 544170 409614 544226
rect 409682 544170 409738 544226
rect 409558 544046 409614 544102
rect 409682 544046 409738 544102
rect 409558 543922 409614 543978
rect 409682 543922 409738 543978
rect 440278 544294 440334 544350
rect 440402 544294 440458 544350
rect 440278 544170 440334 544226
rect 440402 544170 440458 544226
rect 440278 544046 440334 544102
rect 440402 544046 440458 544102
rect 440278 543922 440334 543978
rect 440402 543922 440458 543978
rect 470998 544294 471054 544350
rect 471122 544294 471178 544350
rect 470998 544170 471054 544226
rect 471122 544170 471178 544226
rect 470998 544046 471054 544102
rect 471122 544046 471178 544102
rect 470998 543922 471054 543978
rect 471122 543922 471178 543978
rect 501718 544294 501774 544350
rect 501842 544294 501898 544350
rect 501718 544170 501774 544226
rect 501842 544170 501898 544226
rect 501718 544046 501774 544102
rect 501842 544046 501898 544102
rect 501718 543922 501774 543978
rect 501842 543922 501898 543978
rect 532438 544294 532494 544350
rect 532562 544294 532618 544350
rect 532438 544170 532494 544226
rect 532562 544170 532618 544226
rect 532438 544046 532494 544102
rect 532562 544046 532618 544102
rect 532438 543922 532494 543978
rect 532562 543922 532618 543978
rect 209878 532294 209934 532350
rect 210002 532294 210058 532350
rect 209878 532170 209934 532226
rect 210002 532170 210058 532226
rect 209878 532046 209934 532102
rect 210002 532046 210058 532102
rect 209878 531922 209934 531978
rect 210002 531922 210058 531978
rect 240598 532294 240654 532350
rect 240722 532294 240778 532350
rect 240598 532170 240654 532226
rect 240722 532170 240778 532226
rect 240598 532046 240654 532102
rect 240722 532046 240778 532102
rect 240598 531922 240654 531978
rect 240722 531922 240778 531978
rect 271318 532294 271374 532350
rect 271442 532294 271498 532350
rect 271318 532170 271374 532226
rect 271442 532170 271498 532226
rect 271318 532046 271374 532102
rect 271442 532046 271498 532102
rect 271318 531922 271374 531978
rect 271442 531922 271498 531978
rect 302038 532294 302094 532350
rect 302162 532294 302218 532350
rect 302038 532170 302094 532226
rect 302162 532170 302218 532226
rect 302038 532046 302094 532102
rect 302162 532046 302218 532102
rect 302038 531922 302094 531978
rect 302162 531922 302218 531978
rect 332758 532294 332814 532350
rect 332882 532294 332938 532350
rect 332758 532170 332814 532226
rect 332882 532170 332938 532226
rect 332758 532046 332814 532102
rect 332882 532046 332938 532102
rect 332758 531922 332814 531978
rect 332882 531922 332938 531978
rect 363478 532294 363534 532350
rect 363602 532294 363658 532350
rect 363478 532170 363534 532226
rect 363602 532170 363658 532226
rect 363478 532046 363534 532102
rect 363602 532046 363658 532102
rect 363478 531922 363534 531978
rect 363602 531922 363658 531978
rect 394198 532294 394254 532350
rect 394322 532294 394378 532350
rect 394198 532170 394254 532226
rect 394322 532170 394378 532226
rect 394198 532046 394254 532102
rect 394322 532046 394378 532102
rect 394198 531922 394254 531978
rect 394322 531922 394378 531978
rect 424918 532294 424974 532350
rect 425042 532294 425098 532350
rect 424918 532170 424974 532226
rect 425042 532170 425098 532226
rect 424918 532046 424974 532102
rect 425042 532046 425098 532102
rect 424918 531922 424974 531978
rect 425042 531922 425098 531978
rect 455638 532294 455694 532350
rect 455762 532294 455818 532350
rect 455638 532170 455694 532226
rect 455762 532170 455818 532226
rect 455638 532046 455694 532102
rect 455762 532046 455818 532102
rect 455638 531922 455694 531978
rect 455762 531922 455818 531978
rect 486358 532294 486414 532350
rect 486482 532294 486538 532350
rect 486358 532170 486414 532226
rect 486482 532170 486538 532226
rect 486358 532046 486414 532102
rect 486482 532046 486538 532102
rect 486358 531922 486414 531978
rect 486482 531922 486538 531978
rect 517078 532294 517134 532350
rect 517202 532294 517258 532350
rect 517078 532170 517134 532226
rect 517202 532170 517258 532226
rect 517078 532046 517134 532102
rect 517202 532046 517258 532102
rect 517078 531922 517134 531978
rect 517202 531922 517258 531978
rect 194518 526294 194574 526350
rect 194642 526294 194698 526350
rect 194518 526170 194574 526226
rect 194642 526170 194698 526226
rect 194518 526046 194574 526102
rect 194642 526046 194698 526102
rect 194518 525922 194574 525978
rect 194642 525922 194698 525978
rect 225238 526294 225294 526350
rect 225362 526294 225418 526350
rect 225238 526170 225294 526226
rect 225362 526170 225418 526226
rect 225238 526046 225294 526102
rect 225362 526046 225418 526102
rect 225238 525922 225294 525978
rect 225362 525922 225418 525978
rect 255958 526294 256014 526350
rect 256082 526294 256138 526350
rect 255958 526170 256014 526226
rect 256082 526170 256138 526226
rect 255958 526046 256014 526102
rect 256082 526046 256138 526102
rect 255958 525922 256014 525978
rect 256082 525922 256138 525978
rect 286678 526294 286734 526350
rect 286802 526294 286858 526350
rect 286678 526170 286734 526226
rect 286802 526170 286858 526226
rect 286678 526046 286734 526102
rect 286802 526046 286858 526102
rect 286678 525922 286734 525978
rect 286802 525922 286858 525978
rect 317398 526294 317454 526350
rect 317522 526294 317578 526350
rect 317398 526170 317454 526226
rect 317522 526170 317578 526226
rect 317398 526046 317454 526102
rect 317522 526046 317578 526102
rect 317398 525922 317454 525978
rect 317522 525922 317578 525978
rect 348118 526294 348174 526350
rect 348242 526294 348298 526350
rect 348118 526170 348174 526226
rect 348242 526170 348298 526226
rect 348118 526046 348174 526102
rect 348242 526046 348298 526102
rect 348118 525922 348174 525978
rect 348242 525922 348298 525978
rect 378838 526294 378894 526350
rect 378962 526294 379018 526350
rect 378838 526170 378894 526226
rect 378962 526170 379018 526226
rect 378838 526046 378894 526102
rect 378962 526046 379018 526102
rect 378838 525922 378894 525978
rect 378962 525922 379018 525978
rect 409558 526294 409614 526350
rect 409682 526294 409738 526350
rect 409558 526170 409614 526226
rect 409682 526170 409738 526226
rect 409558 526046 409614 526102
rect 409682 526046 409738 526102
rect 409558 525922 409614 525978
rect 409682 525922 409738 525978
rect 440278 526294 440334 526350
rect 440402 526294 440458 526350
rect 440278 526170 440334 526226
rect 440402 526170 440458 526226
rect 440278 526046 440334 526102
rect 440402 526046 440458 526102
rect 440278 525922 440334 525978
rect 440402 525922 440458 525978
rect 470998 526294 471054 526350
rect 471122 526294 471178 526350
rect 470998 526170 471054 526226
rect 471122 526170 471178 526226
rect 470998 526046 471054 526102
rect 471122 526046 471178 526102
rect 470998 525922 471054 525978
rect 471122 525922 471178 525978
rect 501718 526294 501774 526350
rect 501842 526294 501898 526350
rect 501718 526170 501774 526226
rect 501842 526170 501898 526226
rect 501718 526046 501774 526102
rect 501842 526046 501898 526102
rect 501718 525922 501774 525978
rect 501842 525922 501898 525978
rect 532438 526294 532494 526350
rect 532562 526294 532618 526350
rect 532438 526170 532494 526226
rect 532562 526170 532618 526226
rect 532438 526046 532494 526102
rect 532562 526046 532618 526102
rect 532438 525922 532494 525978
rect 532562 525922 532618 525978
rect 209878 514294 209934 514350
rect 210002 514294 210058 514350
rect 209878 514170 209934 514226
rect 210002 514170 210058 514226
rect 209878 514046 209934 514102
rect 210002 514046 210058 514102
rect 209878 513922 209934 513978
rect 210002 513922 210058 513978
rect 240598 514294 240654 514350
rect 240722 514294 240778 514350
rect 240598 514170 240654 514226
rect 240722 514170 240778 514226
rect 240598 514046 240654 514102
rect 240722 514046 240778 514102
rect 240598 513922 240654 513978
rect 240722 513922 240778 513978
rect 271318 514294 271374 514350
rect 271442 514294 271498 514350
rect 271318 514170 271374 514226
rect 271442 514170 271498 514226
rect 271318 514046 271374 514102
rect 271442 514046 271498 514102
rect 271318 513922 271374 513978
rect 271442 513922 271498 513978
rect 302038 514294 302094 514350
rect 302162 514294 302218 514350
rect 302038 514170 302094 514226
rect 302162 514170 302218 514226
rect 302038 514046 302094 514102
rect 302162 514046 302218 514102
rect 302038 513922 302094 513978
rect 302162 513922 302218 513978
rect 332758 514294 332814 514350
rect 332882 514294 332938 514350
rect 332758 514170 332814 514226
rect 332882 514170 332938 514226
rect 332758 514046 332814 514102
rect 332882 514046 332938 514102
rect 332758 513922 332814 513978
rect 332882 513922 332938 513978
rect 363478 514294 363534 514350
rect 363602 514294 363658 514350
rect 363478 514170 363534 514226
rect 363602 514170 363658 514226
rect 363478 514046 363534 514102
rect 363602 514046 363658 514102
rect 363478 513922 363534 513978
rect 363602 513922 363658 513978
rect 394198 514294 394254 514350
rect 394322 514294 394378 514350
rect 394198 514170 394254 514226
rect 394322 514170 394378 514226
rect 394198 514046 394254 514102
rect 394322 514046 394378 514102
rect 394198 513922 394254 513978
rect 394322 513922 394378 513978
rect 424918 514294 424974 514350
rect 425042 514294 425098 514350
rect 424918 514170 424974 514226
rect 425042 514170 425098 514226
rect 424918 514046 424974 514102
rect 425042 514046 425098 514102
rect 424918 513922 424974 513978
rect 425042 513922 425098 513978
rect 455638 514294 455694 514350
rect 455762 514294 455818 514350
rect 455638 514170 455694 514226
rect 455762 514170 455818 514226
rect 455638 514046 455694 514102
rect 455762 514046 455818 514102
rect 455638 513922 455694 513978
rect 455762 513922 455818 513978
rect 486358 514294 486414 514350
rect 486482 514294 486538 514350
rect 486358 514170 486414 514226
rect 486482 514170 486538 514226
rect 486358 514046 486414 514102
rect 486482 514046 486538 514102
rect 486358 513922 486414 513978
rect 486482 513922 486538 513978
rect 517078 514294 517134 514350
rect 517202 514294 517258 514350
rect 517078 514170 517134 514226
rect 517202 514170 517258 514226
rect 517078 514046 517134 514102
rect 517202 514046 517258 514102
rect 517078 513922 517134 513978
rect 517202 513922 517258 513978
rect 194518 508294 194574 508350
rect 194642 508294 194698 508350
rect 194518 508170 194574 508226
rect 194642 508170 194698 508226
rect 194518 508046 194574 508102
rect 194642 508046 194698 508102
rect 194518 507922 194574 507978
rect 194642 507922 194698 507978
rect 225238 508294 225294 508350
rect 225362 508294 225418 508350
rect 225238 508170 225294 508226
rect 225362 508170 225418 508226
rect 225238 508046 225294 508102
rect 225362 508046 225418 508102
rect 225238 507922 225294 507978
rect 225362 507922 225418 507978
rect 255958 508294 256014 508350
rect 256082 508294 256138 508350
rect 255958 508170 256014 508226
rect 256082 508170 256138 508226
rect 255958 508046 256014 508102
rect 256082 508046 256138 508102
rect 255958 507922 256014 507978
rect 256082 507922 256138 507978
rect 286678 508294 286734 508350
rect 286802 508294 286858 508350
rect 286678 508170 286734 508226
rect 286802 508170 286858 508226
rect 286678 508046 286734 508102
rect 286802 508046 286858 508102
rect 286678 507922 286734 507978
rect 286802 507922 286858 507978
rect 317398 508294 317454 508350
rect 317522 508294 317578 508350
rect 317398 508170 317454 508226
rect 317522 508170 317578 508226
rect 317398 508046 317454 508102
rect 317522 508046 317578 508102
rect 317398 507922 317454 507978
rect 317522 507922 317578 507978
rect 348118 508294 348174 508350
rect 348242 508294 348298 508350
rect 348118 508170 348174 508226
rect 348242 508170 348298 508226
rect 348118 508046 348174 508102
rect 348242 508046 348298 508102
rect 348118 507922 348174 507978
rect 348242 507922 348298 507978
rect 378838 508294 378894 508350
rect 378962 508294 379018 508350
rect 378838 508170 378894 508226
rect 378962 508170 379018 508226
rect 378838 508046 378894 508102
rect 378962 508046 379018 508102
rect 378838 507922 378894 507978
rect 378962 507922 379018 507978
rect 409558 508294 409614 508350
rect 409682 508294 409738 508350
rect 409558 508170 409614 508226
rect 409682 508170 409738 508226
rect 409558 508046 409614 508102
rect 409682 508046 409738 508102
rect 409558 507922 409614 507978
rect 409682 507922 409738 507978
rect 440278 508294 440334 508350
rect 440402 508294 440458 508350
rect 440278 508170 440334 508226
rect 440402 508170 440458 508226
rect 440278 508046 440334 508102
rect 440402 508046 440458 508102
rect 440278 507922 440334 507978
rect 440402 507922 440458 507978
rect 470998 508294 471054 508350
rect 471122 508294 471178 508350
rect 470998 508170 471054 508226
rect 471122 508170 471178 508226
rect 470998 508046 471054 508102
rect 471122 508046 471178 508102
rect 470998 507922 471054 507978
rect 471122 507922 471178 507978
rect 501718 508294 501774 508350
rect 501842 508294 501898 508350
rect 501718 508170 501774 508226
rect 501842 508170 501898 508226
rect 501718 508046 501774 508102
rect 501842 508046 501898 508102
rect 501718 507922 501774 507978
rect 501842 507922 501898 507978
rect 532438 508294 532494 508350
rect 532562 508294 532618 508350
rect 532438 508170 532494 508226
rect 532562 508170 532618 508226
rect 532438 508046 532494 508102
rect 532562 508046 532618 508102
rect 532438 507922 532494 507978
rect 532562 507922 532618 507978
rect 209878 496294 209934 496350
rect 210002 496294 210058 496350
rect 209878 496170 209934 496226
rect 210002 496170 210058 496226
rect 209878 496046 209934 496102
rect 210002 496046 210058 496102
rect 209878 495922 209934 495978
rect 210002 495922 210058 495978
rect 240598 496294 240654 496350
rect 240722 496294 240778 496350
rect 240598 496170 240654 496226
rect 240722 496170 240778 496226
rect 240598 496046 240654 496102
rect 240722 496046 240778 496102
rect 240598 495922 240654 495978
rect 240722 495922 240778 495978
rect 271318 496294 271374 496350
rect 271442 496294 271498 496350
rect 271318 496170 271374 496226
rect 271442 496170 271498 496226
rect 271318 496046 271374 496102
rect 271442 496046 271498 496102
rect 271318 495922 271374 495978
rect 271442 495922 271498 495978
rect 302038 496294 302094 496350
rect 302162 496294 302218 496350
rect 302038 496170 302094 496226
rect 302162 496170 302218 496226
rect 302038 496046 302094 496102
rect 302162 496046 302218 496102
rect 302038 495922 302094 495978
rect 302162 495922 302218 495978
rect 332758 496294 332814 496350
rect 332882 496294 332938 496350
rect 332758 496170 332814 496226
rect 332882 496170 332938 496226
rect 332758 496046 332814 496102
rect 332882 496046 332938 496102
rect 332758 495922 332814 495978
rect 332882 495922 332938 495978
rect 363478 496294 363534 496350
rect 363602 496294 363658 496350
rect 363478 496170 363534 496226
rect 363602 496170 363658 496226
rect 363478 496046 363534 496102
rect 363602 496046 363658 496102
rect 363478 495922 363534 495978
rect 363602 495922 363658 495978
rect 394198 496294 394254 496350
rect 394322 496294 394378 496350
rect 394198 496170 394254 496226
rect 394322 496170 394378 496226
rect 394198 496046 394254 496102
rect 394322 496046 394378 496102
rect 394198 495922 394254 495978
rect 394322 495922 394378 495978
rect 424918 496294 424974 496350
rect 425042 496294 425098 496350
rect 424918 496170 424974 496226
rect 425042 496170 425098 496226
rect 424918 496046 424974 496102
rect 425042 496046 425098 496102
rect 424918 495922 424974 495978
rect 425042 495922 425098 495978
rect 455638 496294 455694 496350
rect 455762 496294 455818 496350
rect 455638 496170 455694 496226
rect 455762 496170 455818 496226
rect 455638 496046 455694 496102
rect 455762 496046 455818 496102
rect 455638 495922 455694 495978
rect 455762 495922 455818 495978
rect 486358 496294 486414 496350
rect 486482 496294 486538 496350
rect 486358 496170 486414 496226
rect 486482 496170 486538 496226
rect 486358 496046 486414 496102
rect 486482 496046 486538 496102
rect 486358 495922 486414 495978
rect 486482 495922 486538 495978
rect 517078 496294 517134 496350
rect 517202 496294 517258 496350
rect 517078 496170 517134 496226
rect 517202 496170 517258 496226
rect 517078 496046 517134 496102
rect 517202 496046 517258 496102
rect 517078 495922 517134 495978
rect 517202 495922 517258 495978
rect 194518 490294 194574 490350
rect 194642 490294 194698 490350
rect 194518 490170 194574 490226
rect 194642 490170 194698 490226
rect 194518 490046 194574 490102
rect 194642 490046 194698 490102
rect 194518 489922 194574 489978
rect 194642 489922 194698 489978
rect 225238 490294 225294 490350
rect 225362 490294 225418 490350
rect 225238 490170 225294 490226
rect 225362 490170 225418 490226
rect 225238 490046 225294 490102
rect 225362 490046 225418 490102
rect 225238 489922 225294 489978
rect 225362 489922 225418 489978
rect 255958 490294 256014 490350
rect 256082 490294 256138 490350
rect 255958 490170 256014 490226
rect 256082 490170 256138 490226
rect 255958 490046 256014 490102
rect 256082 490046 256138 490102
rect 255958 489922 256014 489978
rect 256082 489922 256138 489978
rect 286678 490294 286734 490350
rect 286802 490294 286858 490350
rect 286678 490170 286734 490226
rect 286802 490170 286858 490226
rect 286678 490046 286734 490102
rect 286802 490046 286858 490102
rect 286678 489922 286734 489978
rect 286802 489922 286858 489978
rect 317398 490294 317454 490350
rect 317522 490294 317578 490350
rect 317398 490170 317454 490226
rect 317522 490170 317578 490226
rect 317398 490046 317454 490102
rect 317522 490046 317578 490102
rect 317398 489922 317454 489978
rect 317522 489922 317578 489978
rect 348118 490294 348174 490350
rect 348242 490294 348298 490350
rect 348118 490170 348174 490226
rect 348242 490170 348298 490226
rect 348118 490046 348174 490102
rect 348242 490046 348298 490102
rect 348118 489922 348174 489978
rect 348242 489922 348298 489978
rect 378838 490294 378894 490350
rect 378962 490294 379018 490350
rect 378838 490170 378894 490226
rect 378962 490170 379018 490226
rect 378838 490046 378894 490102
rect 378962 490046 379018 490102
rect 378838 489922 378894 489978
rect 378962 489922 379018 489978
rect 409558 490294 409614 490350
rect 409682 490294 409738 490350
rect 409558 490170 409614 490226
rect 409682 490170 409738 490226
rect 409558 490046 409614 490102
rect 409682 490046 409738 490102
rect 409558 489922 409614 489978
rect 409682 489922 409738 489978
rect 440278 490294 440334 490350
rect 440402 490294 440458 490350
rect 440278 490170 440334 490226
rect 440402 490170 440458 490226
rect 440278 490046 440334 490102
rect 440402 490046 440458 490102
rect 440278 489922 440334 489978
rect 440402 489922 440458 489978
rect 470998 490294 471054 490350
rect 471122 490294 471178 490350
rect 470998 490170 471054 490226
rect 471122 490170 471178 490226
rect 470998 490046 471054 490102
rect 471122 490046 471178 490102
rect 470998 489922 471054 489978
rect 471122 489922 471178 489978
rect 501718 490294 501774 490350
rect 501842 490294 501898 490350
rect 501718 490170 501774 490226
rect 501842 490170 501898 490226
rect 501718 490046 501774 490102
rect 501842 490046 501898 490102
rect 501718 489922 501774 489978
rect 501842 489922 501898 489978
rect 532438 490294 532494 490350
rect 532562 490294 532618 490350
rect 532438 490170 532494 490226
rect 532562 490170 532618 490226
rect 532438 490046 532494 490102
rect 532562 490046 532618 490102
rect 532438 489922 532494 489978
rect 532562 489922 532618 489978
rect 209878 478294 209934 478350
rect 210002 478294 210058 478350
rect 209878 478170 209934 478226
rect 210002 478170 210058 478226
rect 209878 478046 209934 478102
rect 210002 478046 210058 478102
rect 209878 477922 209934 477978
rect 210002 477922 210058 477978
rect 240598 478294 240654 478350
rect 240722 478294 240778 478350
rect 240598 478170 240654 478226
rect 240722 478170 240778 478226
rect 240598 478046 240654 478102
rect 240722 478046 240778 478102
rect 240598 477922 240654 477978
rect 240722 477922 240778 477978
rect 271318 478294 271374 478350
rect 271442 478294 271498 478350
rect 271318 478170 271374 478226
rect 271442 478170 271498 478226
rect 271318 478046 271374 478102
rect 271442 478046 271498 478102
rect 271318 477922 271374 477978
rect 271442 477922 271498 477978
rect 302038 478294 302094 478350
rect 302162 478294 302218 478350
rect 302038 478170 302094 478226
rect 302162 478170 302218 478226
rect 302038 478046 302094 478102
rect 302162 478046 302218 478102
rect 302038 477922 302094 477978
rect 302162 477922 302218 477978
rect 332758 478294 332814 478350
rect 332882 478294 332938 478350
rect 332758 478170 332814 478226
rect 332882 478170 332938 478226
rect 332758 478046 332814 478102
rect 332882 478046 332938 478102
rect 332758 477922 332814 477978
rect 332882 477922 332938 477978
rect 363478 478294 363534 478350
rect 363602 478294 363658 478350
rect 363478 478170 363534 478226
rect 363602 478170 363658 478226
rect 363478 478046 363534 478102
rect 363602 478046 363658 478102
rect 363478 477922 363534 477978
rect 363602 477922 363658 477978
rect 394198 478294 394254 478350
rect 394322 478294 394378 478350
rect 394198 478170 394254 478226
rect 394322 478170 394378 478226
rect 394198 478046 394254 478102
rect 394322 478046 394378 478102
rect 394198 477922 394254 477978
rect 394322 477922 394378 477978
rect 424918 478294 424974 478350
rect 425042 478294 425098 478350
rect 424918 478170 424974 478226
rect 425042 478170 425098 478226
rect 424918 478046 424974 478102
rect 425042 478046 425098 478102
rect 424918 477922 424974 477978
rect 425042 477922 425098 477978
rect 455638 478294 455694 478350
rect 455762 478294 455818 478350
rect 455638 478170 455694 478226
rect 455762 478170 455818 478226
rect 455638 478046 455694 478102
rect 455762 478046 455818 478102
rect 455638 477922 455694 477978
rect 455762 477922 455818 477978
rect 486358 478294 486414 478350
rect 486482 478294 486538 478350
rect 486358 478170 486414 478226
rect 486482 478170 486538 478226
rect 486358 478046 486414 478102
rect 486482 478046 486538 478102
rect 486358 477922 486414 477978
rect 486482 477922 486538 477978
rect 517078 478294 517134 478350
rect 517202 478294 517258 478350
rect 517078 478170 517134 478226
rect 517202 478170 517258 478226
rect 517078 478046 517134 478102
rect 517202 478046 517258 478102
rect 517078 477922 517134 477978
rect 517202 477922 517258 477978
rect 194518 472294 194574 472350
rect 194642 472294 194698 472350
rect 194518 472170 194574 472226
rect 194642 472170 194698 472226
rect 194518 472046 194574 472102
rect 194642 472046 194698 472102
rect 194518 471922 194574 471978
rect 194642 471922 194698 471978
rect 225238 472294 225294 472350
rect 225362 472294 225418 472350
rect 225238 472170 225294 472226
rect 225362 472170 225418 472226
rect 225238 472046 225294 472102
rect 225362 472046 225418 472102
rect 225238 471922 225294 471978
rect 225362 471922 225418 471978
rect 255958 472294 256014 472350
rect 256082 472294 256138 472350
rect 255958 472170 256014 472226
rect 256082 472170 256138 472226
rect 255958 472046 256014 472102
rect 256082 472046 256138 472102
rect 255958 471922 256014 471978
rect 256082 471922 256138 471978
rect 286678 472294 286734 472350
rect 286802 472294 286858 472350
rect 286678 472170 286734 472226
rect 286802 472170 286858 472226
rect 286678 472046 286734 472102
rect 286802 472046 286858 472102
rect 286678 471922 286734 471978
rect 286802 471922 286858 471978
rect 317398 472294 317454 472350
rect 317522 472294 317578 472350
rect 317398 472170 317454 472226
rect 317522 472170 317578 472226
rect 317398 472046 317454 472102
rect 317522 472046 317578 472102
rect 317398 471922 317454 471978
rect 317522 471922 317578 471978
rect 348118 472294 348174 472350
rect 348242 472294 348298 472350
rect 348118 472170 348174 472226
rect 348242 472170 348298 472226
rect 348118 472046 348174 472102
rect 348242 472046 348298 472102
rect 348118 471922 348174 471978
rect 348242 471922 348298 471978
rect 378838 472294 378894 472350
rect 378962 472294 379018 472350
rect 378838 472170 378894 472226
rect 378962 472170 379018 472226
rect 378838 472046 378894 472102
rect 378962 472046 379018 472102
rect 378838 471922 378894 471978
rect 378962 471922 379018 471978
rect 409558 472294 409614 472350
rect 409682 472294 409738 472350
rect 409558 472170 409614 472226
rect 409682 472170 409738 472226
rect 409558 472046 409614 472102
rect 409682 472046 409738 472102
rect 409558 471922 409614 471978
rect 409682 471922 409738 471978
rect 440278 472294 440334 472350
rect 440402 472294 440458 472350
rect 440278 472170 440334 472226
rect 440402 472170 440458 472226
rect 440278 472046 440334 472102
rect 440402 472046 440458 472102
rect 440278 471922 440334 471978
rect 440402 471922 440458 471978
rect 470998 472294 471054 472350
rect 471122 472294 471178 472350
rect 470998 472170 471054 472226
rect 471122 472170 471178 472226
rect 470998 472046 471054 472102
rect 471122 472046 471178 472102
rect 470998 471922 471054 471978
rect 471122 471922 471178 471978
rect 501718 472294 501774 472350
rect 501842 472294 501898 472350
rect 501718 472170 501774 472226
rect 501842 472170 501898 472226
rect 501718 472046 501774 472102
rect 501842 472046 501898 472102
rect 501718 471922 501774 471978
rect 501842 471922 501898 471978
rect 532438 472294 532494 472350
rect 532562 472294 532618 472350
rect 532438 472170 532494 472226
rect 532562 472170 532618 472226
rect 532438 472046 532494 472102
rect 532562 472046 532618 472102
rect 532438 471922 532494 471978
rect 532562 471922 532618 471978
rect 209878 460294 209934 460350
rect 210002 460294 210058 460350
rect 209878 460170 209934 460226
rect 210002 460170 210058 460226
rect 209878 460046 209934 460102
rect 210002 460046 210058 460102
rect 209878 459922 209934 459978
rect 210002 459922 210058 459978
rect 240598 460294 240654 460350
rect 240722 460294 240778 460350
rect 240598 460170 240654 460226
rect 240722 460170 240778 460226
rect 240598 460046 240654 460102
rect 240722 460046 240778 460102
rect 240598 459922 240654 459978
rect 240722 459922 240778 459978
rect 271318 460294 271374 460350
rect 271442 460294 271498 460350
rect 271318 460170 271374 460226
rect 271442 460170 271498 460226
rect 271318 460046 271374 460102
rect 271442 460046 271498 460102
rect 271318 459922 271374 459978
rect 271442 459922 271498 459978
rect 302038 460294 302094 460350
rect 302162 460294 302218 460350
rect 302038 460170 302094 460226
rect 302162 460170 302218 460226
rect 302038 460046 302094 460102
rect 302162 460046 302218 460102
rect 302038 459922 302094 459978
rect 302162 459922 302218 459978
rect 332758 460294 332814 460350
rect 332882 460294 332938 460350
rect 332758 460170 332814 460226
rect 332882 460170 332938 460226
rect 332758 460046 332814 460102
rect 332882 460046 332938 460102
rect 332758 459922 332814 459978
rect 332882 459922 332938 459978
rect 363478 460294 363534 460350
rect 363602 460294 363658 460350
rect 363478 460170 363534 460226
rect 363602 460170 363658 460226
rect 363478 460046 363534 460102
rect 363602 460046 363658 460102
rect 363478 459922 363534 459978
rect 363602 459922 363658 459978
rect 394198 460294 394254 460350
rect 394322 460294 394378 460350
rect 394198 460170 394254 460226
rect 394322 460170 394378 460226
rect 394198 460046 394254 460102
rect 394322 460046 394378 460102
rect 394198 459922 394254 459978
rect 394322 459922 394378 459978
rect 424918 460294 424974 460350
rect 425042 460294 425098 460350
rect 424918 460170 424974 460226
rect 425042 460170 425098 460226
rect 424918 460046 424974 460102
rect 425042 460046 425098 460102
rect 424918 459922 424974 459978
rect 425042 459922 425098 459978
rect 455638 460294 455694 460350
rect 455762 460294 455818 460350
rect 455638 460170 455694 460226
rect 455762 460170 455818 460226
rect 455638 460046 455694 460102
rect 455762 460046 455818 460102
rect 455638 459922 455694 459978
rect 455762 459922 455818 459978
rect 486358 460294 486414 460350
rect 486482 460294 486538 460350
rect 486358 460170 486414 460226
rect 486482 460170 486538 460226
rect 486358 460046 486414 460102
rect 486482 460046 486538 460102
rect 486358 459922 486414 459978
rect 486482 459922 486538 459978
rect 517078 460294 517134 460350
rect 517202 460294 517258 460350
rect 517078 460170 517134 460226
rect 517202 460170 517258 460226
rect 517078 460046 517134 460102
rect 517202 460046 517258 460102
rect 517078 459922 517134 459978
rect 517202 459922 517258 459978
rect 194518 454294 194574 454350
rect 194642 454294 194698 454350
rect 194518 454170 194574 454226
rect 194642 454170 194698 454226
rect 194518 454046 194574 454102
rect 194642 454046 194698 454102
rect 194518 453922 194574 453978
rect 194642 453922 194698 453978
rect 225238 454294 225294 454350
rect 225362 454294 225418 454350
rect 225238 454170 225294 454226
rect 225362 454170 225418 454226
rect 225238 454046 225294 454102
rect 225362 454046 225418 454102
rect 225238 453922 225294 453978
rect 225362 453922 225418 453978
rect 255958 454294 256014 454350
rect 256082 454294 256138 454350
rect 255958 454170 256014 454226
rect 256082 454170 256138 454226
rect 255958 454046 256014 454102
rect 256082 454046 256138 454102
rect 255958 453922 256014 453978
rect 256082 453922 256138 453978
rect 286678 454294 286734 454350
rect 286802 454294 286858 454350
rect 286678 454170 286734 454226
rect 286802 454170 286858 454226
rect 286678 454046 286734 454102
rect 286802 454046 286858 454102
rect 286678 453922 286734 453978
rect 286802 453922 286858 453978
rect 317398 454294 317454 454350
rect 317522 454294 317578 454350
rect 317398 454170 317454 454226
rect 317522 454170 317578 454226
rect 317398 454046 317454 454102
rect 317522 454046 317578 454102
rect 317398 453922 317454 453978
rect 317522 453922 317578 453978
rect 348118 454294 348174 454350
rect 348242 454294 348298 454350
rect 348118 454170 348174 454226
rect 348242 454170 348298 454226
rect 348118 454046 348174 454102
rect 348242 454046 348298 454102
rect 348118 453922 348174 453978
rect 348242 453922 348298 453978
rect 378838 454294 378894 454350
rect 378962 454294 379018 454350
rect 378838 454170 378894 454226
rect 378962 454170 379018 454226
rect 378838 454046 378894 454102
rect 378962 454046 379018 454102
rect 378838 453922 378894 453978
rect 378962 453922 379018 453978
rect 409558 454294 409614 454350
rect 409682 454294 409738 454350
rect 409558 454170 409614 454226
rect 409682 454170 409738 454226
rect 409558 454046 409614 454102
rect 409682 454046 409738 454102
rect 409558 453922 409614 453978
rect 409682 453922 409738 453978
rect 440278 454294 440334 454350
rect 440402 454294 440458 454350
rect 440278 454170 440334 454226
rect 440402 454170 440458 454226
rect 440278 454046 440334 454102
rect 440402 454046 440458 454102
rect 440278 453922 440334 453978
rect 440402 453922 440458 453978
rect 470998 454294 471054 454350
rect 471122 454294 471178 454350
rect 470998 454170 471054 454226
rect 471122 454170 471178 454226
rect 470998 454046 471054 454102
rect 471122 454046 471178 454102
rect 470998 453922 471054 453978
rect 471122 453922 471178 453978
rect 501718 454294 501774 454350
rect 501842 454294 501898 454350
rect 501718 454170 501774 454226
rect 501842 454170 501898 454226
rect 501718 454046 501774 454102
rect 501842 454046 501898 454102
rect 501718 453922 501774 453978
rect 501842 453922 501898 453978
rect 532438 454294 532494 454350
rect 532562 454294 532618 454350
rect 532438 454170 532494 454226
rect 532562 454170 532618 454226
rect 532438 454046 532494 454102
rect 532562 454046 532618 454102
rect 532438 453922 532494 453978
rect 532562 453922 532618 453978
rect 209878 442294 209934 442350
rect 210002 442294 210058 442350
rect 209878 442170 209934 442226
rect 210002 442170 210058 442226
rect 209878 442046 209934 442102
rect 210002 442046 210058 442102
rect 209878 441922 209934 441978
rect 210002 441922 210058 441978
rect 240598 442294 240654 442350
rect 240722 442294 240778 442350
rect 240598 442170 240654 442226
rect 240722 442170 240778 442226
rect 240598 442046 240654 442102
rect 240722 442046 240778 442102
rect 240598 441922 240654 441978
rect 240722 441922 240778 441978
rect 271318 442294 271374 442350
rect 271442 442294 271498 442350
rect 271318 442170 271374 442226
rect 271442 442170 271498 442226
rect 271318 442046 271374 442102
rect 271442 442046 271498 442102
rect 271318 441922 271374 441978
rect 271442 441922 271498 441978
rect 302038 442294 302094 442350
rect 302162 442294 302218 442350
rect 302038 442170 302094 442226
rect 302162 442170 302218 442226
rect 302038 442046 302094 442102
rect 302162 442046 302218 442102
rect 302038 441922 302094 441978
rect 302162 441922 302218 441978
rect 332758 442294 332814 442350
rect 332882 442294 332938 442350
rect 332758 442170 332814 442226
rect 332882 442170 332938 442226
rect 332758 442046 332814 442102
rect 332882 442046 332938 442102
rect 332758 441922 332814 441978
rect 332882 441922 332938 441978
rect 363478 442294 363534 442350
rect 363602 442294 363658 442350
rect 363478 442170 363534 442226
rect 363602 442170 363658 442226
rect 363478 442046 363534 442102
rect 363602 442046 363658 442102
rect 363478 441922 363534 441978
rect 363602 441922 363658 441978
rect 394198 442294 394254 442350
rect 394322 442294 394378 442350
rect 394198 442170 394254 442226
rect 394322 442170 394378 442226
rect 394198 442046 394254 442102
rect 394322 442046 394378 442102
rect 394198 441922 394254 441978
rect 394322 441922 394378 441978
rect 424918 442294 424974 442350
rect 425042 442294 425098 442350
rect 424918 442170 424974 442226
rect 425042 442170 425098 442226
rect 424918 442046 424974 442102
rect 425042 442046 425098 442102
rect 424918 441922 424974 441978
rect 425042 441922 425098 441978
rect 455638 442294 455694 442350
rect 455762 442294 455818 442350
rect 455638 442170 455694 442226
rect 455762 442170 455818 442226
rect 455638 442046 455694 442102
rect 455762 442046 455818 442102
rect 455638 441922 455694 441978
rect 455762 441922 455818 441978
rect 486358 442294 486414 442350
rect 486482 442294 486538 442350
rect 486358 442170 486414 442226
rect 486482 442170 486538 442226
rect 486358 442046 486414 442102
rect 486482 442046 486538 442102
rect 486358 441922 486414 441978
rect 486482 441922 486538 441978
rect 517078 442294 517134 442350
rect 517202 442294 517258 442350
rect 517078 442170 517134 442226
rect 517202 442170 517258 442226
rect 517078 442046 517134 442102
rect 517202 442046 517258 442102
rect 517078 441922 517134 441978
rect 517202 441922 517258 441978
rect 194518 436294 194574 436350
rect 194642 436294 194698 436350
rect 194518 436170 194574 436226
rect 194642 436170 194698 436226
rect 194518 436046 194574 436102
rect 194642 436046 194698 436102
rect 194518 435922 194574 435978
rect 194642 435922 194698 435978
rect 225238 436294 225294 436350
rect 225362 436294 225418 436350
rect 225238 436170 225294 436226
rect 225362 436170 225418 436226
rect 225238 436046 225294 436102
rect 225362 436046 225418 436102
rect 225238 435922 225294 435978
rect 225362 435922 225418 435978
rect 255958 436294 256014 436350
rect 256082 436294 256138 436350
rect 255958 436170 256014 436226
rect 256082 436170 256138 436226
rect 255958 436046 256014 436102
rect 256082 436046 256138 436102
rect 255958 435922 256014 435978
rect 256082 435922 256138 435978
rect 286678 436294 286734 436350
rect 286802 436294 286858 436350
rect 286678 436170 286734 436226
rect 286802 436170 286858 436226
rect 286678 436046 286734 436102
rect 286802 436046 286858 436102
rect 286678 435922 286734 435978
rect 286802 435922 286858 435978
rect 317398 436294 317454 436350
rect 317522 436294 317578 436350
rect 317398 436170 317454 436226
rect 317522 436170 317578 436226
rect 317398 436046 317454 436102
rect 317522 436046 317578 436102
rect 317398 435922 317454 435978
rect 317522 435922 317578 435978
rect 348118 436294 348174 436350
rect 348242 436294 348298 436350
rect 348118 436170 348174 436226
rect 348242 436170 348298 436226
rect 348118 436046 348174 436102
rect 348242 436046 348298 436102
rect 348118 435922 348174 435978
rect 348242 435922 348298 435978
rect 378838 436294 378894 436350
rect 378962 436294 379018 436350
rect 378838 436170 378894 436226
rect 378962 436170 379018 436226
rect 378838 436046 378894 436102
rect 378962 436046 379018 436102
rect 378838 435922 378894 435978
rect 378962 435922 379018 435978
rect 409558 436294 409614 436350
rect 409682 436294 409738 436350
rect 409558 436170 409614 436226
rect 409682 436170 409738 436226
rect 409558 436046 409614 436102
rect 409682 436046 409738 436102
rect 409558 435922 409614 435978
rect 409682 435922 409738 435978
rect 440278 436294 440334 436350
rect 440402 436294 440458 436350
rect 440278 436170 440334 436226
rect 440402 436170 440458 436226
rect 440278 436046 440334 436102
rect 440402 436046 440458 436102
rect 440278 435922 440334 435978
rect 440402 435922 440458 435978
rect 470998 436294 471054 436350
rect 471122 436294 471178 436350
rect 470998 436170 471054 436226
rect 471122 436170 471178 436226
rect 470998 436046 471054 436102
rect 471122 436046 471178 436102
rect 470998 435922 471054 435978
rect 471122 435922 471178 435978
rect 501718 436294 501774 436350
rect 501842 436294 501898 436350
rect 501718 436170 501774 436226
rect 501842 436170 501898 436226
rect 501718 436046 501774 436102
rect 501842 436046 501898 436102
rect 501718 435922 501774 435978
rect 501842 435922 501898 435978
rect 532438 436294 532494 436350
rect 532562 436294 532618 436350
rect 532438 436170 532494 436226
rect 532562 436170 532618 436226
rect 532438 436046 532494 436102
rect 532562 436046 532618 436102
rect 532438 435922 532494 435978
rect 532562 435922 532618 435978
rect 209878 424294 209934 424350
rect 210002 424294 210058 424350
rect 209878 424170 209934 424226
rect 210002 424170 210058 424226
rect 209878 424046 209934 424102
rect 210002 424046 210058 424102
rect 209878 423922 209934 423978
rect 210002 423922 210058 423978
rect 240598 424294 240654 424350
rect 240722 424294 240778 424350
rect 240598 424170 240654 424226
rect 240722 424170 240778 424226
rect 240598 424046 240654 424102
rect 240722 424046 240778 424102
rect 240598 423922 240654 423978
rect 240722 423922 240778 423978
rect 271318 424294 271374 424350
rect 271442 424294 271498 424350
rect 271318 424170 271374 424226
rect 271442 424170 271498 424226
rect 271318 424046 271374 424102
rect 271442 424046 271498 424102
rect 271318 423922 271374 423978
rect 271442 423922 271498 423978
rect 302038 424294 302094 424350
rect 302162 424294 302218 424350
rect 302038 424170 302094 424226
rect 302162 424170 302218 424226
rect 302038 424046 302094 424102
rect 302162 424046 302218 424102
rect 302038 423922 302094 423978
rect 302162 423922 302218 423978
rect 332758 424294 332814 424350
rect 332882 424294 332938 424350
rect 332758 424170 332814 424226
rect 332882 424170 332938 424226
rect 332758 424046 332814 424102
rect 332882 424046 332938 424102
rect 332758 423922 332814 423978
rect 332882 423922 332938 423978
rect 363478 424294 363534 424350
rect 363602 424294 363658 424350
rect 363478 424170 363534 424226
rect 363602 424170 363658 424226
rect 363478 424046 363534 424102
rect 363602 424046 363658 424102
rect 363478 423922 363534 423978
rect 363602 423922 363658 423978
rect 394198 424294 394254 424350
rect 394322 424294 394378 424350
rect 394198 424170 394254 424226
rect 394322 424170 394378 424226
rect 394198 424046 394254 424102
rect 394322 424046 394378 424102
rect 394198 423922 394254 423978
rect 394322 423922 394378 423978
rect 424918 424294 424974 424350
rect 425042 424294 425098 424350
rect 424918 424170 424974 424226
rect 425042 424170 425098 424226
rect 424918 424046 424974 424102
rect 425042 424046 425098 424102
rect 424918 423922 424974 423978
rect 425042 423922 425098 423978
rect 455638 424294 455694 424350
rect 455762 424294 455818 424350
rect 455638 424170 455694 424226
rect 455762 424170 455818 424226
rect 455638 424046 455694 424102
rect 455762 424046 455818 424102
rect 455638 423922 455694 423978
rect 455762 423922 455818 423978
rect 486358 424294 486414 424350
rect 486482 424294 486538 424350
rect 486358 424170 486414 424226
rect 486482 424170 486538 424226
rect 486358 424046 486414 424102
rect 486482 424046 486538 424102
rect 486358 423922 486414 423978
rect 486482 423922 486538 423978
rect 517078 424294 517134 424350
rect 517202 424294 517258 424350
rect 517078 424170 517134 424226
rect 517202 424170 517258 424226
rect 517078 424046 517134 424102
rect 517202 424046 517258 424102
rect 517078 423922 517134 423978
rect 517202 423922 517258 423978
rect 194518 418294 194574 418350
rect 194642 418294 194698 418350
rect 194518 418170 194574 418226
rect 194642 418170 194698 418226
rect 194518 418046 194574 418102
rect 194642 418046 194698 418102
rect 194518 417922 194574 417978
rect 194642 417922 194698 417978
rect 225238 418294 225294 418350
rect 225362 418294 225418 418350
rect 225238 418170 225294 418226
rect 225362 418170 225418 418226
rect 225238 418046 225294 418102
rect 225362 418046 225418 418102
rect 225238 417922 225294 417978
rect 225362 417922 225418 417978
rect 255958 418294 256014 418350
rect 256082 418294 256138 418350
rect 255958 418170 256014 418226
rect 256082 418170 256138 418226
rect 255958 418046 256014 418102
rect 256082 418046 256138 418102
rect 255958 417922 256014 417978
rect 256082 417922 256138 417978
rect 286678 418294 286734 418350
rect 286802 418294 286858 418350
rect 286678 418170 286734 418226
rect 286802 418170 286858 418226
rect 286678 418046 286734 418102
rect 286802 418046 286858 418102
rect 286678 417922 286734 417978
rect 286802 417922 286858 417978
rect 317398 418294 317454 418350
rect 317522 418294 317578 418350
rect 317398 418170 317454 418226
rect 317522 418170 317578 418226
rect 317398 418046 317454 418102
rect 317522 418046 317578 418102
rect 317398 417922 317454 417978
rect 317522 417922 317578 417978
rect 348118 418294 348174 418350
rect 348242 418294 348298 418350
rect 348118 418170 348174 418226
rect 348242 418170 348298 418226
rect 348118 418046 348174 418102
rect 348242 418046 348298 418102
rect 348118 417922 348174 417978
rect 348242 417922 348298 417978
rect 378838 418294 378894 418350
rect 378962 418294 379018 418350
rect 378838 418170 378894 418226
rect 378962 418170 379018 418226
rect 378838 418046 378894 418102
rect 378962 418046 379018 418102
rect 378838 417922 378894 417978
rect 378962 417922 379018 417978
rect 409558 418294 409614 418350
rect 409682 418294 409738 418350
rect 409558 418170 409614 418226
rect 409682 418170 409738 418226
rect 409558 418046 409614 418102
rect 409682 418046 409738 418102
rect 409558 417922 409614 417978
rect 409682 417922 409738 417978
rect 440278 418294 440334 418350
rect 440402 418294 440458 418350
rect 440278 418170 440334 418226
rect 440402 418170 440458 418226
rect 440278 418046 440334 418102
rect 440402 418046 440458 418102
rect 440278 417922 440334 417978
rect 440402 417922 440458 417978
rect 470998 418294 471054 418350
rect 471122 418294 471178 418350
rect 470998 418170 471054 418226
rect 471122 418170 471178 418226
rect 470998 418046 471054 418102
rect 471122 418046 471178 418102
rect 470998 417922 471054 417978
rect 471122 417922 471178 417978
rect 501718 418294 501774 418350
rect 501842 418294 501898 418350
rect 501718 418170 501774 418226
rect 501842 418170 501898 418226
rect 501718 418046 501774 418102
rect 501842 418046 501898 418102
rect 501718 417922 501774 417978
rect 501842 417922 501898 417978
rect 532438 418294 532494 418350
rect 532562 418294 532618 418350
rect 532438 418170 532494 418226
rect 532562 418170 532618 418226
rect 532438 418046 532494 418102
rect 532562 418046 532618 418102
rect 532438 417922 532494 417978
rect 532562 417922 532618 417978
rect 308028 409202 308084 409258
rect 302652 409022 302708 409078
rect 193554 406294 193610 406350
rect 193678 406294 193734 406350
rect 193802 406294 193858 406350
rect 193926 406294 193982 406350
rect 193554 406170 193610 406226
rect 193678 406170 193734 406226
rect 193802 406170 193858 406226
rect 193926 406170 193982 406226
rect 193554 406046 193610 406102
rect 193678 406046 193734 406102
rect 193802 406046 193858 406102
rect 193926 406046 193982 406102
rect 193554 405922 193610 405978
rect 193678 405922 193734 405978
rect 193802 405922 193858 405978
rect 193926 405922 193982 405978
rect 220554 400294 220610 400350
rect 220678 400294 220734 400350
rect 220802 400294 220858 400350
rect 220926 400294 220982 400350
rect 220554 400170 220610 400226
rect 220678 400170 220734 400226
rect 220802 400170 220858 400226
rect 220926 400170 220982 400226
rect 220554 400046 220610 400102
rect 220678 400046 220734 400102
rect 220802 400046 220858 400102
rect 220926 400046 220982 400102
rect 220554 399922 220610 399978
rect 220678 399922 220734 399978
rect 220802 399922 220858 399978
rect 220926 399922 220982 399978
rect 193554 388294 193610 388350
rect 193678 388294 193734 388350
rect 193802 388294 193858 388350
rect 193926 388294 193982 388350
rect 193554 388170 193610 388226
rect 193678 388170 193734 388226
rect 193802 388170 193858 388226
rect 193926 388170 193982 388226
rect 193554 388046 193610 388102
rect 193678 388046 193734 388102
rect 193802 388046 193858 388102
rect 193926 388046 193982 388102
rect 193554 387922 193610 387978
rect 193678 387922 193734 387978
rect 193802 387922 193858 387978
rect 193926 387922 193982 387978
rect 212492 388862 212548 388918
rect 193554 370294 193610 370350
rect 193678 370294 193734 370350
rect 193802 370294 193858 370350
rect 193926 370294 193982 370350
rect 193554 370170 193610 370226
rect 193678 370170 193734 370226
rect 193802 370170 193858 370226
rect 193926 370170 193982 370226
rect 193554 370046 193610 370102
rect 193678 370046 193734 370102
rect 193802 370046 193858 370102
rect 193926 370046 193982 370102
rect 193554 369922 193610 369978
rect 193678 369922 193734 369978
rect 193802 369922 193858 369978
rect 193926 369922 193982 369978
rect 193554 352294 193610 352350
rect 193678 352294 193734 352350
rect 193802 352294 193858 352350
rect 193926 352294 193982 352350
rect 193554 352170 193610 352226
rect 193678 352170 193734 352226
rect 193802 352170 193858 352226
rect 193926 352170 193982 352226
rect 193554 352046 193610 352102
rect 193678 352046 193734 352102
rect 193802 352046 193858 352102
rect 193926 352046 193982 352102
rect 193554 351922 193610 351978
rect 193678 351922 193734 351978
rect 193802 351922 193858 351978
rect 193926 351922 193982 351978
rect 193554 334294 193610 334350
rect 193678 334294 193734 334350
rect 193802 334294 193858 334350
rect 193926 334294 193982 334350
rect 193554 334170 193610 334226
rect 193678 334170 193734 334226
rect 193802 334170 193858 334226
rect 193926 334170 193982 334226
rect 193554 334046 193610 334102
rect 193678 334046 193734 334102
rect 193802 334046 193858 334102
rect 193926 334046 193982 334102
rect 193554 333922 193610 333978
rect 193678 333922 193734 333978
rect 193802 333922 193858 333978
rect 193926 333922 193982 333978
rect 193554 316294 193610 316350
rect 193678 316294 193734 316350
rect 193802 316294 193858 316350
rect 193926 316294 193982 316350
rect 193554 316170 193610 316226
rect 193678 316170 193734 316226
rect 193802 316170 193858 316226
rect 193926 316170 193982 316226
rect 193554 316046 193610 316102
rect 193678 316046 193734 316102
rect 193802 316046 193858 316102
rect 193926 316046 193982 316102
rect 193554 315922 193610 315978
rect 193678 315922 193734 315978
rect 193802 315922 193858 315978
rect 193926 315922 193982 315978
rect 193554 298294 193610 298350
rect 193678 298294 193734 298350
rect 193802 298294 193858 298350
rect 193926 298294 193982 298350
rect 193554 298170 193610 298226
rect 193678 298170 193734 298226
rect 193802 298170 193858 298226
rect 193926 298170 193982 298226
rect 193554 298046 193610 298102
rect 193678 298046 193734 298102
rect 193802 298046 193858 298102
rect 193926 298046 193982 298102
rect 193554 297922 193610 297978
rect 193678 297922 193734 297978
rect 193802 297922 193858 297978
rect 193926 297922 193982 297978
rect 189834 274294 189890 274350
rect 189958 274294 190014 274350
rect 190082 274294 190138 274350
rect 190206 274294 190262 274350
rect 189834 274170 189890 274226
rect 189958 274170 190014 274226
rect 190082 274170 190138 274226
rect 190206 274170 190262 274226
rect 189834 274046 189890 274102
rect 189958 274046 190014 274102
rect 190082 274046 190138 274102
rect 190206 274046 190262 274102
rect 189834 273922 189890 273978
rect 189958 273922 190014 273978
rect 190082 273922 190138 273978
rect 190206 273922 190262 273978
rect 189532 268802 189588 268858
rect 189834 256294 189890 256350
rect 189958 256294 190014 256350
rect 190082 256294 190138 256350
rect 190206 256294 190262 256350
rect 189834 256170 189890 256226
rect 189958 256170 190014 256226
rect 190082 256170 190138 256226
rect 190206 256170 190262 256226
rect 189834 256046 189890 256102
rect 189958 256046 190014 256102
rect 190082 256046 190138 256102
rect 190206 256046 190262 256102
rect 189834 255922 189890 255978
rect 189958 255922 190014 255978
rect 190082 255922 190138 255978
rect 190206 255922 190262 255978
rect 162834 244294 162890 244350
rect 162958 244294 163014 244350
rect 163082 244294 163138 244350
rect 163206 244294 163262 244350
rect 162834 244170 162890 244226
rect 162958 244170 163014 244226
rect 163082 244170 163138 244226
rect 163206 244170 163262 244226
rect 162834 244046 162890 244102
rect 162958 244046 163014 244102
rect 163082 244046 163138 244102
rect 163206 244046 163262 244102
rect 162834 243922 162890 243978
rect 162958 243922 163014 243978
rect 163082 243922 163138 243978
rect 163206 243922 163262 243978
rect 162834 226294 162890 226350
rect 162958 226294 163014 226350
rect 163082 226294 163138 226350
rect 163206 226294 163262 226350
rect 162834 226170 162890 226226
rect 162958 226170 163014 226226
rect 163082 226170 163138 226226
rect 163206 226170 163262 226226
rect 162834 226046 162890 226102
rect 162958 226046 163014 226102
rect 163082 226046 163138 226102
rect 163206 226046 163262 226102
rect 162834 225922 162890 225978
rect 162958 225922 163014 225978
rect 163082 225922 163138 225978
rect 163206 225922 163262 225978
rect 189834 238294 189890 238350
rect 189958 238294 190014 238350
rect 190082 238294 190138 238350
rect 190206 238294 190262 238350
rect 189834 238170 189890 238226
rect 189958 238170 190014 238226
rect 190082 238170 190138 238226
rect 190206 238170 190262 238226
rect 189834 238046 189890 238102
rect 189958 238046 190014 238102
rect 190082 238046 190138 238102
rect 190206 238046 190262 238102
rect 189834 237922 189890 237978
rect 189958 237922 190014 237978
rect 190082 237922 190138 237978
rect 190206 237922 190262 237978
rect 189834 220294 189890 220350
rect 189958 220294 190014 220350
rect 190082 220294 190138 220350
rect 190206 220294 190262 220350
rect 189834 220170 189890 220226
rect 189958 220170 190014 220226
rect 190082 220170 190138 220226
rect 190206 220170 190262 220226
rect 189834 220046 189890 220102
rect 189958 220046 190014 220102
rect 190082 220046 190138 220102
rect 190206 220046 190262 220102
rect 189834 219922 189890 219978
rect 189958 219922 190014 219978
rect 190082 219922 190138 219978
rect 190206 219922 190262 219978
rect 193554 280294 193610 280350
rect 193678 280294 193734 280350
rect 193802 280294 193858 280350
rect 193926 280294 193982 280350
rect 193554 280170 193610 280226
rect 193678 280170 193734 280226
rect 193802 280170 193858 280226
rect 193926 280170 193982 280226
rect 193554 280046 193610 280102
rect 193678 280046 193734 280102
rect 193802 280046 193858 280102
rect 193926 280046 193982 280102
rect 193554 279922 193610 279978
rect 193678 279922 193734 279978
rect 193802 279922 193858 279978
rect 193926 279922 193982 279978
rect 193554 262294 193610 262350
rect 193678 262294 193734 262350
rect 193802 262294 193858 262350
rect 193926 262294 193982 262350
rect 193554 262170 193610 262226
rect 193678 262170 193734 262226
rect 193802 262170 193858 262226
rect 193926 262170 193982 262226
rect 193554 262046 193610 262102
rect 193678 262046 193734 262102
rect 193802 262046 193858 262102
rect 193926 262046 193982 262102
rect 193554 261922 193610 261978
rect 193678 261922 193734 261978
rect 193802 261922 193858 261978
rect 193926 261922 193982 261978
rect 193554 244294 193610 244350
rect 193678 244294 193734 244350
rect 193802 244294 193858 244350
rect 193926 244294 193982 244350
rect 193554 244170 193610 244226
rect 193678 244170 193734 244226
rect 193802 244170 193858 244226
rect 193926 244170 193982 244226
rect 193554 244046 193610 244102
rect 193678 244046 193734 244102
rect 193802 244046 193858 244102
rect 193926 244046 193982 244102
rect 193554 243922 193610 243978
rect 193678 243922 193734 243978
rect 193802 243922 193858 243978
rect 193926 243922 193982 243978
rect 220554 382294 220610 382350
rect 220678 382294 220734 382350
rect 220802 382294 220858 382350
rect 220926 382294 220982 382350
rect 220554 382170 220610 382226
rect 220678 382170 220734 382226
rect 220802 382170 220858 382226
rect 220926 382170 220982 382226
rect 220554 382046 220610 382102
rect 220678 382046 220734 382102
rect 220802 382046 220858 382102
rect 220926 382046 220982 382102
rect 220554 381922 220610 381978
rect 220678 381922 220734 381978
rect 220802 381922 220858 381978
rect 220926 381922 220982 381978
rect 220554 364294 220610 364350
rect 220678 364294 220734 364350
rect 220802 364294 220858 364350
rect 220926 364294 220982 364350
rect 220554 364170 220610 364226
rect 220678 364170 220734 364226
rect 220802 364170 220858 364226
rect 220926 364170 220982 364226
rect 220554 364046 220610 364102
rect 220678 364046 220734 364102
rect 220802 364046 220858 364102
rect 220926 364046 220982 364102
rect 220554 363922 220610 363978
rect 220678 363922 220734 363978
rect 220802 363922 220858 363978
rect 220926 363922 220982 363978
rect 220554 346294 220610 346350
rect 220678 346294 220734 346350
rect 220802 346294 220858 346350
rect 220926 346294 220982 346350
rect 220554 346170 220610 346226
rect 220678 346170 220734 346226
rect 220802 346170 220858 346226
rect 220926 346170 220982 346226
rect 220554 346046 220610 346102
rect 220678 346046 220734 346102
rect 220802 346046 220858 346102
rect 220926 346046 220982 346102
rect 220554 345922 220610 345978
rect 220678 345922 220734 345978
rect 220802 345922 220858 345978
rect 220926 345922 220982 345978
rect 193554 226294 193610 226350
rect 193678 226294 193734 226350
rect 193802 226294 193858 226350
rect 193926 226294 193982 226350
rect 193554 226170 193610 226226
rect 193678 226170 193734 226226
rect 193802 226170 193858 226226
rect 193926 226170 193982 226226
rect 193554 226046 193610 226102
rect 193678 226046 193734 226102
rect 193802 226046 193858 226102
rect 193926 226046 193982 226102
rect 193554 225922 193610 225978
rect 193678 225922 193734 225978
rect 193802 225922 193858 225978
rect 193926 225922 193982 225978
rect 245196 407596 245252 407638
rect 245196 407582 245252 407596
rect 238140 407402 238196 407458
rect 224274 406294 224330 406350
rect 224398 406294 224454 406350
rect 224522 406294 224578 406350
rect 224646 406294 224702 406350
rect 224274 406170 224330 406226
rect 224398 406170 224454 406226
rect 224522 406170 224578 406226
rect 224646 406170 224702 406226
rect 224274 406046 224330 406102
rect 224398 406046 224454 406102
rect 224522 406046 224578 406102
rect 224646 406046 224702 406102
rect 224274 405922 224330 405978
rect 224398 405922 224454 405978
rect 224522 405922 224578 405978
rect 224646 405922 224702 405978
rect 224274 388294 224330 388350
rect 224398 388294 224454 388350
rect 224522 388294 224578 388350
rect 224646 388294 224702 388350
rect 224274 388170 224330 388226
rect 224398 388170 224454 388226
rect 224522 388170 224578 388226
rect 224646 388170 224702 388226
rect 224274 388046 224330 388102
rect 224398 388046 224454 388102
rect 224522 388046 224578 388102
rect 224646 388046 224702 388102
rect 224274 387922 224330 387978
rect 224398 387922 224454 387978
rect 224522 387922 224578 387978
rect 224646 387922 224702 387978
rect 224274 370294 224330 370350
rect 224398 370294 224454 370350
rect 224522 370294 224578 370350
rect 224646 370294 224702 370350
rect 224274 370170 224330 370226
rect 224398 370170 224454 370226
rect 224522 370170 224578 370226
rect 224646 370170 224702 370226
rect 224274 370046 224330 370102
rect 224398 370046 224454 370102
rect 224522 370046 224578 370102
rect 224646 370046 224702 370102
rect 224274 369922 224330 369978
rect 224398 369922 224454 369978
rect 224522 369922 224578 369978
rect 224646 369922 224702 369978
rect 224274 352294 224330 352350
rect 224398 352294 224454 352350
rect 224522 352294 224578 352350
rect 224646 352294 224702 352350
rect 224274 352170 224330 352226
rect 224398 352170 224454 352226
rect 224522 352170 224578 352226
rect 224646 352170 224702 352226
rect 224274 352046 224330 352102
rect 224398 352046 224454 352102
rect 224522 352046 224578 352102
rect 224646 352046 224702 352102
rect 224274 351922 224330 351978
rect 224398 351922 224454 351978
rect 224522 351922 224578 351978
rect 224646 351922 224702 351978
rect 224274 334294 224330 334350
rect 224398 334294 224454 334350
rect 224522 334294 224578 334350
rect 224646 334294 224702 334350
rect 224274 334170 224330 334226
rect 224398 334170 224454 334226
rect 224522 334170 224578 334226
rect 224646 334170 224702 334226
rect 224274 334046 224330 334102
rect 224398 334046 224454 334102
rect 224522 334046 224578 334102
rect 224646 334046 224702 334102
rect 224274 333922 224330 333978
rect 224398 333922 224454 333978
rect 224522 333922 224578 333978
rect 224646 333922 224702 333978
rect 220554 328294 220610 328350
rect 220678 328294 220734 328350
rect 220802 328294 220858 328350
rect 220926 328294 220982 328350
rect 220554 328170 220610 328226
rect 220678 328170 220734 328226
rect 220802 328170 220858 328226
rect 220926 328170 220982 328226
rect 220554 328046 220610 328102
rect 220678 328046 220734 328102
rect 220802 328046 220858 328102
rect 220926 328046 220982 328102
rect 220554 327922 220610 327978
rect 220678 327922 220734 327978
rect 220802 327922 220858 327978
rect 220926 327922 220982 327978
rect 220554 310294 220610 310350
rect 220678 310294 220734 310350
rect 220802 310294 220858 310350
rect 220926 310294 220982 310350
rect 220554 310170 220610 310226
rect 220678 310170 220734 310226
rect 220802 310170 220858 310226
rect 220926 310170 220982 310226
rect 220554 310046 220610 310102
rect 220678 310046 220734 310102
rect 220802 310046 220858 310102
rect 220926 310046 220982 310102
rect 220554 309922 220610 309978
rect 220678 309922 220734 309978
rect 220802 309922 220858 309978
rect 220926 309922 220982 309978
rect 220554 292294 220610 292350
rect 220678 292294 220734 292350
rect 220802 292294 220858 292350
rect 220926 292294 220982 292350
rect 220554 292170 220610 292226
rect 220678 292170 220734 292226
rect 220802 292170 220858 292226
rect 220926 292170 220982 292226
rect 220554 292046 220610 292102
rect 220678 292046 220734 292102
rect 220802 292046 220858 292102
rect 220926 292046 220982 292102
rect 220554 291922 220610 291978
rect 220678 291922 220734 291978
rect 220802 291922 220858 291978
rect 220926 291922 220982 291978
rect 220554 274294 220610 274350
rect 220678 274294 220734 274350
rect 220802 274294 220858 274350
rect 220926 274294 220982 274350
rect 220554 274170 220610 274226
rect 220678 274170 220734 274226
rect 220802 274170 220858 274226
rect 220926 274170 220982 274226
rect 220554 274046 220610 274102
rect 220678 274046 220734 274102
rect 220802 274046 220858 274102
rect 220926 274046 220982 274102
rect 220554 273922 220610 273978
rect 220678 273922 220734 273978
rect 220802 273922 220858 273978
rect 220926 273922 220982 273978
rect 220554 256294 220610 256350
rect 220678 256294 220734 256350
rect 220802 256294 220858 256350
rect 220926 256294 220982 256350
rect 220554 256170 220610 256226
rect 220678 256170 220734 256226
rect 220802 256170 220858 256226
rect 220926 256170 220982 256226
rect 220554 256046 220610 256102
rect 220678 256046 220734 256102
rect 220802 256046 220858 256102
rect 220926 256046 220982 256102
rect 220554 255922 220610 255978
rect 220678 255922 220734 255978
rect 220802 255922 220858 255978
rect 220926 255922 220982 255978
rect 220554 238294 220610 238350
rect 220678 238294 220734 238350
rect 220802 238294 220858 238350
rect 220926 238294 220982 238350
rect 220554 238170 220610 238226
rect 220678 238170 220734 238226
rect 220802 238170 220858 238226
rect 220926 238170 220982 238226
rect 220554 238046 220610 238102
rect 220678 238046 220734 238102
rect 220802 238046 220858 238102
rect 220926 238046 220982 238102
rect 220554 237922 220610 237978
rect 220678 237922 220734 237978
rect 220802 237922 220858 237978
rect 220926 237922 220982 237978
rect 224274 316294 224330 316350
rect 224398 316294 224454 316350
rect 224522 316294 224578 316350
rect 224646 316294 224702 316350
rect 224274 316170 224330 316226
rect 224398 316170 224454 316226
rect 224522 316170 224578 316226
rect 224646 316170 224702 316226
rect 224274 316046 224330 316102
rect 224398 316046 224454 316102
rect 224522 316046 224578 316102
rect 224646 316046 224702 316102
rect 224274 315922 224330 315978
rect 224398 315922 224454 315978
rect 224522 315922 224578 315978
rect 224646 315922 224702 315978
rect 224274 298294 224330 298350
rect 224398 298294 224454 298350
rect 224522 298294 224578 298350
rect 224646 298294 224702 298350
rect 224274 298170 224330 298226
rect 224398 298170 224454 298226
rect 224522 298170 224578 298226
rect 224646 298170 224702 298226
rect 224274 298046 224330 298102
rect 224398 298046 224454 298102
rect 224522 298046 224578 298102
rect 224646 298046 224702 298102
rect 224274 297922 224330 297978
rect 224398 297922 224454 297978
rect 224522 297922 224578 297978
rect 224646 297922 224702 297978
rect 224274 280294 224330 280350
rect 224398 280294 224454 280350
rect 224522 280294 224578 280350
rect 224646 280294 224702 280350
rect 224274 280170 224330 280226
rect 224398 280170 224454 280226
rect 224522 280170 224578 280226
rect 224646 280170 224702 280226
rect 224274 280046 224330 280102
rect 224398 280046 224454 280102
rect 224522 280046 224578 280102
rect 224646 280046 224702 280102
rect 224274 279922 224330 279978
rect 224398 279922 224454 279978
rect 224522 279922 224578 279978
rect 224646 279922 224702 279978
rect 224274 262294 224330 262350
rect 224398 262294 224454 262350
rect 224522 262294 224578 262350
rect 224646 262294 224702 262350
rect 224274 262170 224330 262226
rect 224398 262170 224454 262226
rect 224522 262170 224578 262226
rect 224646 262170 224702 262226
rect 224274 262046 224330 262102
rect 224398 262046 224454 262102
rect 224522 262046 224578 262102
rect 224646 262046 224702 262102
rect 224274 261922 224330 261978
rect 224398 261922 224454 261978
rect 224522 261922 224578 261978
rect 224646 261922 224702 261978
rect 224274 244294 224330 244350
rect 224398 244294 224454 244350
rect 224522 244294 224578 244350
rect 224646 244294 224702 244350
rect 224274 244170 224330 244226
rect 224398 244170 224454 244226
rect 224522 244170 224578 244226
rect 224646 244170 224702 244226
rect 224274 244046 224330 244102
rect 224398 244046 224454 244102
rect 224522 244046 224578 244102
rect 224646 244046 224702 244102
rect 224274 243922 224330 243978
rect 224398 243922 224454 243978
rect 224522 243922 224578 243978
rect 224646 243922 224702 243978
rect 220554 220294 220610 220350
rect 220678 220294 220734 220350
rect 220802 220294 220858 220350
rect 220926 220294 220982 220350
rect 220554 220170 220610 220226
rect 220678 220170 220734 220226
rect 220802 220170 220858 220226
rect 220926 220170 220982 220226
rect 220554 220046 220610 220102
rect 220678 220046 220734 220102
rect 220802 220046 220858 220102
rect 220926 220046 220982 220102
rect 220554 219922 220610 219978
rect 220678 219922 220734 219978
rect 220802 219922 220858 219978
rect 220926 219922 220982 219978
rect 224274 226294 224330 226350
rect 224398 226294 224454 226350
rect 224522 226294 224578 226350
rect 224646 226294 224702 226350
rect 224274 226170 224330 226226
rect 224398 226170 224454 226226
rect 224522 226170 224578 226226
rect 224646 226170 224702 226226
rect 224274 226046 224330 226102
rect 224398 226046 224454 226102
rect 224522 226046 224578 226102
rect 224646 226046 224702 226102
rect 224274 225922 224330 225978
rect 224398 225922 224454 225978
rect 224522 225922 224578 225978
rect 224646 225922 224702 225978
rect 231756 403982 231812 404038
rect 230972 249362 231028 249418
rect 231868 246122 231924 246178
rect 235900 382562 235956 382618
rect 237692 385622 237748 385678
rect 237580 268802 237636 268858
rect 236236 211022 236292 211078
rect 238252 389762 238308 389818
rect 254994 406294 255050 406350
rect 255118 406294 255174 406350
rect 255242 406294 255298 406350
rect 255366 406294 255422 406350
rect 254994 406170 255050 406226
rect 255118 406170 255174 406226
rect 255242 406170 255298 406226
rect 255366 406170 255422 406226
rect 254994 406046 255050 406102
rect 255118 406046 255174 406102
rect 255242 406046 255298 406102
rect 255366 406046 255422 406102
rect 254994 405922 255050 405978
rect 255118 405922 255174 405978
rect 255242 405922 255298 405978
rect 255366 405922 255422 405978
rect 285714 406294 285770 406350
rect 285838 406294 285894 406350
rect 285962 406294 286018 406350
rect 286086 406294 286142 406350
rect 285714 406170 285770 406226
rect 285838 406170 285894 406226
rect 285962 406170 286018 406226
rect 286086 406170 286142 406226
rect 285714 406046 285770 406102
rect 285838 406046 285894 406102
rect 285962 406046 286018 406102
rect 286086 406046 286142 406102
rect 285714 405922 285770 405978
rect 285838 405922 285894 405978
rect 285962 405922 286018 405978
rect 286086 405922 286142 405978
rect 254994 388294 255050 388350
rect 255118 388294 255174 388350
rect 255242 388294 255298 388350
rect 255366 388294 255422 388350
rect 254994 388170 255050 388226
rect 255118 388170 255174 388226
rect 255242 388170 255298 388226
rect 255366 388170 255422 388226
rect 254994 388046 255050 388102
rect 255118 388046 255174 388102
rect 255242 388046 255298 388102
rect 255366 388046 255422 388102
rect 282156 388682 282212 388738
rect 285714 388294 285770 388350
rect 285838 388294 285894 388350
rect 285962 388294 286018 388350
rect 286086 388294 286142 388350
rect 285714 388170 285770 388226
rect 285838 388170 285894 388226
rect 285962 388170 286018 388226
rect 286086 388170 286142 388226
rect 254994 387922 255050 387978
rect 255118 387922 255174 387978
rect 255242 387922 255298 387978
rect 255366 387922 255422 387978
rect 285714 388046 285770 388102
rect 285838 388046 285894 388102
rect 285962 388046 286018 388102
rect 286086 388046 286142 388102
rect 285714 387922 285770 387978
rect 285838 387922 285894 387978
rect 285962 387922 286018 387978
rect 286086 387922 286142 387978
rect 267820 385476 267876 385498
rect 267820 385442 267876 385476
rect 273196 385476 273252 385498
rect 273196 385442 273252 385476
rect 269612 385308 269668 385318
rect 269612 385262 269668 385308
rect 271404 385308 271460 385318
rect 271404 385262 271460 385308
rect 297388 388862 297444 388918
rect 286300 385622 286356 385678
rect 303996 385622 304052 385678
rect 316434 406294 316490 406350
rect 316558 406294 316614 406350
rect 316682 406294 316738 406350
rect 316806 406294 316862 406350
rect 316434 406170 316490 406226
rect 316558 406170 316614 406226
rect 316682 406170 316738 406226
rect 316806 406170 316862 406226
rect 316434 406046 316490 406102
rect 316558 406046 316614 406102
rect 316682 406046 316738 406102
rect 316806 406046 316862 406102
rect 316434 405922 316490 405978
rect 316558 405922 316614 405978
rect 316682 405922 316738 405978
rect 316806 405922 316862 405978
rect 316434 388294 316490 388350
rect 316558 388294 316614 388350
rect 316682 388294 316738 388350
rect 316806 388294 316862 388350
rect 316434 388170 316490 388226
rect 316558 388170 316614 388226
rect 316682 388170 316738 388226
rect 316806 388170 316862 388226
rect 316434 388046 316490 388102
rect 316558 388046 316614 388102
rect 316682 388046 316738 388102
rect 316806 388046 316862 388102
rect 316434 387922 316490 387978
rect 316558 387922 316614 387978
rect 316682 387922 316738 387978
rect 316806 387922 316862 387978
rect 287532 384362 287588 384418
rect 288428 384182 288484 384238
rect 290220 384002 290276 384058
rect 289324 383822 289380 383878
rect 347154 406294 347210 406350
rect 347278 406294 347334 406350
rect 347402 406294 347458 406350
rect 347526 406294 347582 406350
rect 347154 406170 347210 406226
rect 347278 406170 347334 406226
rect 347402 406170 347458 406226
rect 347526 406170 347582 406226
rect 347154 406046 347210 406102
rect 347278 406046 347334 406102
rect 347402 406046 347458 406102
rect 347526 406046 347582 406102
rect 347154 405922 347210 405978
rect 347278 405922 347334 405978
rect 347402 405922 347458 405978
rect 347526 405922 347582 405978
rect 347154 388294 347210 388350
rect 347278 388294 347334 388350
rect 347402 388294 347458 388350
rect 347526 388294 347582 388350
rect 347154 388170 347210 388226
rect 347278 388170 347334 388226
rect 347402 388170 347458 388226
rect 347526 388170 347582 388226
rect 347154 388046 347210 388102
rect 347278 388046 347334 388102
rect 347402 388046 347458 388102
rect 347526 388046 347582 388102
rect 347154 387922 347210 387978
rect 347278 387922 347334 387978
rect 347402 387922 347458 387978
rect 347526 387922 347582 387978
rect 240518 382213 240574 382269
rect 240642 382213 240698 382269
rect 240518 382089 240574 382145
rect 240642 382089 240698 382145
rect 240518 381965 240574 382021
rect 240642 381965 240698 382021
rect 240518 381841 240574 381897
rect 240642 381841 240698 381897
rect 271238 382213 271294 382269
rect 271362 382213 271418 382269
rect 271238 382089 271294 382145
rect 271362 382089 271418 382145
rect 271238 381965 271294 382021
rect 271362 381965 271418 382021
rect 271238 381841 271294 381897
rect 271362 381841 271418 381897
rect 301958 382213 302014 382269
rect 302082 382213 302138 382269
rect 301958 382089 302014 382145
rect 302082 382089 302138 382145
rect 301958 381965 302014 382021
rect 302082 381965 302138 382021
rect 301958 381841 302014 381897
rect 302082 381841 302138 381897
rect 332678 382213 332734 382269
rect 332802 382213 332858 382269
rect 332678 382089 332734 382145
rect 332802 382089 332858 382145
rect 332678 381965 332734 382021
rect 332802 381965 332858 382021
rect 332678 381841 332734 381897
rect 332802 381841 332858 381897
rect 363398 382213 363454 382269
rect 363522 382213 363578 382269
rect 363398 382089 363454 382145
rect 363522 382089 363578 382145
rect 363398 381965 363454 382021
rect 363522 381965 363578 382021
rect 363398 381841 363454 381897
rect 363522 381841 363578 381897
rect 255878 370294 255934 370350
rect 256002 370294 256058 370350
rect 255878 370170 255934 370226
rect 256002 370170 256058 370226
rect 255878 370046 255934 370102
rect 256002 370046 256058 370102
rect 255878 369922 255934 369978
rect 256002 369922 256058 369978
rect 286598 370294 286654 370350
rect 286722 370294 286778 370350
rect 286598 370170 286654 370226
rect 286722 370170 286778 370226
rect 286598 370046 286654 370102
rect 286722 370046 286778 370102
rect 286598 369922 286654 369978
rect 286722 369922 286778 369978
rect 317318 370294 317374 370350
rect 317442 370294 317498 370350
rect 317318 370170 317374 370226
rect 317442 370170 317498 370226
rect 317318 370046 317374 370102
rect 317442 370046 317498 370102
rect 317318 369922 317374 369978
rect 317442 369922 317498 369978
rect 348038 370294 348094 370350
rect 348162 370294 348218 370350
rect 348038 370170 348094 370226
rect 348162 370170 348218 370226
rect 348038 370046 348094 370102
rect 348162 370046 348218 370102
rect 348038 369922 348094 369978
rect 348162 369922 348218 369978
rect 240518 364294 240574 364350
rect 240642 364294 240698 364350
rect 240518 364170 240574 364226
rect 240642 364170 240698 364226
rect 240518 364046 240574 364102
rect 240642 364046 240698 364102
rect 240518 363922 240574 363978
rect 240642 363922 240698 363978
rect 271238 364294 271294 364350
rect 271362 364294 271418 364350
rect 271238 364170 271294 364226
rect 271362 364170 271418 364226
rect 271238 364046 271294 364102
rect 271362 364046 271418 364102
rect 271238 363922 271294 363978
rect 271362 363922 271418 363978
rect 301958 364294 302014 364350
rect 302082 364294 302138 364350
rect 301958 364170 302014 364226
rect 302082 364170 302138 364226
rect 301958 364046 302014 364102
rect 302082 364046 302138 364102
rect 301958 363922 302014 363978
rect 302082 363922 302138 363978
rect 332678 364294 332734 364350
rect 332802 364294 332858 364350
rect 332678 364170 332734 364226
rect 332802 364170 332858 364226
rect 332678 364046 332734 364102
rect 332802 364046 332858 364102
rect 332678 363922 332734 363978
rect 332802 363922 332858 363978
rect 363398 364294 363454 364350
rect 363522 364294 363578 364350
rect 363398 364170 363454 364226
rect 363522 364170 363578 364226
rect 363398 364046 363454 364102
rect 363522 364046 363578 364102
rect 363398 363922 363454 363978
rect 363522 363922 363578 363978
rect 255878 352294 255934 352350
rect 256002 352294 256058 352350
rect 255878 352170 255934 352226
rect 256002 352170 256058 352226
rect 255878 352046 255934 352102
rect 256002 352046 256058 352102
rect 255878 351922 255934 351978
rect 256002 351922 256058 351978
rect 286598 352294 286654 352350
rect 286722 352294 286778 352350
rect 286598 352170 286654 352226
rect 286722 352170 286778 352226
rect 286598 352046 286654 352102
rect 286722 352046 286778 352102
rect 286598 351922 286654 351978
rect 286722 351922 286778 351978
rect 317318 352294 317374 352350
rect 317442 352294 317498 352350
rect 317318 352170 317374 352226
rect 317442 352170 317498 352226
rect 317318 352046 317374 352102
rect 317442 352046 317498 352102
rect 317318 351922 317374 351978
rect 317442 351922 317498 351978
rect 348038 352294 348094 352350
rect 348162 352294 348218 352350
rect 348038 352170 348094 352226
rect 348162 352170 348218 352226
rect 348038 352046 348094 352102
rect 348162 352046 348218 352102
rect 348038 351922 348094 351978
rect 348162 351922 348218 351978
rect 240518 346294 240574 346350
rect 240642 346294 240698 346350
rect 240518 346170 240574 346226
rect 240642 346170 240698 346226
rect 240518 346046 240574 346102
rect 240642 346046 240698 346102
rect 240518 345922 240574 345978
rect 240642 345922 240698 345978
rect 271238 346294 271294 346350
rect 271362 346294 271418 346350
rect 271238 346170 271294 346226
rect 271362 346170 271418 346226
rect 271238 346046 271294 346102
rect 271362 346046 271418 346102
rect 271238 345922 271294 345978
rect 271362 345922 271418 345978
rect 301958 346294 302014 346350
rect 302082 346294 302138 346350
rect 301958 346170 302014 346226
rect 302082 346170 302138 346226
rect 301958 346046 302014 346102
rect 302082 346046 302138 346102
rect 301958 345922 302014 345978
rect 302082 345922 302138 345978
rect 332678 346294 332734 346350
rect 332802 346294 332858 346350
rect 332678 346170 332734 346226
rect 332802 346170 332858 346226
rect 332678 346046 332734 346102
rect 332802 346046 332858 346102
rect 332678 345922 332734 345978
rect 332802 345922 332858 345978
rect 363398 346294 363454 346350
rect 363522 346294 363578 346350
rect 363398 346170 363454 346226
rect 363522 346170 363578 346226
rect 363398 346046 363454 346102
rect 363522 346046 363578 346102
rect 363398 345922 363454 345978
rect 363522 345922 363578 345978
rect 255878 334294 255934 334350
rect 256002 334294 256058 334350
rect 255878 334170 255934 334226
rect 256002 334170 256058 334226
rect 255878 334046 255934 334102
rect 256002 334046 256058 334102
rect 255878 333922 255934 333978
rect 256002 333922 256058 333978
rect 286598 334294 286654 334350
rect 286722 334294 286778 334350
rect 286598 334170 286654 334226
rect 286722 334170 286778 334226
rect 286598 334046 286654 334102
rect 286722 334046 286778 334102
rect 286598 333922 286654 333978
rect 286722 333922 286778 333978
rect 317318 334294 317374 334350
rect 317442 334294 317498 334350
rect 317318 334170 317374 334226
rect 317442 334170 317498 334226
rect 317318 334046 317374 334102
rect 317442 334046 317498 334102
rect 317318 333922 317374 333978
rect 317442 333922 317498 333978
rect 348038 334294 348094 334350
rect 348162 334294 348218 334350
rect 348038 334170 348094 334226
rect 348162 334170 348218 334226
rect 348038 334046 348094 334102
rect 348162 334046 348218 334102
rect 348038 333922 348094 333978
rect 348162 333922 348218 333978
rect 240518 328294 240574 328350
rect 240642 328294 240698 328350
rect 240518 328170 240574 328226
rect 240642 328170 240698 328226
rect 240518 328046 240574 328102
rect 240642 328046 240698 328102
rect 240518 327922 240574 327978
rect 240642 327922 240698 327978
rect 271238 328294 271294 328350
rect 271362 328294 271418 328350
rect 271238 328170 271294 328226
rect 271362 328170 271418 328226
rect 271238 328046 271294 328102
rect 271362 328046 271418 328102
rect 271238 327922 271294 327978
rect 271362 327922 271418 327978
rect 301958 328294 302014 328350
rect 302082 328294 302138 328350
rect 301958 328170 302014 328226
rect 302082 328170 302138 328226
rect 301958 328046 302014 328102
rect 302082 328046 302138 328102
rect 301958 327922 302014 327978
rect 302082 327922 302138 327978
rect 332678 328294 332734 328350
rect 332802 328294 332858 328350
rect 332678 328170 332734 328226
rect 332802 328170 332858 328226
rect 332678 328046 332734 328102
rect 332802 328046 332858 328102
rect 332678 327922 332734 327978
rect 332802 327922 332858 327978
rect 363398 328294 363454 328350
rect 363522 328294 363578 328350
rect 363398 328170 363454 328226
rect 363522 328170 363578 328226
rect 363398 328046 363454 328102
rect 363522 328046 363578 328102
rect 363398 327922 363454 327978
rect 363522 327922 363578 327978
rect 255878 316294 255934 316350
rect 256002 316294 256058 316350
rect 255878 316170 255934 316226
rect 256002 316170 256058 316226
rect 255878 316046 255934 316102
rect 256002 316046 256058 316102
rect 255878 315922 255934 315978
rect 256002 315922 256058 315978
rect 286598 316294 286654 316350
rect 286722 316294 286778 316350
rect 286598 316170 286654 316226
rect 286722 316170 286778 316226
rect 286598 316046 286654 316102
rect 286722 316046 286778 316102
rect 286598 315922 286654 315978
rect 286722 315922 286778 315978
rect 317318 316294 317374 316350
rect 317442 316294 317498 316350
rect 317318 316170 317374 316226
rect 317442 316170 317498 316226
rect 317318 316046 317374 316102
rect 317442 316046 317498 316102
rect 317318 315922 317374 315978
rect 317442 315922 317498 315978
rect 348038 316294 348094 316350
rect 348162 316294 348218 316350
rect 348038 316170 348094 316226
rect 348162 316170 348218 316226
rect 348038 316046 348094 316102
rect 348162 316046 348218 316102
rect 348038 315922 348094 315978
rect 348162 315922 348218 315978
rect 240518 310294 240574 310350
rect 240642 310294 240698 310350
rect 240518 310170 240574 310226
rect 240642 310170 240698 310226
rect 240518 310046 240574 310102
rect 240642 310046 240698 310102
rect 240518 309922 240574 309978
rect 240642 309922 240698 309978
rect 271238 310294 271294 310350
rect 271362 310294 271418 310350
rect 271238 310170 271294 310226
rect 271362 310170 271418 310226
rect 271238 310046 271294 310102
rect 271362 310046 271418 310102
rect 271238 309922 271294 309978
rect 271362 309922 271418 309978
rect 301958 310294 302014 310350
rect 302082 310294 302138 310350
rect 301958 310170 302014 310226
rect 302082 310170 302138 310226
rect 301958 310046 302014 310102
rect 302082 310046 302138 310102
rect 301958 309922 302014 309978
rect 302082 309922 302138 309978
rect 332678 310294 332734 310350
rect 332802 310294 332858 310350
rect 332678 310170 332734 310226
rect 332802 310170 332858 310226
rect 332678 310046 332734 310102
rect 332802 310046 332858 310102
rect 332678 309922 332734 309978
rect 332802 309922 332858 309978
rect 363398 310294 363454 310350
rect 363522 310294 363578 310350
rect 363398 310170 363454 310226
rect 363522 310170 363578 310226
rect 363398 310046 363454 310102
rect 363522 310046 363578 310102
rect 363398 309922 363454 309978
rect 363522 309922 363578 309978
rect 255878 298294 255934 298350
rect 256002 298294 256058 298350
rect 255878 298170 255934 298226
rect 256002 298170 256058 298226
rect 255878 298046 255934 298102
rect 256002 298046 256058 298102
rect 255878 297922 255934 297978
rect 256002 297922 256058 297978
rect 286598 298294 286654 298350
rect 286722 298294 286778 298350
rect 286598 298170 286654 298226
rect 286722 298170 286778 298226
rect 286598 298046 286654 298102
rect 286722 298046 286778 298102
rect 286598 297922 286654 297978
rect 286722 297922 286778 297978
rect 317318 298294 317374 298350
rect 317442 298294 317498 298350
rect 317318 298170 317374 298226
rect 317442 298170 317498 298226
rect 317318 298046 317374 298102
rect 317442 298046 317498 298102
rect 317318 297922 317374 297978
rect 317442 297922 317498 297978
rect 348038 298294 348094 298350
rect 348162 298294 348218 298350
rect 348038 298170 348094 298226
rect 348162 298170 348218 298226
rect 348038 298046 348094 298102
rect 348162 298046 348218 298102
rect 348038 297922 348094 297978
rect 348162 297922 348218 297978
rect 240518 292294 240574 292350
rect 240642 292294 240698 292350
rect 240518 292170 240574 292226
rect 240642 292170 240698 292226
rect 240518 292046 240574 292102
rect 240642 292046 240698 292102
rect 240518 291922 240574 291978
rect 240642 291922 240698 291978
rect 271238 292294 271294 292350
rect 271362 292294 271418 292350
rect 271238 292170 271294 292226
rect 271362 292170 271418 292226
rect 271238 292046 271294 292102
rect 271362 292046 271418 292102
rect 271238 291922 271294 291978
rect 271362 291922 271418 291978
rect 301958 292294 302014 292350
rect 302082 292294 302138 292350
rect 301958 292170 302014 292226
rect 302082 292170 302138 292226
rect 301958 292046 302014 292102
rect 302082 292046 302138 292102
rect 301958 291922 302014 291978
rect 302082 291922 302138 291978
rect 332678 292294 332734 292350
rect 332802 292294 332858 292350
rect 332678 292170 332734 292226
rect 332802 292170 332858 292226
rect 332678 292046 332734 292102
rect 332802 292046 332858 292102
rect 332678 291922 332734 291978
rect 332802 291922 332858 291978
rect 363398 292294 363454 292350
rect 363522 292294 363578 292350
rect 363398 292170 363454 292226
rect 363522 292170 363578 292226
rect 363398 292046 363454 292102
rect 363522 292046 363578 292102
rect 363398 291922 363454 291978
rect 363522 291922 363578 291978
rect 255878 280294 255934 280350
rect 256002 280294 256058 280350
rect 255878 280170 255934 280226
rect 256002 280170 256058 280226
rect 255878 280046 255934 280102
rect 256002 280046 256058 280102
rect 255878 279922 255934 279978
rect 256002 279922 256058 279978
rect 286598 280294 286654 280350
rect 286722 280294 286778 280350
rect 286598 280170 286654 280226
rect 286722 280170 286778 280226
rect 286598 280046 286654 280102
rect 286722 280046 286778 280102
rect 286598 279922 286654 279978
rect 286722 279922 286778 279978
rect 317318 280294 317374 280350
rect 317442 280294 317498 280350
rect 317318 280170 317374 280226
rect 317442 280170 317498 280226
rect 317318 280046 317374 280102
rect 317442 280046 317498 280102
rect 317318 279922 317374 279978
rect 317442 279922 317498 279978
rect 348038 280294 348094 280350
rect 348162 280294 348218 280350
rect 348038 280170 348094 280226
rect 348162 280170 348218 280226
rect 348038 280046 348094 280102
rect 348162 280046 348218 280102
rect 348038 279922 348094 279978
rect 348162 279922 348218 279978
rect 240518 274294 240574 274350
rect 240642 274294 240698 274350
rect 240518 274170 240574 274226
rect 240642 274170 240698 274226
rect 240518 274046 240574 274102
rect 240642 274046 240698 274102
rect 240518 273922 240574 273978
rect 240642 273922 240698 273978
rect 271238 274294 271294 274350
rect 271362 274294 271418 274350
rect 271238 274170 271294 274226
rect 271362 274170 271418 274226
rect 271238 274046 271294 274102
rect 271362 274046 271418 274102
rect 271238 273922 271294 273978
rect 271362 273922 271418 273978
rect 301958 274294 302014 274350
rect 302082 274294 302138 274350
rect 301958 274170 302014 274226
rect 302082 274170 302138 274226
rect 301958 274046 302014 274102
rect 302082 274046 302138 274102
rect 301958 273922 302014 273978
rect 302082 273922 302138 273978
rect 332678 274294 332734 274350
rect 332802 274294 332858 274350
rect 332678 274170 332734 274226
rect 332802 274170 332858 274226
rect 332678 274046 332734 274102
rect 332802 274046 332858 274102
rect 332678 273922 332734 273978
rect 332802 273922 332858 273978
rect 363398 274294 363454 274350
rect 363522 274294 363578 274350
rect 363398 274170 363454 274226
rect 363522 274170 363578 274226
rect 363398 274046 363454 274102
rect 363522 274046 363578 274102
rect 363398 273922 363454 273978
rect 363522 273922 363578 273978
rect 255878 262294 255934 262350
rect 256002 262294 256058 262350
rect 255878 262170 255934 262226
rect 256002 262170 256058 262226
rect 255878 262046 255934 262102
rect 256002 262046 256058 262102
rect 255878 261922 255934 261978
rect 256002 261922 256058 261978
rect 286598 262294 286654 262350
rect 286722 262294 286778 262350
rect 286598 262170 286654 262226
rect 286722 262170 286778 262226
rect 286598 262046 286654 262102
rect 286722 262046 286778 262102
rect 286598 261922 286654 261978
rect 286722 261922 286778 261978
rect 317318 262294 317374 262350
rect 317442 262294 317498 262350
rect 317318 262170 317374 262226
rect 317442 262170 317498 262226
rect 317318 262046 317374 262102
rect 317442 262046 317498 262102
rect 317318 261922 317374 261978
rect 317442 261922 317498 261978
rect 348038 262294 348094 262350
rect 348162 262294 348218 262350
rect 348038 262170 348094 262226
rect 348162 262170 348218 262226
rect 348038 262046 348094 262102
rect 348162 262046 348218 262102
rect 348038 261922 348094 261978
rect 348162 261922 348218 261978
rect 358652 257822 358708 257878
rect 237916 210842 237972 210898
rect 251274 256294 251330 256350
rect 251398 256294 251454 256350
rect 251522 256294 251578 256350
rect 251646 256294 251702 256350
rect 251274 256170 251330 256226
rect 251398 256170 251454 256226
rect 251522 256170 251578 256226
rect 251646 256170 251702 256226
rect 251274 256046 251330 256102
rect 251398 256046 251454 256102
rect 251522 256046 251578 256102
rect 251646 256046 251702 256102
rect 251274 255922 251330 255978
rect 251398 255922 251454 255978
rect 251522 255922 251578 255978
rect 251646 255922 251702 255978
rect 251916 252782 251972 252838
rect 252588 252422 252644 252478
rect 251274 238294 251330 238350
rect 251398 238294 251454 238350
rect 251522 238294 251578 238350
rect 251646 238294 251702 238350
rect 251274 238170 251330 238226
rect 251398 238170 251454 238226
rect 251522 238170 251578 238226
rect 251646 238170 251702 238226
rect 251274 238046 251330 238102
rect 251398 238046 251454 238102
rect 251522 238046 251578 238102
rect 251646 238046 251702 238102
rect 251274 237922 251330 237978
rect 251398 237922 251454 237978
rect 251522 237922 251578 237978
rect 251646 237922 251702 237978
rect 251274 220294 251330 220350
rect 251398 220294 251454 220350
rect 251522 220294 251578 220350
rect 251646 220294 251702 220350
rect 251274 220170 251330 220226
rect 251398 220170 251454 220226
rect 251522 220170 251578 220226
rect 251646 220170 251702 220226
rect 251274 220046 251330 220102
rect 251398 220046 251454 220102
rect 251522 220046 251578 220102
rect 251646 220046 251702 220102
rect 251274 219922 251330 219978
rect 251398 219922 251454 219978
rect 251522 219922 251578 219978
rect 251646 219922 251702 219978
rect 258860 252602 258916 252658
rect 259756 252242 259812 252298
rect 260652 252062 260708 252118
rect 254994 244294 255050 244350
rect 255118 244294 255174 244350
rect 255242 244294 255298 244350
rect 255366 244294 255422 244350
rect 254994 244170 255050 244226
rect 255118 244170 255174 244226
rect 255242 244170 255298 244226
rect 255366 244170 255422 244226
rect 254994 244046 255050 244102
rect 255118 244046 255174 244102
rect 255242 244046 255298 244102
rect 255366 244046 255422 244102
rect 254994 243922 255050 243978
rect 255118 243922 255174 243978
rect 255242 243922 255298 243978
rect 255366 243922 255422 243978
rect 254994 226294 255050 226350
rect 255118 226294 255174 226350
rect 255242 226294 255298 226350
rect 255366 226294 255422 226350
rect 254994 226170 255050 226226
rect 255118 226170 255174 226226
rect 255242 226170 255298 226226
rect 255366 226170 255422 226226
rect 254994 226046 255050 226102
rect 255118 226046 255174 226102
rect 255242 226046 255298 226102
rect 255366 226046 255422 226102
rect 254994 225922 255050 225978
rect 255118 225922 255174 225978
rect 255242 225922 255298 225978
rect 255366 225922 255422 225978
rect 75238 202294 75294 202350
rect 75362 202294 75418 202350
rect 75238 202170 75294 202226
rect 75362 202170 75418 202226
rect 75238 202046 75294 202102
rect 75362 202046 75418 202102
rect 75238 201922 75294 201978
rect 75362 201922 75418 201978
rect 105958 202294 106014 202350
rect 106082 202294 106138 202350
rect 105958 202170 106014 202226
rect 106082 202170 106138 202226
rect 105958 202046 106014 202102
rect 106082 202046 106138 202102
rect 105958 201922 106014 201978
rect 106082 201922 106138 201978
rect 136678 202294 136734 202350
rect 136802 202294 136858 202350
rect 136678 202170 136734 202226
rect 136802 202170 136858 202226
rect 136678 202046 136734 202102
rect 136802 202046 136858 202102
rect 136678 201922 136734 201978
rect 136802 201922 136858 201978
rect 167398 202294 167454 202350
rect 167522 202294 167578 202350
rect 167398 202170 167454 202226
rect 167522 202170 167578 202226
rect 167398 202046 167454 202102
rect 167522 202046 167578 202102
rect 167398 201922 167454 201978
rect 167522 201922 167578 201978
rect 198118 202294 198174 202350
rect 198242 202294 198298 202350
rect 198118 202170 198174 202226
rect 198242 202170 198298 202226
rect 198118 202046 198174 202102
rect 198242 202046 198298 202102
rect 198118 201922 198174 201978
rect 198242 201922 198298 201978
rect 228838 202294 228894 202350
rect 228962 202294 229018 202350
rect 228838 202170 228894 202226
rect 228962 202170 229018 202226
rect 228838 202046 228894 202102
rect 228962 202046 229018 202102
rect 228838 201922 228894 201978
rect 228962 201922 229018 201978
rect 259558 202294 259614 202350
rect 259682 202294 259738 202350
rect 259558 202170 259614 202226
rect 259682 202170 259738 202226
rect 259558 202046 259614 202102
rect 259682 202046 259738 202102
rect 259558 201922 259614 201978
rect 259682 201922 259738 201978
rect 59878 190294 59934 190350
rect 60002 190294 60058 190350
rect 59878 190170 59934 190226
rect 60002 190170 60058 190226
rect 59878 190046 59934 190102
rect 60002 190046 60058 190102
rect 59878 189922 59934 189978
rect 60002 189922 60058 189978
rect 90598 190294 90654 190350
rect 90722 190294 90778 190350
rect 90598 190170 90654 190226
rect 90722 190170 90778 190226
rect 90598 190046 90654 190102
rect 90722 190046 90778 190102
rect 90598 189922 90654 189978
rect 90722 189922 90778 189978
rect 121318 190294 121374 190350
rect 121442 190294 121498 190350
rect 121318 190170 121374 190226
rect 121442 190170 121498 190226
rect 121318 190046 121374 190102
rect 121442 190046 121498 190102
rect 121318 189922 121374 189978
rect 121442 189922 121498 189978
rect 152038 190294 152094 190350
rect 152162 190294 152218 190350
rect 152038 190170 152094 190226
rect 152162 190170 152218 190226
rect 152038 190046 152094 190102
rect 152162 190046 152218 190102
rect 152038 189922 152094 189978
rect 152162 189922 152218 189978
rect 182758 190294 182814 190350
rect 182882 190294 182938 190350
rect 182758 190170 182814 190226
rect 182882 190170 182938 190226
rect 182758 190046 182814 190102
rect 182882 190046 182938 190102
rect 182758 189922 182814 189978
rect 182882 189922 182938 189978
rect 213478 190294 213534 190350
rect 213602 190294 213658 190350
rect 213478 190170 213534 190226
rect 213602 190170 213658 190226
rect 213478 190046 213534 190102
rect 213602 190046 213658 190102
rect 213478 189922 213534 189978
rect 213602 189922 213658 189978
rect 244198 190294 244254 190350
rect 244322 190294 244378 190350
rect 244198 190170 244254 190226
rect 244322 190170 244378 190226
rect 244198 190046 244254 190102
rect 244322 190046 244378 190102
rect 244198 189922 244254 189978
rect 244322 189922 244378 189978
rect 75238 184294 75294 184350
rect 75362 184294 75418 184350
rect 75238 184170 75294 184226
rect 75362 184170 75418 184226
rect 75238 184046 75294 184102
rect 75362 184046 75418 184102
rect 75238 183922 75294 183978
rect 75362 183922 75418 183978
rect 105958 184294 106014 184350
rect 106082 184294 106138 184350
rect 105958 184170 106014 184226
rect 106082 184170 106138 184226
rect 105958 184046 106014 184102
rect 106082 184046 106138 184102
rect 105958 183922 106014 183978
rect 106082 183922 106138 183978
rect 136678 184294 136734 184350
rect 136802 184294 136858 184350
rect 136678 184170 136734 184226
rect 136802 184170 136858 184226
rect 136678 184046 136734 184102
rect 136802 184046 136858 184102
rect 136678 183922 136734 183978
rect 136802 183922 136858 183978
rect 167398 184294 167454 184350
rect 167522 184294 167578 184350
rect 167398 184170 167454 184226
rect 167522 184170 167578 184226
rect 167398 184046 167454 184102
rect 167522 184046 167578 184102
rect 167398 183922 167454 183978
rect 167522 183922 167578 183978
rect 198118 184294 198174 184350
rect 198242 184294 198298 184350
rect 198118 184170 198174 184226
rect 198242 184170 198298 184226
rect 198118 184046 198174 184102
rect 198242 184046 198298 184102
rect 198118 183922 198174 183978
rect 198242 183922 198298 183978
rect 228838 184294 228894 184350
rect 228962 184294 229018 184350
rect 228838 184170 228894 184226
rect 228962 184170 229018 184226
rect 228838 184046 228894 184102
rect 228962 184046 229018 184102
rect 228838 183922 228894 183978
rect 228962 183922 229018 183978
rect 259558 184294 259614 184350
rect 259682 184294 259738 184350
rect 259558 184170 259614 184226
rect 259682 184170 259738 184226
rect 259558 184046 259614 184102
rect 259682 184046 259738 184102
rect 259558 183922 259614 183978
rect 259682 183922 259738 183978
rect 59878 172294 59934 172350
rect 60002 172294 60058 172350
rect 59878 172170 59934 172226
rect 60002 172170 60058 172226
rect 59878 172046 59934 172102
rect 60002 172046 60058 172102
rect 59878 171922 59934 171978
rect 60002 171922 60058 171978
rect 90598 172294 90654 172350
rect 90722 172294 90778 172350
rect 90598 172170 90654 172226
rect 90722 172170 90778 172226
rect 90598 172046 90654 172102
rect 90722 172046 90778 172102
rect 90598 171922 90654 171978
rect 90722 171922 90778 171978
rect 121318 172294 121374 172350
rect 121442 172294 121498 172350
rect 121318 172170 121374 172226
rect 121442 172170 121498 172226
rect 121318 172046 121374 172102
rect 121442 172046 121498 172102
rect 121318 171922 121374 171978
rect 121442 171922 121498 171978
rect 152038 172294 152094 172350
rect 152162 172294 152218 172350
rect 152038 172170 152094 172226
rect 152162 172170 152218 172226
rect 152038 172046 152094 172102
rect 152162 172046 152218 172102
rect 152038 171922 152094 171978
rect 152162 171922 152218 171978
rect 182758 172294 182814 172350
rect 182882 172294 182938 172350
rect 182758 172170 182814 172226
rect 182882 172170 182938 172226
rect 182758 172046 182814 172102
rect 182882 172046 182938 172102
rect 182758 171922 182814 171978
rect 182882 171922 182938 171978
rect 213478 172294 213534 172350
rect 213602 172294 213658 172350
rect 213478 172170 213534 172226
rect 213602 172170 213658 172226
rect 213478 172046 213534 172102
rect 213602 172046 213658 172102
rect 213478 171922 213534 171978
rect 213602 171922 213658 171978
rect 244198 172294 244254 172350
rect 244322 172294 244378 172350
rect 244198 172170 244254 172226
rect 244322 172170 244378 172226
rect 244198 172046 244254 172102
rect 244322 172046 244378 172102
rect 244198 171922 244254 171978
rect 244322 171922 244378 171978
rect 75238 166294 75294 166350
rect 75362 166294 75418 166350
rect 75238 166170 75294 166226
rect 75362 166170 75418 166226
rect 75238 166046 75294 166102
rect 75362 166046 75418 166102
rect 75238 165922 75294 165978
rect 75362 165922 75418 165978
rect 105958 166294 106014 166350
rect 106082 166294 106138 166350
rect 105958 166170 106014 166226
rect 106082 166170 106138 166226
rect 105958 166046 106014 166102
rect 106082 166046 106138 166102
rect 105958 165922 106014 165978
rect 106082 165922 106138 165978
rect 136678 166294 136734 166350
rect 136802 166294 136858 166350
rect 136678 166170 136734 166226
rect 136802 166170 136858 166226
rect 136678 166046 136734 166102
rect 136802 166046 136858 166102
rect 136678 165922 136734 165978
rect 136802 165922 136858 165978
rect 167398 166294 167454 166350
rect 167522 166294 167578 166350
rect 167398 166170 167454 166226
rect 167522 166170 167578 166226
rect 167398 166046 167454 166102
rect 167522 166046 167578 166102
rect 167398 165922 167454 165978
rect 167522 165922 167578 165978
rect 198118 166294 198174 166350
rect 198242 166294 198298 166350
rect 198118 166170 198174 166226
rect 198242 166170 198298 166226
rect 198118 166046 198174 166102
rect 198242 166046 198298 166102
rect 198118 165922 198174 165978
rect 198242 165922 198298 165978
rect 228838 166294 228894 166350
rect 228962 166294 229018 166350
rect 228838 166170 228894 166226
rect 228962 166170 229018 166226
rect 228838 166046 228894 166102
rect 228962 166046 229018 166102
rect 228838 165922 228894 165978
rect 228962 165922 229018 165978
rect 259558 166294 259614 166350
rect 259682 166294 259738 166350
rect 259558 166170 259614 166226
rect 259682 166170 259738 166226
rect 259558 166046 259614 166102
rect 259682 166046 259738 166102
rect 259558 165922 259614 165978
rect 259682 165922 259738 165978
rect 59878 154294 59934 154350
rect 60002 154294 60058 154350
rect 59878 154170 59934 154226
rect 60002 154170 60058 154226
rect 59878 154046 59934 154102
rect 60002 154046 60058 154102
rect 59878 153922 59934 153978
rect 60002 153922 60058 153978
rect 90598 154294 90654 154350
rect 90722 154294 90778 154350
rect 90598 154170 90654 154226
rect 90722 154170 90778 154226
rect 90598 154046 90654 154102
rect 90722 154046 90778 154102
rect 90598 153922 90654 153978
rect 90722 153922 90778 153978
rect 121318 154294 121374 154350
rect 121442 154294 121498 154350
rect 121318 154170 121374 154226
rect 121442 154170 121498 154226
rect 121318 154046 121374 154102
rect 121442 154046 121498 154102
rect 121318 153922 121374 153978
rect 121442 153922 121498 153978
rect 152038 154294 152094 154350
rect 152162 154294 152218 154350
rect 152038 154170 152094 154226
rect 152162 154170 152218 154226
rect 152038 154046 152094 154102
rect 152162 154046 152218 154102
rect 152038 153922 152094 153978
rect 152162 153922 152218 153978
rect 182758 154294 182814 154350
rect 182882 154294 182938 154350
rect 182758 154170 182814 154226
rect 182882 154170 182938 154226
rect 182758 154046 182814 154102
rect 182882 154046 182938 154102
rect 182758 153922 182814 153978
rect 182882 153922 182938 153978
rect 213478 154294 213534 154350
rect 213602 154294 213658 154350
rect 213478 154170 213534 154226
rect 213602 154170 213658 154226
rect 213478 154046 213534 154102
rect 213602 154046 213658 154102
rect 213478 153922 213534 153978
rect 213602 153922 213658 153978
rect 244198 154294 244254 154350
rect 244322 154294 244378 154350
rect 244198 154170 244254 154226
rect 244322 154170 244378 154226
rect 244198 154046 244254 154102
rect 244322 154046 244378 154102
rect 244198 153922 244254 153978
rect 244322 153922 244378 153978
rect 75238 148294 75294 148350
rect 75362 148294 75418 148350
rect 75238 148170 75294 148226
rect 75362 148170 75418 148226
rect 75238 148046 75294 148102
rect 75362 148046 75418 148102
rect 75238 147922 75294 147978
rect 75362 147922 75418 147978
rect 105958 148294 106014 148350
rect 106082 148294 106138 148350
rect 105958 148170 106014 148226
rect 106082 148170 106138 148226
rect 105958 148046 106014 148102
rect 106082 148046 106138 148102
rect 105958 147922 106014 147978
rect 106082 147922 106138 147978
rect 136678 148294 136734 148350
rect 136802 148294 136858 148350
rect 136678 148170 136734 148226
rect 136802 148170 136858 148226
rect 136678 148046 136734 148102
rect 136802 148046 136858 148102
rect 136678 147922 136734 147978
rect 136802 147922 136858 147978
rect 167398 148294 167454 148350
rect 167522 148294 167578 148350
rect 167398 148170 167454 148226
rect 167522 148170 167578 148226
rect 167398 148046 167454 148102
rect 167522 148046 167578 148102
rect 167398 147922 167454 147978
rect 167522 147922 167578 147978
rect 198118 148294 198174 148350
rect 198242 148294 198298 148350
rect 198118 148170 198174 148226
rect 198242 148170 198298 148226
rect 198118 148046 198174 148102
rect 198242 148046 198298 148102
rect 198118 147922 198174 147978
rect 198242 147922 198298 147978
rect 228838 148294 228894 148350
rect 228962 148294 229018 148350
rect 228838 148170 228894 148226
rect 228962 148170 229018 148226
rect 228838 148046 228894 148102
rect 228962 148046 229018 148102
rect 228838 147922 228894 147978
rect 228962 147922 229018 147978
rect 259558 148294 259614 148350
rect 259682 148294 259738 148350
rect 259558 148170 259614 148226
rect 259682 148170 259738 148226
rect 259558 148046 259614 148102
rect 259682 148046 259738 148102
rect 259558 147922 259614 147978
rect 259682 147922 259738 147978
rect 59878 136294 59934 136350
rect 60002 136294 60058 136350
rect 59878 136170 59934 136226
rect 60002 136170 60058 136226
rect 59878 136046 59934 136102
rect 60002 136046 60058 136102
rect 59878 135922 59934 135978
rect 60002 135922 60058 135978
rect 90598 136294 90654 136350
rect 90722 136294 90778 136350
rect 90598 136170 90654 136226
rect 90722 136170 90778 136226
rect 90598 136046 90654 136102
rect 90722 136046 90778 136102
rect 90598 135922 90654 135978
rect 90722 135922 90778 135978
rect 121318 136294 121374 136350
rect 121442 136294 121498 136350
rect 121318 136170 121374 136226
rect 121442 136170 121498 136226
rect 121318 136046 121374 136102
rect 121442 136046 121498 136102
rect 121318 135922 121374 135978
rect 121442 135922 121498 135978
rect 152038 136294 152094 136350
rect 152162 136294 152218 136350
rect 152038 136170 152094 136226
rect 152162 136170 152218 136226
rect 152038 136046 152094 136102
rect 152162 136046 152218 136102
rect 152038 135922 152094 135978
rect 152162 135922 152218 135978
rect 182758 136294 182814 136350
rect 182882 136294 182938 136350
rect 182758 136170 182814 136226
rect 182882 136170 182938 136226
rect 182758 136046 182814 136102
rect 182882 136046 182938 136102
rect 182758 135922 182814 135978
rect 182882 135922 182938 135978
rect 213478 136294 213534 136350
rect 213602 136294 213658 136350
rect 213478 136170 213534 136226
rect 213602 136170 213658 136226
rect 213478 136046 213534 136102
rect 213602 136046 213658 136102
rect 213478 135922 213534 135978
rect 213602 135922 213658 135978
rect 244198 136294 244254 136350
rect 244322 136294 244378 136350
rect 244198 136170 244254 136226
rect 244322 136170 244378 136226
rect 244198 136046 244254 136102
rect 244322 136046 244378 136102
rect 244198 135922 244254 135978
rect 244322 135922 244378 135978
rect 75238 130294 75294 130350
rect 75362 130294 75418 130350
rect 75238 130170 75294 130226
rect 75362 130170 75418 130226
rect 75238 130046 75294 130102
rect 75362 130046 75418 130102
rect 75238 129922 75294 129978
rect 75362 129922 75418 129978
rect 105958 130294 106014 130350
rect 106082 130294 106138 130350
rect 105958 130170 106014 130226
rect 106082 130170 106138 130226
rect 105958 130046 106014 130102
rect 106082 130046 106138 130102
rect 105958 129922 106014 129978
rect 106082 129922 106138 129978
rect 136678 130294 136734 130350
rect 136802 130294 136858 130350
rect 136678 130170 136734 130226
rect 136802 130170 136858 130226
rect 136678 130046 136734 130102
rect 136802 130046 136858 130102
rect 136678 129922 136734 129978
rect 136802 129922 136858 129978
rect 167398 130294 167454 130350
rect 167522 130294 167578 130350
rect 167398 130170 167454 130226
rect 167522 130170 167578 130226
rect 167398 130046 167454 130102
rect 167522 130046 167578 130102
rect 167398 129922 167454 129978
rect 167522 129922 167578 129978
rect 198118 130294 198174 130350
rect 198242 130294 198298 130350
rect 198118 130170 198174 130226
rect 198242 130170 198298 130226
rect 198118 130046 198174 130102
rect 198242 130046 198298 130102
rect 198118 129922 198174 129978
rect 198242 129922 198298 129978
rect 228838 130294 228894 130350
rect 228962 130294 229018 130350
rect 228838 130170 228894 130226
rect 228962 130170 229018 130226
rect 228838 130046 228894 130102
rect 228962 130046 229018 130102
rect 228838 129922 228894 129978
rect 228962 129922 229018 129978
rect 259558 130294 259614 130350
rect 259682 130294 259738 130350
rect 259558 130170 259614 130226
rect 259682 130170 259738 130226
rect 259558 130046 259614 130102
rect 259682 130046 259738 130102
rect 259558 129922 259614 129978
rect 259682 129922 259738 129978
rect 59878 118294 59934 118350
rect 60002 118294 60058 118350
rect 59878 118170 59934 118226
rect 60002 118170 60058 118226
rect 59878 118046 59934 118102
rect 60002 118046 60058 118102
rect 59878 117922 59934 117978
rect 60002 117922 60058 117978
rect 90598 118294 90654 118350
rect 90722 118294 90778 118350
rect 90598 118170 90654 118226
rect 90722 118170 90778 118226
rect 90598 118046 90654 118102
rect 90722 118046 90778 118102
rect 90598 117922 90654 117978
rect 90722 117922 90778 117978
rect 121318 118294 121374 118350
rect 121442 118294 121498 118350
rect 121318 118170 121374 118226
rect 121442 118170 121498 118226
rect 121318 118046 121374 118102
rect 121442 118046 121498 118102
rect 121318 117922 121374 117978
rect 121442 117922 121498 117978
rect 152038 118294 152094 118350
rect 152162 118294 152218 118350
rect 152038 118170 152094 118226
rect 152162 118170 152218 118226
rect 152038 118046 152094 118102
rect 152162 118046 152218 118102
rect 152038 117922 152094 117978
rect 152162 117922 152218 117978
rect 182758 118294 182814 118350
rect 182882 118294 182938 118350
rect 182758 118170 182814 118226
rect 182882 118170 182938 118226
rect 182758 118046 182814 118102
rect 182882 118046 182938 118102
rect 182758 117922 182814 117978
rect 182882 117922 182938 117978
rect 213478 118294 213534 118350
rect 213602 118294 213658 118350
rect 213478 118170 213534 118226
rect 213602 118170 213658 118226
rect 213478 118046 213534 118102
rect 213602 118046 213658 118102
rect 213478 117922 213534 117978
rect 213602 117922 213658 117978
rect 244198 118294 244254 118350
rect 244322 118294 244378 118350
rect 244198 118170 244254 118226
rect 244322 118170 244378 118226
rect 244198 118046 244254 118102
rect 244322 118046 244378 118102
rect 244198 117922 244254 117978
rect 244322 117922 244378 117978
rect 75238 112294 75294 112350
rect 75362 112294 75418 112350
rect 75238 112170 75294 112226
rect 75362 112170 75418 112226
rect 75238 112046 75294 112102
rect 75362 112046 75418 112102
rect 75238 111922 75294 111978
rect 75362 111922 75418 111978
rect 105958 112294 106014 112350
rect 106082 112294 106138 112350
rect 105958 112170 106014 112226
rect 106082 112170 106138 112226
rect 105958 112046 106014 112102
rect 106082 112046 106138 112102
rect 105958 111922 106014 111978
rect 106082 111922 106138 111978
rect 136678 112294 136734 112350
rect 136802 112294 136858 112350
rect 136678 112170 136734 112226
rect 136802 112170 136858 112226
rect 136678 112046 136734 112102
rect 136802 112046 136858 112102
rect 136678 111922 136734 111978
rect 136802 111922 136858 111978
rect 167398 112294 167454 112350
rect 167522 112294 167578 112350
rect 167398 112170 167454 112226
rect 167522 112170 167578 112226
rect 167398 112046 167454 112102
rect 167522 112046 167578 112102
rect 167398 111922 167454 111978
rect 167522 111922 167578 111978
rect 198118 112294 198174 112350
rect 198242 112294 198298 112350
rect 198118 112170 198174 112226
rect 198242 112170 198298 112226
rect 198118 112046 198174 112102
rect 198242 112046 198298 112102
rect 198118 111922 198174 111978
rect 198242 111922 198298 111978
rect 228838 112294 228894 112350
rect 228962 112294 229018 112350
rect 228838 112170 228894 112226
rect 228962 112170 229018 112226
rect 228838 112046 228894 112102
rect 228962 112046 229018 112102
rect 228838 111922 228894 111978
rect 228962 111922 229018 111978
rect 259558 112294 259614 112350
rect 259682 112294 259738 112350
rect 259558 112170 259614 112226
rect 259682 112170 259738 112226
rect 259558 112046 259614 112102
rect 259682 112046 259738 112102
rect 259558 111922 259614 111978
rect 259682 111922 259738 111978
rect 59878 100294 59934 100350
rect 60002 100294 60058 100350
rect 59878 100170 59934 100226
rect 60002 100170 60058 100226
rect 59878 100046 59934 100102
rect 60002 100046 60058 100102
rect 59878 99922 59934 99978
rect 60002 99922 60058 99978
rect 90598 100294 90654 100350
rect 90722 100294 90778 100350
rect 90598 100170 90654 100226
rect 90722 100170 90778 100226
rect 90598 100046 90654 100102
rect 90722 100046 90778 100102
rect 90598 99922 90654 99978
rect 90722 99922 90778 99978
rect 121318 100294 121374 100350
rect 121442 100294 121498 100350
rect 121318 100170 121374 100226
rect 121442 100170 121498 100226
rect 121318 100046 121374 100102
rect 121442 100046 121498 100102
rect 121318 99922 121374 99978
rect 121442 99922 121498 99978
rect 152038 100294 152094 100350
rect 152162 100294 152218 100350
rect 152038 100170 152094 100226
rect 152162 100170 152218 100226
rect 152038 100046 152094 100102
rect 152162 100046 152218 100102
rect 152038 99922 152094 99978
rect 152162 99922 152218 99978
rect 182758 100294 182814 100350
rect 182882 100294 182938 100350
rect 182758 100170 182814 100226
rect 182882 100170 182938 100226
rect 182758 100046 182814 100102
rect 182882 100046 182938 100102
rect 182758 99922 182814 99978
rect 182882 99922 182938 99978
rect 213478 100294 213534 100350
rect 213602 100294 213658 100350
rect 213478 100170 213534 100226
rect 213602 100170 213658 100226
rect 213478 100046 213534 100102
rect 213602 100046 213658 100102
rect 213478 99922 213534 99978
rect 213602 99922 213658 99978
rect 244198 100294 244254 100350
rect 244322 100294 244378 100350
rect 244198 100170 244254 100226
rect 244322 100170 244378 100226
rect 244198 100046 244254 100102
rect 244322 100046 244378 100102
rect 244198 99922 244254 99978
rect 244322 99922 244378 99978
rect 75238 94294 75294 94350
rect 75362 94294 75418 94350
rect 75238 94170 75294 94226
rect 75362 94170 75418 94226
rect 75238 94046 75294 94102
rect 75362 94046 75418 94102
rect 75238 93922 75294 93978
rect 75362 93922 75418 93978
rect 105958 94294 106014 94350
rect 106082 94294 106138 94350
rect 105958 94170 106014 94226
rect 106082 94170 106138 94226
rect 105958 94046 106014 94102
rect 106082 94046 106138 94102
rect 105958 93922 106014 93978
rect 106082 93922 106138 93978
rect 136678 94294 136734 94350
rect 136802 94294 136858 94350
rect 136678 94170 136734 94226
rect 136802 94170 136858 94226
rect 136678 94046 136734 94102
rect 136802 94046 136858 94102
rect 136678 93922 136734 93978
rect 136802 93922 136858 93978
rect 167398 94294 167454 94350
rect 167522 94294 167578 94350
rect 167398 94170 167454 94226
rect 167522 94170 167578 94226
rect 167398 94046 167454 94102
rect 167522 94046 167578 94102
rect 167398 93922 167454 93978
rect 167522 93922 167578 93978
rect 198118 94294 198174 94350
rect 198242 94294 198298 94350
rect 198118 94170 198174 94226
rect 198242 94170 198298 94226
rect 198118 94046 198174 94102
rect 198242 94046 198298 94102
rect 198118 93922 198174 93978
rect 198242 93922 198298 93978
rect 228838 94294 228894 94350
rect 228962 94294 229018 94350
rect 228838 94170 228894 94226
rect 228962 94170 229018 94226
rect 228838 94046 228894 94102
rect 228962 94046 229018 94102
rect 228838 93922 228894 93978
rect 228962 93922 229018 93978
rect 259558 94294 259614 94350
rect 259682 94294 259738 94350
rect 259558 94170 259614 94226
rect 259682 94170 259738 94226
rect 259558 94046 259614 94102
rect 259682 94046 259738 94102
rect 259558 93922 259614 93978
rect 259682 93922 259738 93978
rect 59878 82294 59934 82350
rect 60002 82294 60058 82350
rect 59878 82170 59934 82226
rect 60002 82170 60058 82226
rect 59878 82046 59934 82102
rect 60002 82046 60058 82102
rect 59878 81922 59934 81978
rect 60002 81922 60058 81978
rect 90598 82294 90654 82350
rect 90722 82294 90778 82350
rect 90598 82170 90654 82226
rect 90722 82170 90778 82226
rect 90598 82046 90654 82102
rect 90722 82046 90778 82102
rect 90598 81922 90654 81978
rect 90722 81922 90778 81978
rect 121318 82294 121374 82350
rect 121442 82294 121498 82350
rect 121318 82170 121374 82226
rect 121442 82170 121498 82226
rect 121318 82046 121374 82102
rect 121442 82046 121498 82102
rect 121318 81922 121374 81978
rect 121442 81922 121498 81978
rect 152038 82294 152094 82350
rect 152162 82294 152218 82350
rect 152038 82170 152094 82226
rect 152162 82170 152218 82226
rect 152038 82046 152094 82102
rect 152162 82046 152218 82102
rect 152038 81922 152094 81978
rect 152162 81922 152218 81978
rect 182758 82294 182814 82350
rect 182882 82294 182938 82350
rect 182758 82170 182814 82226
rect 182882 82170 182938 82226
rect 182758 82046 182814 82102
rect 182882 82046 182938 82102
rect 182758 81922 182814 81978
rect 182882 81922 182938 81978
rect 213478 82294 213534 82350
rect 213602 82294 213658 82350
rect 213478 82170 213534 82226
rect 213602 82170 213658 82226
rect 213478 82046 213534 82102
rect 213602 82046 213658 82102
rect 213478 81922 213534 81978
rect 213602 81922 213658 81978
rect 244198 82294 244254 82350
rect 244322 82294 244378 82350
rect 244198 82170 244254 82226
rect 244322 82170 244378 82226
rect 244198 82046 244254 82102
rect 244322 82046 244378 82102
rect 244198 81922 244254 81978
rect 244322 81922 244378 81978
rect 75238 76294 75294 76350
rect 75362 76294 75418 76350
rect 75238 76170 75294 76226
rect 75362 76170 75418 76226
rect 75238 76046 75294 76102
rect 75362 76046 75418 76102
rect 75238 75922 75294 75978
rect 75362 75922 75418 75978
rect 105958 76294 106014 76350
rect 106082 76294 106138 76350
rect 105958 76170 106014 76226
rect 106082 76170 106138 76226
rect 105958 76046 106014 76102
rect 106082 76046 106138 76102
rect 105958 75922 106014 75978
rect 106082 75922 106138 75978
rect 136678 76294 136734 76350
rect 136802 76294 136858 76350
rect 136678 76170 136734 76226
rect 136802 76170 136858 76226
rect 136678 76046 136734 76102
rect 136802 76046 136858 76102
rect 136678 75922 136734 75978
rect 136802 75922 136858 75978
rect 167398 76294 167454 76350
rect 167522 76294 167578 76350
rect 167398 76170 167454 76226
rect 167522 76170 167578 76226
rect 167398 76046 167454 76102
rect 167522 76046 167578 76102
rect 167398 75922 167454 75978
rect 167522 75922 167578 75978
rect 198118 76294 198174 76350
rect 198242 76294 198298 76350
rect 198118 76170 198174 76226
rect 198242 76170 198298 76226
rect 198118 76046 198174 76102
rect 198242 76046 198298 76102
rect 198118 75922 198174 75978
rect 198242 75922 198298 75978
rect 228838 76294 228894 76350
rect 228962 76294 229018 76350
rect 228838 76170 228894 76226
rect 228962 76170 229018 76226
rect 228838 76046 228894 76102
rect 228962 76046 229018 76102
rect 228838 75922 228894 75978
rect 228962 75922 229018 75978
rect 259558 76294 259614 76350
rect 259682 76294 259738 76350
rect 259558 76170 259614 76226
rect 259682 76170 259738 76226
rect 259558 76046 259614 76102
rect 259682 76046 259738 76102
rect 259558 75922 259614 75978
rect 259682 75922 259738 75978
rect 59878 64294 59934 64350
rect 60002 64294 60058 64350
rect 59878 64170 59934 64226
rect 60002 64170 60058 64226
rect 59878 64046 59934 64102
rect 60002 64046 60058 64102
rect 59878 63922 59934 63978
rect 60002 63922 60058 63978
rect 90598 64294 90654 64350
rect 90722 64294 90778 64350
rect 90598 64170 90654 64226
rect 90722 64170 90778 64226
rect 90598 64046 90654 64102
rect 90722 64046 90778 64102
rect 90598 63922 90654 63978
rect 90722 63922 90778 63978
rect 121318 64294 121374 64350
rect 121442 64294 121498 64350
rect 121318 64170 121374 64226
rect 121442 64170 121498 64226
rect 121318 64046 121374 64102
rect 121442 64046 121498 64102
rect 121318 63922 121374 63978
rect 121442 63922 121498 63978
rect 152038 64294 152094 64350
rect 152162 64294 152218 64350
rect 152038 64170 152094 64226
rect 152162 64170 152218 64226
rect 152038 64046 152094 64102
rect 152162 64046 152218 64102
rect 152038 63922 152094 63978
rect 152162 63922 152218 63978
rect 182758 64294 182814 64350
rect 182882 64294 182938 64350
rect 182758 64170 182814 64226
rect 182882 64170 182938 64226
rect 182758 64046 182814 64102
rect 182882 64046 182938 64102
rect 182758 63922 182814 63978
rect 182882 63922 182938 63978
rect 213478 64294 213534 64350
rect 213602 64294 213658 64350
rect 213478 64170 213534 64226
rect 213602 64170 213658 64226
rect 213478 64046 213534 64102
rect 213602 64046 213658 64102
rect 213478 63922 213534 63978
rect 213602 63922 213658 63978
rect 244198 64294 244254 64350
rect 244322 64294 244378 64350
rect 244198 64170 244254 64226
rect 244322 64170 244378 64226
rect 244198 64046 244254 64102
rect 244322 64046 244378 64102
rect 244198 63922 244254 63978
rect 244322 63922 244378 63978
rect 75238 58294 75294 58350
rect 75362 58294 75418 58350
rect 75238 58170 75294 58226
rect 75362 58170 75418 58226
rect 75238 58046 75294 58102
rect 75362 58046 75418 58102
rect 75238 57922 75294 57978
rect 75362 57922 75418 57978
rect 105958 58294 106014 58350
rect 106082 58294 106138 58350
rect 105958 58170 106014 58226
rect 106082 58170 106138 58226
rect 105958 58046 106014 58102
rect 106082 58046 106138 58102
rect 105958 57922 106014 57978
rect 106082 57922 106138 57978
rect 136678 58294 136734 58350
rect 136802 58294 136858 58350
rect 136678 58170 136734 58226
rect 136802 58170 136858 58226
rect 136678 58046 136734 58102
rect 136802 58046 136858 58102
rect 136678 57922 136734 57978
rect 136802 57922 136858 57978
rect 167398 58294 167454 58350
rect 167522 58294 167578 58350
rect 167398 58170 167454 58226
rect 167522 58170 167578 58226
rect 167398 58046 167454 58102
rect 167522 58046 167578 58102
rect 167398 57922 167454 57978
rect 167522 57922 167578 57978
rect 198118 58294 198174 58350
rect 198242 58294 198298 58350
rect 198118 58170 198174 58226
rect 198242 58170 198298 58226
rect 198118 58046 198174 58102
rect 198242 58046 198298 58102
rect 198118 57922 198174 57978
rect 198242 57922 198298 57978
rect 228838 58294 228894 58350
rect 228962 58294 229018 58350
rect 228838 58170 228894 58226
rect 228962 58170 229018 58226
rect 228838 58046 228894 58102
rect 228962 58046 229018 58102
rect 228838 57922 228894 57978
rect 228962 57922 229018 57978
rect 259558 58294 259614 58350
rect 259682 58294 259738 58350
rect 259558 58170 259614 58226
rect 259682 58170 259738 58226
rect 259558 58046 259614 58102
rect 259682 58046 259738 58102
rect 259558 57922 259614 57978
rect 259682 57922 259738 57978
rect 66954 40294 67010 40350
rect 67078 40294 67134 40350
rect 67202 40294 67258 40350
rect 67326 40294 67382 40350
rect 66954 40170 67010 40226
rect 67078 40170 67134 40226
rect 67202 40170 67258 40226
rect 67326 40170 67382 40226
rect 66954 40046 67010 40102
rect 67078 40046 67134 40102
rect 67202 40046 67258 40102
rect 67326 40046 67382 40102
rect 66954 39922 67010 39978
rect 67078 39922 67134 39978
rect 67202 39922 67258 39978
rect 67326 39922 67382 39978
rect 66954 22294 67010 22350
rect 67078 22294 67134 22350
rect 67202 22294 67258 22350
rect 67326 22294 67382 22350
rect 66954 22170 67010 22226
rect 67078 22170 67134 22226
rect 67202 22170 67258 22226
rect 67326 22170 67382 22226
rect 66954 22046 67010 22102
rect 67078 22046 67134 22102
rect 67202 22046 67258 22102
rect 67326 22046 67382 22102
rect 66954 21922 67010 21978
rect 67078 21922 67134 21978
rect 67202 21922 67258 21978
rect 67326 21922 67382 21978
rect 39954 -1176 40010 -1120
rect 40078 -1176 40134 -1120
rect 40202 -1176 40258 -1120
rect 40326 -1176 40382 -1120
rect 39954 -1300 40010 -1244
rect 40078 -1300 40134 -1244
rect 40202 -1300 40258 -1244
rect 40326 -1300 40382 -1244
rect 39954 -1424 40010 -1368
rect 40078 -1424 40134 -1368
rect 40202 -1424 40258 -1368
rect 40326 -1424 40382 -1368
rect 39954 -1548 40010 -1492
rect 40078 -1548 40134 -1492
rect 40202 -1548 40258 -1492
rect 40326 -1548 40382 -1492
rect 66954 4294 67010 4350
rect 67078 4294 67134 4350
rect 67202 4294 67258 4350
rect 67326 4294 67382 4350
rect 66954 4170 67010 4226
rect 67078 4170 67134 4226
rect 67202 4170 67258 4226
rect 67326 4170 67382 4226
rect 66954 4046 67010 4102
rect 67078 4046 67134 4102
rect 67202 4046 67258 4102
rect 67326 4046 67382 4102
rect 66954 3922 67010 3978
rect 67078 3922 67134 3978
rect 67202 3922 67258 3978
rect 67326 3922 67382 3978
rect 66954 -216 67010 -160
rect 67078 -216 67134 -160
rect 67202 -216 67258 -160
rect 67326 -216 67382 -160
rect 66954 -340 67010 -284
rect 67078 -340 67134 -284
rect 67202 -340 67258 -284
rect 67326 -340 67382 -284
rect 66954 -464 67010 -408
rect 67078 -464 67134 -408
rect 67202 -464 67258 -408
rect 67326 -464 67382 -408
rect 66954 -588 67010 -532
rect 67078 -588 67134 -532
rect 67202 -588 67258 -532
rect 67326 -588 67382 -532
rect 70674 46294 70730 46350
rect 70798 46294 70854 46350
rect 70922 46294 70978 46350
rect 71046 46294 71102 46350
rect 70674 46170 70730 46226
rect 70798 46170 70854 46226
rect 70922 46170 70978 46226
rect 71046 46170 71102 46226
rect 70674 46046 70730 46102
rect 70798 46046 70854 46102
rect 70922 46046 70978 46102
rect 71046 46046 71102 46102
rect 70674 45922 70730 45978
rect 70798 45922 70854 45978
rect 70922 45922 70978 45978
rect 71046 45922 71102 45978
rect 70674 28294 70730 28350
rect 70798 28294 70854 28350
rect 70922 28294 70978 28350
rect 71046 28294 71102 28350
rect 70674 28170 70730 28226
rect 70798 28170 70854 28226
rect 70922 28170 70978 28226
rect 71046 28170 71102 28226
rect 70674 28046 70730 28102
rect 70798 28046 70854 28102
rect 70922 28046 70978 28102
rect 71046 28046 71102 28102
rect 70674 27922 70730 27978
rect 70798 27922 70854 27978
rect 70922 27922 70978 27978
rect 71046 27922 71102 27978
rect 70674 10294 70730 10350
rect 70798 10294 70854 10350
rect 70922 10294 70978 10350
rect 71046 10294 71102 10350
rect 70674 10170 70730 10226
rect 70798 10170 70854 10226
rect 70922 10170 70978 10226
rect 71046 10170 71102 10226
rect 70674 10046 70730 10102
rect 70798 10046 70854 10102
rect 70922 10046 70978 10102
rect 71046 10046 71102 10102
rect 70674 9922 70730 9978
rect 70798 9922 70854 9978
rect 70922 9922 70978 9978
rect 71046 9922 71102 9978
rect 70674 -1176 70730 -1120
rect 70798 -1176 70854 -1120
rect 70922 -1176 70978 -1120
rect 71046 -1176 71102 -1120
rect 70674 -1300 70730 -1244
rect 70798 -1300 70854 -1244
rect 70922 -1300 70978 -1244
rect 71046 -1300 71102 -1244
rect 70674 -1424 70730 -1368
rect 70798 -1424 70854 -1368
rect 70922 -1424 70978 -1368
rect 71046 -1424 71102 -1368
rect 70674 -1548 70730 -1492
rect 70798 -1548 70854 -1492
rect 70922 -1548 70978 -1492
rect 71046 -1548 71102 -1492
rect 97674 40294 97730 40350
rect 97798 40294 97854 40350
rect 97922 40294 97978 40350
rect 98046 40294 98102 40350
rect 97674 40170 97730 40226
rect 97798 40170 97854 40226
rect 97922 40170 97978 40226
rect 98046 40170 98102 40226
rect 97674 40046 97730 40102
rect 97798 40046 97854 40102
rect 97922 40046 97978 40102
rect 98046 40046 98102 40102
rect 97674 39922 97730 39978
rect 97798 39922 97854 39978
rect 97922 39922 97978 39978
rect 98046 39922 98102 39978
rect 97674 22294 97730 22350
rect 97798 22294 97854 22350
rect 97922 22294 97978 22350
rect 98046 22294 98102 22350
rect 97674 22170 97730 22226
rect 97798 22170 97854 22226
rect 97922 22170 97978 22226
rect 98046 22170 98102 22226
rect 97674 22046 97730 22102
rect 97798 22046 97854 22102
rect 97922 22046 97978 22102
rect 98046 22046 98102 22102
rect 97674 21922 97730 21978
rect 97798 21922 97854 21978
rect 97922 21922 97978 21978
rect 98046 21922 98102 21978
rect 97674 4294 97730 4350
rect 97798 4294 97854 4350
rect 97922 4294 97978 4350
rect 98046 4294 98102 4350
rect 97674 4170 97730 4226
rect 97798 4170 97854 4226
rect 97922 4170 97978 4226
rect 98046 4170 98102 4226
rect 97674 4046 97730 4102
rect 97798 4046 97854 4102
rect 97922 4046 97978 4102
rect 98046 4046 98102 4102
rect 97674 3922 97730 3978
rect 97798 3922 97854 3978
rect 97922 3922 97978 3978
rect 98046 3922 98102 3978
rect 97674 -216 97730 -160
rect 97798 -216 97854 -160
rect 97922 -216 97978 -160
rect 98046 -216 98102 -160
rect 97674 -340 97730 -284
rect 97798 -340 97854 -284
rect 97922 -340 97978 -284
rect 98046 -340 98102 -284
rect 97674 -464 97730 -408
rect 97798 -464 97854 -408
rect 97922 -464 97978 -408
rect 98046 -464 98102 -408
rect 97674 -588 97730 -532
rect 97798 -588 97854 -532
rect 97922 -588 97978 -532
rect 98046 -588 98102 -532
rect 101394 46294 101450 46350
rect 101518 46294 101574 46350
rect 101642 46294 101698 46350
rect 101766 46294 101822 46350
rect 101394 46170 101450 46226
rect 101518 46170 101574 46226
rect 101642 46170 101698 46226
rect 101766 46170 101822 46226
rect 101394 46046 101450 46102
rect 101518 46046 101574 46102
rect 101642 46046 101698 46102
rect 101766 46046 101822 46102
rect 101394 45922 101450 45978
rect 101518 45922 101574 45978
rect 101642 45922 101698 45978
rect 101766 45922 101822 45978
rect 101394 28294 101450 28350
rect 101518 28294 101574 28350
rect 101642 28294 101698 28350
rect 101766 28294 101822 28350
rect 101394 28170 101450 28226
rect 101518 28170 101574 28226
rect 101642 28170 101698 28226
rect 101766 28170 101822 28226
rect 101394 28046 101450 28102
rect 101518 28046 101574 28102
rect 101642 28046 101698 28102
rect 101766 28046 101822 28102
rect 101394 27922 101450 27978
rect 101518 27922 101574 27978
rect 101642 27922 101698 27978
rect 101766 27922 101822 27978
rect 101394 10294 101450 10350
rect 101518 10294 101574 10350
rect 101642 10294 101698 10350
rect 101766 10294 101822 10350
rect 101394 10170 101450 10226
rect 101518 10170 101574 10226
rect 101642 10170 101698 10226
rect 101766 10170 101822 10226
rect 101394 10046 101450 10102
rect 101518 10046 101574 10102
rect 101642 10046 101698 10102
rect 101766 10046 101822 10102
rect 101394 9922 101450 9978
rect 101518 9922 101574 9978
rect 101642 9922 101698 9978
rect 101766 9922 101822 9978
rect 101394 -1176 101450 -1120
rect 101518 -1176 101574 -1120
rect 101642 -1176 101698 -1120
rect 101766 -1176 101822 -1120
rect 101394 -1300 101450 -1244
rect 101518 -1300 101574 -1244
rect 101642 -1300 101698 -1244
rect 101766 -1300 101822 -1244
rect 101394 -1424 101450 -1368
rect 101518 -1424 101574 -1368
rect 101642 -1424 101698 -1368
rect 101766 -1424 101822 -1368
rect 101394 -1548 101450 -1492
rect 101518 -1548 101574 -1492
rect 101642 -1548 101698 -1492
rect 101766 -1548 101822 -1492
rect 128394 40294 128450 40350
rect 128518 40294 128574 40350
rect 128642 40294 128698 40350
rect 128766 40294 128822 40350
rect 128394 40170 128450 40226
rect 128518 40170 128574 40226
rect 128642 40170 128698 40226
rect 128766 40170 128822 40226
rect 128394 40046 128450 40102
rect 128518 40046 128574 40102
rect 128642 40046 128698 40102
rect 128766 40046 128822 40102
rect 128394 39922 128450 39978
rect 128518 39922 128574 39978
rect 128642 39922 128698 39978
rect 128766 39922 128822 39978
rect 128394 22294 128450 22350
rect 128518 22294 128574 22350
rect 128642 22294 128698 22350
rect 128766 22294 128822 22350
rect 128394 22170 128450 22226
rect 128518 22170 128574 22226
rect 128642 22170 128698 22226
rect 128766 22170 128822 22226
rect 128394 22046 128450 22102
rect 128518 22046 128574 22102
rect 128642 22046 128698 22102
rect 128766 22046 128822 22102
rect 128394 21922 128450 21978
rect 128518 21922 128574 21978
rect 128642 21922 128698 21978
rect 128766 21922 128822 21978
rect 128394 4294 128450 4350
rect 128518 4294 128574 4350
rect 128642 4294 128698 4350
rect 128766 4294 128822 4350
rect 128394 4170 128450 4226
rect 128518 4170 128574 4226
rect 128642 4170 128698 4226
rect 128766 4170 128822 4226
rect 128394 4046 128450 4102
rect 128518 4046 128574 4102
rect 128642 4046 128698 4102
rect 128766 4046 128822 4102
rect 128394 3922 128450 3978
rect 128518 3922 128574 3978
rect 128642 3922 128698 3978
rect 128766 3922 128822 3978
rect 128394 -216 128450 -160
rect 128518 -216 128574 -160
rect 128642 -216 128698 -160
rect 128766 -216 128822 -160
rect 128394 -340 128450 -284
rect 128518 -340 128574 -284
rect 128642 -340 128698 -284
rect 128766 -340 128822 -284
rect 128394 -464 128450 -408
rect 128518 -464 128574 -408
rect 128642 -464 128698 -408
rect 128766 -464 128822 -408
rect 128394 -588 128450 -532
rect 128518 -588 128574 -532
rect 128642 -588 128698 -532
rect 128766 -588 128822 -532
rect 132114 46294 132170 46350
rect 132238 46294 132294 46350
rect 132362 46294 132418 46350
rect 132486 46294 132542 46350
rect 132114 46170 132170 46226
rect 132238 46170 132294 46226
rect 132362 46170 132418 46226
rect 132486 46170 132542 46226
rect 132114 46046 132170 46102
rect 132238 46046 132294 46102
rect 132362 46046 132418 46102
rect 132486 46046 132542 46102
rect 132114 45922 132170 45978
rect 132238 45922 132294 45978
rect 132362 45922 132418 45978
rect 132486 45922 132542 45978
rect 132114 28294 132170 28350
rect 132238 28294 132294 28350
rect 132362 28294 132418 28350
rect 132486 28294 132542 28350
rect 132114 28170 132170 28226
rect 132238 28170 132294 28226
rect 132362 28170 132418 28226
rect 132486 28170 132542 28226
rect 132114 28046 132170 28102
rect 132238 28046 132294 28102
rect 132362 28046 132418 28102
rect 132486 28046 132542 28102
rect 132114 27922 132170 27978
rect 132238 27922 132294 27978
rect 132362 27922 132418 27978
rect 132486 27922 132542 27978
rect 132114 10294 132170 10350
rect 132238 10294 132294 10350
rect 132362 10294 132418 10350
rect 132486 10294 132542 10350
rect 132114 10170 132170 10226
rect 132238 10170 132294 10226
rect 132362 10170 132418 10226
rect 132486 10170 132542 10226
rect 132114 10046 132170 10102
rect 132238 10046 132294 10102
rect 132362 10046 132418 10102
rect 132486 10046 132542 10102
rect 132114 9922 132170 9978
rect 132238 9922 132294 9978
rect 132362 9922 132418 9978
rect 132486 9922 132542 9978
rect 132114 -1176 132170 -1120
rect 132238 -1176 132294 -1120
rect 132362 -1176 132418 -1120
rect 132486 -1176 132542 -1120
rect 132114 -1300 132170 -1244
rect 132238 -1300 132294 -1244
rect 132362 -1300 132418 -1244
rect 132486 -1300 132542 -1244
rect 132114 -1424 132170 -1368
rect 132238 -1424 132294 -1368
rect 132362 -1424 132418 -1368
rect 132486 -1424 132542 -1368
rect 132114 -1548 132170 -1492
rect 132238 -1548 132294 -1492
rect 132362 -1548 132418 -1492
rect 132486 -1548 132542 -1492
rect 159114 40294 159170 40350
rect 159238 40294 159294 40350
rect 159362 40294 159418 40350
rect 159486 40294 159542 40350
rect 159114 40170 159170 40226
rect 159238 40170 159294 40226
rect 159362 40170 159418 40226
rect 159486 40170 159542 40226
rect 159114 40046 159170 40102
rect 159238 40046 159294 40102
rect 159362 40046 159418 40102
rect 159486 40046 159542 40102
rect 159114 39922 159170 39978
rect 159238 39922 159294 39978
rect 159362 39922 159418 39978
rect 159486 39922 159542 39978
rect 159114 22294 159170 22350
rect 159238 22294 159294 22350
rect 159362 22294 159418 22350
rect 159486 22294 159542 22350
rect 159114 22170 159170 22226
rect 159238 22170 159294 22226
rect 159362 22170 159418 22226
rect 159486 22170 159542 22226
rect 159114 22046 159170 22102
rect 159238 22046 159294 22102
rect 159362 22046 159418 22102
rect 159486 22046 159542 22102
rect 159114 21922 159170 21978
rect 159238 21922 159294 21978
rect 159362 21922 159418 21978
rect 159486 21922 159542 21978
rect 159114 4294 159170 4350
rect 159238 4294 159294 4350
rect 159362 4294 159418 4350
rect 159486 4294 159542 4350
rect 159114 4170 159170 4226
rect 159238 4170 159294 4226
rect 159362 4170 159418 4226
rect 159486 4170 159542 4226
rect 159114 4046 159170 4102
rect 159238 4046 159294 4102
rect 159362 4046 159418 4102
rect 159486 4046 159542 4102
rect 159114 3922 159170 3978
rect 159238 3922 159294 3978
rect 159362 3922 159418 3978
rect 159486 3922 159542 3978
rect 159114 -216 159170 -160
rect 159238 -216 159294 -160
rect 159362 -216 159418 -160
rect 159486 -216 159542 -160
rect 159114 -340 159170 -284
rect 159238 -340 159294 -284
rect 159362 -340 159418 -284
rect 159486 -340 159542 -284
rect 159114 -464 159170 -408
rect 159238 -464 159294 -408
rect 159362 -464 159418 -408
rect 159486 -464 159542 -408
rect 159114 -588 159170 -532
rect 159238 -588 159294 -532
rect 159362 -588 159418 -532
rect 159486 -588 159542 -532
rect 162834 46294 162890 46350
rect 162958 46294 163014 46350
rect 163082 46294 163138 46350
rect 163206 46294 163262 46350
rect 162834 46170 162890 46226
rect 162958 46170 163014 46226
rect 163082 46170 163138 46226
rect 163206 46170 163262 46226
rect 162834 46046 162890 46102
rect 162958 46046 163014 46102
rect 163082 46046 163138 46102
rect 163206 46046 163262 46102
rect 162834 45922 162890 45978
rect 162958 45922 163014 45978
rect 163082 45922 163138 45978
rect 163206 45922 163262 45978
rect 162834 28294 162890 28350
rect 162958 28294 163014 28350
rect 163082 28294 163138 28350
rect 163206 28294 163262 28350
rect 162834 28170 162890 28226
rect 162958 28170 163014 28226
rect 163082 28170 163138 28226
rect 163206 28170 163262 28226
rect 162834 28046 162890 28102
rect 162958 28046 163014 28102
rect 163082 28046 163138 28102
rect 163206 28046 163262 28102
rect 162834 27922 162890 27978
rect 162958 27922 163014 27978
rect 163082 27922 163138 27978
rect 163206 27922 163262 27978
rect 162834 10294 162890 10350
rect 162958 10294 163014 10350
rect 163082 10294 163138 10350
rect 163206 10294 163262 10350
rect 162834 10170 162890 10226
rect 162958 10170 163014 10226
rect 163082 10170 163138 10226
rect 163206 10170 163262 10226
rect 162834 10046 162890 10102
rect 162958 10046 163014 10102
rect 163082 10046 163138 10102
rect 163206 10046 163262 10102
rect 162834 9922 162890 9978
rect 162958 9922 163014 9978
rect 163082 9922 163138 9978
rect 163206 9922 163262 9978
rect 162834 -1176 162890 -1120
rect 162958 -1176 163014 -1120
rect 163082 -1176 163138 -1120
rect 163206 -1176 163262 -1120
rect 162834 -1300 162890 -1244
rect 162958 -1300 163014 -1244
rect 163082 -1300 163138 -1244
rect 163206 -1300 163262 -1244
rect 162834 -1424 162890 -1368
rect 162958 -1424 163014 -1368
rect 163082 -1424 163138 -1368
rect 163206 -1424 163262 -1368
rect 162834 -1548 162890 -1492
rect 162958 -1548 163014 -1492
rect 163082 -1548 163138 -1492
rect 163206 -1548 163262 -1492
rect 189834 40294 189890 40350
rect 189958 40294 190014 40350
rect 190082 40294 190138 40350
rect 190206 40294 190262 40350
rect 189834 40170 189890 40226
rect 189958 40170 190014 40226
rect 190082 40170 190138 40226
rect 190206 40170 190262 40226
rect 189834 40046 189890 40102
rect 189958 40046 190014 40102
rect 190082 40046 190138 40102
rect 190206 40046 190262 40102
rect 189834 39922 189890 39978
rect 189958 39922 190014 39978
rect 190082 39922 190138 39978
rect 190206 39922 190262 39978
rect 189834 22294 189890 22350
rect 189958 22294 190014 22350
rect 190082 22294 190138 22350
rect 190206 22294 190262 22350
rect 189834 22170 189890 22226
rect 189958 22170 190014 22226
rect 190082 22170 190138 22226
rect 190206 22170 190262 22226
rect 189834 22046 189890 22102
rect 189958 22046 190014 22102
rect 190082 22046 190138 22102
rect 190206 22046 190262 22102
rect 189834 21922 189890 21978
rect 189958 21922 190014 21978
rect 190082 21922 190138 21978
rect 190206 21922 190262 21978
rect 189834 4294 189890 4350
rect 189958 4294 190014 4350
rect 190082 4294 190138 4350
rect 190206 4294 190262 4350
rect 189834 4170 189890 4226
rect 189958 4170 190014 4226
rect 190082 4170 190138 4226
rect 190206 4170 190262 4226
rect 189834 4046 189890 4102
rect 189958 4046 190014 4102
rect 190082 4046 190138 4102
rect 190206 4046 190262 4102
rect 189834 3922 189890 3978
rect 189958 3922 190014 3978
rect 190082 3922 190138 3978
rect 190206 3922 190262 3978
rect 189834 -216 189890 -160
rect 189958 -216 190014 -160
rect 190082 -216 190138 -160
rect 190206 -216 190262 -160
rect 189834 -340 189890 -284
rect 189958 -340 190014 -284
rect 190082 -340 190138 -284
rect 190206 -340 190262 -284
rect 189834 -464 189890 -408
rect 189958 -464 190014 -408
rect 190082 -464 190138 -408
rect 190206 -464 190262 -408
rect 189834 -588 189890 -532
rect 189958 -588 190014 -532
rect 190082 -588 190138 -532
rect 190206 -588 190262 -532
rect 193554 46294 193610 46350
rect 193678 46294 193734 46350
rect 193802 46294 193858 46350
rect 193926 46294 193982 46350
rect 193554 46170 193610 46226
rect 193678 46170 193734 46226
rect 193802 46170 193858 46226
rect 193926 46170 193982 46226
rect 193554 46046 193610 46102
rect 193678 46046 193734 46102
rect 193802 46046 193858 46102
rect 193926 46046 193982 46102
rect 193554 45922 193610 45978
rect 193678 45922 193734 45978
rect 193802 45922 193858 45978
rect 193926 45922 193982 45978
rect 193554 28294 193610 28350
rect 193678 28294 193734 28350
rect 193802 28294 193858 28350
rect 193926 28294 193982 28350
rect 193554 28170 193610 28226
rect 193678 28170 193734 28226
rect 193802 28170 193858 28226
rect 193926 28170 193982 28226
rect 193554 28046 193610 28102
rect 193678 28046 193734 28102
rect 193802 28046 193858 28102
rect 193926 28046 193982 28102
rect 193554 27922 193610 27978
rect 193678 27922 193734 27978
rect 193802 27922 193858 27978
rect 193926 27922 193982 27978
rect 193554 10294 193610 10350
rect 193678 10294 193734 10350
rect 193802 10294 193858 10350
rect 193926 10294 193982 10350
rect 193554 10170 193610 10226
rect 193678 10170 193734 10226
rect 193802 10170 193858 10226
rect 193926 10170 193982 10226
rect 193554 10046 193610 10102
rect 193678 10046 193734 10102
rect 193802 10046 193858 10102
rect 193926 10046 193982 10102
rect 193554 9922 193610 9978
rect 193678 9922 193734 9978
rect 193802 9922 193858 9978
rect 193926 9922 193982 9978
rect 193554 -1176 193610 -1120
rect 193678 -1176 193734 -1120
rect 193802 -1176 193858 -1120
rect 193926 -1176 193982 -1120
rect 193554 -1300 193610 -1244
rect 193678 -1300 193734 -1244
rect 193802 -1300 193858 -1244
rect 193926 -1300 193982 -1244
rect 193554 -1424 193610 -1368
rect 193678 -1424 193734 -1368
rect 193802 -1424 193858 -1368
rect 193926 -1424 193982 -1368
rect 193554 -1548 193610 -1492
rect 193678 -1548 193734 -1492
rect 193802 -1548 193858 -1492
rect 193926 -1548 193982 -1492
rect 220554 40294 220610 40350
rect 220678 40294 220734 40350
rect 220802 40294 220858 40350
rect 220926 40294 220982 40350
rect 220554 40170 220610 40226
rect 220678 40170 220734 40226
rect 220802 40170 220858 40226
rect 220926 40170 220982 40226
rect 220554 40046 220610 40102
rect 220678 40046 220734 40102
rect 220802 40046 220858 40102
rect 220926 40046 220982 40102
rect 220554 39922 220610 39978
rect 220678 39922 220734 39978
rect 220802 39922 220858 39978
rect 220926 39922 220982 39978
rect 220554 22294 220610 22350
rect 220678 22294 220734 22350
rect 220802 22294 220858 22350
rect 220926 22294 220982 22350
rect 220554 22170 220610 22226
rect 220678 22170 220734 22226
rect 220802 22170 220858 22226
rect 220926 22170 220982 22226
rect 220554 22046 220610 22102
rect 220678 22046 220734 22102
rect 220802 22046 220858 22102
rect 220926 22046 220982 22102
rect 220554 21922 220610 21978
rect 220678 21922 220734 21978
rect 220802 21922 220858 21978
rect 220926 21922 220982 21978
rect 220554 4294 220610 4350
rect 220678 4294 220734 4350
rect 220802 4294 220858 4350
rect 220926 4294 220982 4350
rect 220554 4170 220610 4226
rect 220678 4170 220734 4226
rect 220802 4170 220858 4226
rect 220926 4170 220982 4226
rect 220554 4046 220610 4102
rect 220678 4046 220734 4102
rect 220802 4046 220858 4102
rect 220926 4046 220982 4102
rect 220554 3922 220610 3978
rect 220678 3922 220734 3978
rect 220802 3922 220858 3978
rect 220926 3922 220982 3978
rect 220554 -216 220610 -160
rect 220678 -216 220734 -160
rect 220802 -216 220858 -160
rect 220926 -216 220982 -160
rect 220554 -340 220610 -284
rect 220678 -340 220734 -284
rect 220802 -340 220858 -284
rect 220926 -340 220982 -284
rect 220554 -464 220610 -408
rect 220678 -464 220734 -408
rect 220802 -464 220858 -408
rect 220926 -464 220982 -408
rect 220554 -588 220610 -532
rect 220678 -588 220734 -532
rect 220802 -588 220858 -532
rect 220926 -588 220982 -532
rect 224274 46294 224330 46350
rect 224398 46294 224454 46350
rect 224522 46294 224578 46350
rect 224646 46294 224702 46350
rect 224274 46170 224330 46226
rect 224398 46170 224454 46226
rect 224522 46170 224578 46226
rect 224646 46170 224702 46226
rect 224274 46046 224330 46102
rect 224398 46046 224454 46102
rect 224522 46046 224578 46102
rect 224646 46046 224702 46102
rect 224274 45922 224330 45978
rect 224398 45922 224454 45978
rect 224522 45922 224578 45978
rect 224646 45922 224702 45978
rect 224274 28294 224330 28350
rect 224398 28294 224454 28350
rect 224522 28294 224578 28350
rect 224646 28294 224702 28350
rect 224274 28170 224330 28226
rect 224398 28170 224454 28226
rect 224522 28170 224578 28226
rect 224646 28170 224702 28226
rect 224274 28046 224330 28102
rect 224398 28046 224454 28102
rect 224522 28046 224578 28102
rect 224646 28046 224702 28102
rect 224274 27922 224330 27978
rect 224398 27922 224454 27978
rect 224522 27922 224578 27978
rect 224646 27922 224702 27978
rect 224274 10294 224330 10350
rect 224398 10294 224454 10350
rect 224522 10294 224578 10350
rect 224646 10294 224702 10350
rect 224274 10170 224330 10226
rect 224398 10170 224454 10226
rect 224522 10170 224578 10226
rect 224646 10170 224702 10226
rect 224274 10046 224330 10102
rect 224398 10046 224454 10102
rect 224522 10046 224578 10102
rect 224646 10046 224702 10102
rect 224274 9922 224330 9978
rect 224398 9922 224454 9978
rect 224522 9922 224578 9978
rect 224646 9922 224702 9978
rect 224274 -1176 224330 -1120
rect 224398 -1176 224454 -1120
rect 224522 -1176 224578 -1120
rect 224646 -1176 224702 -1120
rect 224274 -1300 224330 -1244
rect 224398 -1300 224454 -1244
rect 224522 -1300 224578 -1244
rect 224646 -1300 224702 -1244
rect 224274 -1424 224330 -1368
rect 224398 -1424 224454 -1368
rect 224522 -1424 224578 -1368
rect 224646 -1424 224702 -1368
rect 224274 -1548 224330 -1492
rect 224398 -1548 224454 -1492
rect 224522 -1548 224578 -1492
rect 224646 -1548 224702 -1492
rect 251274 40294 251330 40350
rect 251398 40294 251454 40350
rect 251522 40294 251578 40350
rect 251646 40294 251702 40350
rect 251274 40170 251330 40226
rect 251398 40170 251454 40226
rect 251522 40170 251578 40226
rect 251646 40170 251702 40226
rect 251274 40046 251330 40102
rect 251398 40046 251454 40102
rect 251522 40046 251578 40102
rect 251646 40046 251702 40102
rect 251274 39922 251330 39978
rect 251398 39922 251454 39978
rect 251522 39922 251578 39978
rect 251646 39922 251702 39978
rect 251274 22294 251330 22350
rect 251398 22294 251454 22350
rect 251522 22294 251578 22350
rect 251646 22294 251702 22350
rect 251274 22170 251330 22226
rect 251398 22170 251454 22226
rect 251522 22170 251578 22226
rect 251646 22170 251702 22226
rect 251274 22046 251330 22102
rect 251398 22046 251454 22102
rect 251522 22046 251578 22102
rect 251646 22046 251702 22102
rect 251274 21922 251330 21978
rect 251398 21922 251454 21978
rect 251522 21922 251578 21978
rect 251646 21922 251702 21978
rect 251274 4294 251330 4350
rect 251398 4294 251454 4350
rect 251522 4294 251578 4350
rect 251646 4294 251702 4350
rect 251274 4170 251330 4226
rect 251398 4170 251454 4226
rect 251522 4170 251578 4226
rect 251646 4170 251702 4226
rect 251274 4046 251330 4102
rect 251398 4046 251454 4102
rect 251522 4046 251578 4102
rect 251646 4046 251702 4102
rect 251274 3922 251330 3978
rect 251398 3922 251454 3978
rect 251522 3922 251578 3978
rect 251646 3922 251702 3978
rect 251274 -216 251330 -160
rect 251398 -216 251454 -160
rect 251522 -216 251578 -160
rect 251646 -216 251702 -160
rect 251274 -340 251330 -284
rect 251398 -340 251454 -284
rect 251522 -340 251578 -284
rect 251646 -340 251702 -284
rect 251274 -464 251330 -408
rect 251398 -464 251454 -408
rect 251522 -464 251578 -408
rect 251646 -464 251702 -408
rect 251274 -588 251330 -532
rect 251398 -588 251454 -532
rect 251522 -588 251578 -532
rect 251646 -588 251702 -532
rect 268716 246122 268772 246178
rect 281994 256294 282050 256350
rect 282118 256294 282174 256350
rect 282242 256294 282298 256350
rect 282366 256294 282422 256350
rect 270508 252782 270564 252838
rect 269612 252422 269668 252478
rect 269500 252062 269556 252118
rect 254994 46294 255050 46350
rect 255118 46294 255174 46350
rect 255242 46294 255298 46350
rect 255366 46294 255422 46350
rect 254994 46170 255050 46226
rect 255118 46170 255174 46226
rect 255242 46170 255298 46226
rect 255366 46170 255422 46226
rect 254994 46046 255050 46102
rect 255118 46046 255174 46102
rect 255242 46046 255298 46102
rect 255366 46046 255422 46102
rect 254994 45922 255050 45978
rect 255118 45922 255174 45978
rect 255242 45922 255298 45978
rect 255366 45922 255422 45978
rect 281994 256170 282050 256226
rect 282118 256170 282174 256226
rect 282242 256170 282298 256226
rect 282366 256170 282422 256226
rect 281994 256046 282050 256102
rect 282118 256046 282174 256102
rect 282242 256046 282298 256102
rect 282366 256046 282422 256102
rect 281994 255922 282050 255978
rect 282118 255922 282174 255978
rect 282242 255922 282298 255978
rect 282366 255922 282422 255978
rect 275548 252602 275604 252658
rect 274652 249362 274708 249418
rect 273756 152882 273812 152938
rect 275660 252242 275716 252298
rect 281994 238294 282050 238350
rect 282118 238294 282174 238350
rect 282242 238294 282298 238350
rect 282366 238294 282422 238350
rect 281994 238170 282050 238226
rect 282118 238170 282174 238226
rect 282242 238170 282298 238226
rect 282366 238170 282422 238226
rect 281994 238046 282050 238102
rect 282118 238046 282174 238102
rect 282242 238046 282298 238102
rect 282366 238046 282422 238102
rect 281994 237922 282050 237978
rect 282118 237922 282174 237978
rect 282242 237922 282298 237978
rect 282366 237922 282422 237978
rect 281994 220294 282050 220350
rect 282118 220294 282174 220350
rect 282242 220294 282298 220350
rect 282366 220294 282422 220350
rect 281994 220170 282050 220226
rect 282118 220170 282174 220226
rect 282242 220170 282298 220226
rect 282366 220170 282422 220226
rect 281994 220046 282050 220102
rect 282118 220046 282174 220102
rect 282242 220046 282298 220102
rect 282366 220046 282422 220102
rect 281994 219922 282050 219978
rect 282118 219922 282174 219978
rect 282242 219922 282298 219978
rect 282366 219922 282422 219978
rect 281994 202294 282050 202350
rect 282118 202294 282174 202350
rect 282242 202294 282298 202350
rect 282366 202294 282422 202350
rect 281994 202170 282050 202226
rect 282118 202170 282174 202226
rect 282242 202170 282298 202226
rect 282366 202170 282422 202226
rect 281994 202046 282050 202102
rect 282118 202046 282174 202102
rect 282242 202046 282298 202102
rect 282366 202046 282422 202102
rect 281994 201922 282050 201978
rect 282118 201922 282174 201978
rect 282242 201922 282298 201978
rect 282366 201922 282422 201978
rect 281994 184294 282050 184350
rect 282118 184294 282174 184350
rect 282242 184294 282298 184350
rect 282366 184294 282422 184350
rect 281994 184170 282050 184226
rect 282118 184170 282174 184226
rect 282242 184170 282298 184226
rect 282366 184170 282422 184226
rect 281994 184046 282050 184102
rect 282118 184046 282174 184102
rect 282242 184046 282298 184102
rect 282366 184046 282422 184102
rect 281994 183922 282050 183978
rect 282118 183922 282174 183978
rect 282242 183922 282298 183978
rect 282366 183922 282422 183978
rect 281994 166294 282050 166350
rect 282118 166294 282174 166350
rect 282242 166294 282298 166350
rect 282366 166294 282422 166350
rect 281994 166170 282050 166226
rect 282118 166170 282174 166226
rect 282242 166170 282298 166226
rect 282366 166170 282422 166226
rect 281994 166046 282050 166102
rect 282118 166046 282174 166102
rect 282242 166046 282298 166102
rect 282366 166046 282422 166102
rect 281994 165922 282050 165978
rect 282118 165922 282174 165978
rect 282242 165922 282298 165978
rect 282366 165922 282422 165978
rect 281994 148294 282050 148350
rect 282118 148294 282174 148350
rect 282242 148294 282298 148350
rect 282366 148294 282422 148350
rect 281994 148170 282050 148226
rect 282118 148170 282174 148226
rect 282242 148170 282298 148226
rect 282366 148170 282422 148226
rect 281994 148046 282050 148102
rect 282118 148046 282174 148102
rect 282242 148046 282298 148102
rect 282366 148046 282422 148102
rect 281994 147922 282050 147978
rect 282118 147922 282174 147978
rect 282242 147922 282298 147978
rect 282366 147922 282422 147978
rect 281994 130294 282050 130350
rect 282118 130294 282174 130350
rect 282242 130294 282298 130350
rect 282366 130294 282422 130350
rect 281994 130170 282050 130226
rect 282118 130170 282174 130226
rect 282242 130170 282298 130226
rect 282366 130170 282422 130226
rect 281994 130046 282050 130102
rect 282118 130046 282174 130102
rect 282242 130046 282298 130102
rect 282366 130046 282422 130102
rect 281994 129922 282050 129978
rect 282118 129922 282174 129978
rect 282242 129922 282298 129978
rect 282366 129922 282422 129978
rect 281994 112294 282050 112350
rect 282118 112294 282174 112350
rect 282242 112294 282298 112350
rect 282366 112294 282422 112350
rect 281994 112170 282050 112226
rect 282118 112170 282174 112226
rect 282242 112170 282298 112226
rect 282366 112170 282422 112226
rect 281994 112046 282050 112102
rect 282118 112046 282174 112102
rect 282242 112046 282298 112102
rect 282366 112046 282422 112102
rect 281994 111922 282050 111978
rect 282118 111922 282174 111978
rect 282242 111922 282298 111978
rect 282366 111922 282422 111978
rect 281994 94294 282050 94350
rect 282118 94294 282174 94350
rect 282242 94294 282298 94350
rect 282366 94294 282422 94350
rect 281994 94170 282050 94226
rect 282118 94170 282174 94226
rect 282242 94170 282298 94226
rect 282366 94170 282422 94226
rect 281994 94046 282050 94102
rect 282118 94046 282174 94102
rect 282242 94046 282298 94102
rect 282366 94046 282422 94102
rect 281994 93922 282050 93978
rect 282118 93922 282174 93978
rect 282242 93922 282298 93978
rect 282366 93922 282422 93978
rect 281994 76294 282050 76350
rect 282118 76294 282174 76350
rect 282242 76294 282298 76350
rect 282366 76294 282422 76350
rect 281994 76170 282050 76226
rect 282118 76170 282174 76226
rect 282242 76170 282298 76226
rect 282366 76170 282422 76226
rect 281994 76046 282050 76102
rect 282118 76046 282174 76102
rect 282242 76046 282298 76102
rect 282366 76046 282422 76102
rect 281994 75922 282050 75978
rect 282118 75922 282174 75978
rect 282242 75922 282298 75978
rect 282366 75922 282422 75978
rect 281994 58294 282050 58350
rect 282118 58294 282174 58350
rect 282242 58294 282298 58350
rect 282366 58294 282422 58350
rect 281994 58170 282050 58226
rect 282118 58170 282174 58226
rect 282242 58170 282298 58226
rect 282366 58170 282422 58226
rect 281994 58046 282050 58102
rect 282118 58046 282174 58102
rect 282242 58046 282298 58102
rect 282366 58046 282422 58102
rect 281994 57922 282050 57978
rect 282118 57922 282174 57978
rect 282242 57922 282298 57978
rect 282366 57922 282422 57978
rect 281994 40294 282050 40350
rect 282118 40294 282174 40350
rect 282242 40294 282298 40350
rect 282366 40294 282422 40350
rect 281994 40170 282050 40226
rect 282118 40170 282174 40226
rect 282242 40170 282298 40226
rect 282366 40170 282422 40226
rect 281994 40046 282050 40102
rect 282118 40046 282174 40102
rect 282242 40046 282298 40102
rect 282366 40046 282422 40102
rect 281994 39922 282050 39978
rect 282118 39922 282174 39978
rect 282242 39922 282298 39978
rect 282366 39922 282422 39978
rect 254994 28294 255050 28350
rect 255118 28294 255174 28350
rect 255242 28294 255298 28350
rect 255366 28294 255422 28350
rect 254994 28170 255050 28226
rect 255118 28170 255174 28226
rect 255242 28170 255298 28226
rect 255366 28170 255422 28226
rect 254994 28046 255050 28102
rect 255118 28046 255174 28102
rect 255242 28046 255298 28102
rect 255366 28046 255422 28102
rect 254994 27922 255050 27978
rect 255118 27922 255174 27978
rect 255242 27922 255298 27978
rect 255366 27922 255422 27978
rect 254994 10294 255050 10350
rect 255118 10294 255174 10350
rect 255242 10294 255298 10350
rect 255366 10294 255422 10350
rect 254994 10170 255050 10226
rect 255118 10170 255174 10226
rect 255242 10170 255298 10226
rect 255366 10170 255422 10226
rect 254994 10046 255050 10102
rect 255118 10046 255174 10102
rect 255242 10046 255298 10102
rect 255366 10046 255422 10102
rect 254994 9922 255050 9978
rect 255118 9922 255174 9978
rect 255242 9922 255298 9978
rect 255366 9922 255422 9978
rect 254994 -1176 255050 -1120
rect 255118 -1176 255174 -1120
rect 255242 -1176 255298 -1120
rect 255366 -1176 255422 -1120
rect 254994 -1300 255050 -1244
rect 255118 -1300 255174 -1244
rect 255242 -1300 255298 -1244
rect 255366 -1300 255422 -1244
rect 254994 -1424 255050 -1368
rect 255118 -1424 255174 -1368
rect 255242 -1424 255298 -1368
rect 255366 -1424 255422 -1368
rect 254994 -1548 255050 -1492
rect 255118 -1548 255174 -1492
rect 255242 -1548 255298 -1492
rect 255366 -1548 255422 -1492
rect 281994 22294 282050 22350
rect 282118 22294 282174 22350
rect 282242 22294 282298 22350
rect 282366 22294 282422 22350
rect 281994 22170 282050 22226
rect 282118 22170 282174 22226
rect 282242 22170 282298 22226
rect 282366 22170 282422 22226
rect 281994 22046 282050 22102
rect 282118 22046 282174 22102
rect 282242 22046 282298 22102
rect 282366 22046 282422 22102
rect 281994 21922 282050 21978
rect 282118 21922 282174 21978
rect 282242 21922 282298 21978
rect 282366 21922 282422 21978
rect 281994 4294 282050 4350
rect 282118 4294 282174 4350
rect 282242 4294 282298 4350
rect 282366 4294 282422 4350
rect 281994 4170 282050 4226
rect 282118 4170 282174 4226
rect 282242 4170 282298 4226
rect 282366 4170 282422 4226
rect 281994 4046 282050 4102
rect 282118 4046 282174 4102
rect 282242 4046 282298 4102
rect 282366 4046 282422 4102
rect 281994 3922 282050 3978
rect 282118 3922 282174 3978
rect 282242 3922 282298 3978
rect 282366 3922 282422 3978
rect 281994 -216 282050 -160
rect 282118 -216 282174 -160
rect 282242 -216 282298 -160
rect 282366 -216 282422 -160
rect 281994 -340 282050 -284
rect 282118 -340 282174 -284
rect 282242 -340 282298 -284
rect 282366 -340 282422 -284
rect 281994 -464 282050 -408
rect 282118 -464 282174 -408
rect 282242 -464 282298 -408
rect 282366 -464 282422 -408
rect 281994 -588 282050 -532
rect 282118 -588 282174 -532
rect 282242 -588 282298 -532
rect 282366 -588 282422 -532
rect 312714 256294 312770 256350
rect 312838 256294 312894 256350
rect 312962 256294 313018 256350
rect 313086 256294 313142 256350
rect 312714 256170 312770 256226
rect 312838 256170 312894 256226
rect 312962 256170 313018 256226
rect 313086 256170 313142 256226
rect 312714 256046 312770 256102
rect 312838 256046 312894 256102
rect 312962 256046 313018 256102
rect 313086 256046 313142 256102
rect 312714 255922 312770 255978
rect 312838 255922 312894 255978
rect 312962 255922 313018 255978
rect 313086 255922 313142 255978
rect 285714 244294 285770 244350
rect 285838 244294 285894 244350
rect 285962 244294 286018 244350
rect 286086 244294 286142 244350
rect 285714 244170 285770 244226
rect 285838 244170 285894 244226
rect 285962 244170 286018 244226
rect 286086 244170 286142 244226
rect 285714 244046 285770 244102
rect 285838 244046 285894 244102
rect 285962 244046 286018 244102
rect 286086 244046 286142 244102
rect 285714 243922 285770 243978
rect 285838 243922 285894 243978
rect 285962 243922 286018 243978
rect 286086 243922 286142 243978
rect 285714 226294 285770 226350
rect 285838 226294 285894 226350
rect 285962 226294 286018 226350
rect 286086 226294 286142 226350
rect 285714 226170 285770 226226
rect 285838 226170 285894 226226
rect 285962 226170 286018 226226
rect 286086 226170 286142 226226
rect 285714 226046 285770 226102
rect 285838 226046 285894 226102
rect 285962 226046 286018 226102
rect 286086 226046 286142 226102
rect 285714 225922 285770 225978
rect 285838 225922 285894 225978
rect 285962 225922 286018 225978
rect 286086 225922 286142 225978
rect 285714 208294 285770 208350
rect 285838 208294 285894 208350
rect 285962 208294 286018 208350
rect 286086 208294 286142 208350
rect 285714 208170 285770 208226
rect 285838 208170 285894 208226
rect 285962 208170 286018 208226
rect 286086 208170 286142 208226
rect 285714 208046 285770 208102
rect 285838 208046 285894 208102
rect 285962 208046 286018 208102
rect 286086 208046 286142 208102
rect 285714 207922 285770 207978
rect 285838 207922 285894 207978
rect 285962 207922 286018 207978
rect 286086 207922 286142 207978
rect 285714 190294 285770 190350
rect 285838 190294 285894 190350
rect 285962 190294 286018 190350
rect 286086 190294 286142 190350
rect 285714 190170 285770 190226
rect 285838 190170 285894 190226
rect 285962 190170 286018 190226
rect 286086 190170 286142 190226
rect 285714 190046 285770 190102
rect 285838 190046 285894 190102
rect 285962 190046 286018 190102
rect 286086 190046 286142 190102
rect 285714 189922 285770 189978
rect 285838 189922 285894 189978
rect 285962 189922 286018 189978
rect 286086 189922 286142 189978
rect 285714 172294 285770 172350
rect 285838 172294 285894 172350
rect 285962 172294 286018 172350
rect 286086 172294 286142 172350
rect 285714 172170 285770 172226
rect 285838 172170 285894 172226
rect 285962 172170 286018 172226
rect 286086 172170 286142 172226
rect 285714 172046 285770 172102
rect 285838 172046 285894 172102
rect 285962 172046 286018 172102
rect 286086 172046 286142 172102
rect 285714 171922 285770 171978
rect 285838 171922 285894 171978
rect 285962 171922 286018 171978
rect 286086 171922 286142 171978
rect 285714 154294 285770 154350
rect 285838 154294 285894 154350
rect 285962 154294 286018 154350
rect 286086 154294 286142 154350
rect 285714 154170 285770 154226
rect 285838 154170 285894 154226
rect 285962 154170 286018 154226
rect 286086 154170 286142 154226
rect 285714 154046 285770 154102
rect 285838 154046 285894 154102
rect 285962 154046 286018 154102
rect 286086 154046 286142 154102
rect 285714 153922 285770 153978
rect 285838 153922 285894 153978
rect 285962 153922 286018 153978
rect 286086 153922 286142 153978
rect 285714 136294 285770 136350
rect 285838 136294 285894 136350
rect 285962 136294 286018 136350
rect 286086 136294 286142 136350
rect 285714 136170 285770 136226
rect 285838 136170 285894 136226
rect 285962 136170 286018 136226
rect 286086 136170 286142 136226
rect 285714 136046 285770 136102
rect 285838 136046 285894 136102
rect 285962 136046 286018 136102
rect 286086 136046 286142 136102
rect 285714 135922 285770 135978
rect 285838 135922 285894 135978
rect 285962 135922 286018 135978
rect 286086 135922 286142 135978
rect 285714 118294 285770 118350
rect 285838 118294 285894 118350
rect 285962 118294 286018 118350
rect 286086 118294 286142 118350
rect 285714 118170 285770 118226
rect 285838 118170 285894 118226
rect 285962 118170 286018 118226
rect 286086 118170 286142 118226
rect 285714 118046 285770 118102
rect 285838 118046 285894 118102
rect 285962 118046 286018 118102
rect 286086 118046 286142 118102
rect 285714 117922 285770 117978
rect 285838 117922 285894 117978
rect 285962 117922 286018 117978
rect 286086 117922 286142 117978
rect 285714 100294 285770 100350
rect 285838 100294 285894 100350
rect 285962 100294 286018 100350
rect 286086 100294 286142 100350
rect 285714 100170 285770 100226
rect 285838 100170 285894 100226
rect 285962 100170 286018 100226
rect 286086 100170 286142 100226
rect 285714 100046 285770 100102
rect 285838 100046 285894 100102
rect 285962 100046 286018 100102
rect 286086 100046 286142 100102
rect 285714 99922 285770 99978
rect 285838 99922 285894 99978
rect 285962 99922 286018 99978
rect 286086 99922 286142 99978
rect 285714 82294 285770 82350
rect 285838 82294 285894 82350
rect 285962 82294 286018 82350
rect 286086 82294 286142 82350
rect 285714 82170 285770 82226
rect 285838 82170 285894 82226
rect 285962 82170 286018 82226
rect 286086 82170 286142 82226
rect 285714 82046 285770 82102
rect 285838 82046 285894 82102
rect 285962 82046 286018 82102
rect 286086 82046 286142 82102
rect 285714 81922 285770 81978
rect 285838 81922 285894 81978
rect 285962 81922 286018 81978
rect 286086 81922 286142 81978
rect 285714 64294 285770 64350
rect 285838 64294 285894 64350
rect 285962 64294 286018 64350
rect 286086 64294 286142 64350
rect 285714 64170 285770 64226
rect 285838 64170 285894 64226
rect 285962 64170 286018 64226
rect 286086 64170 286142 64226
rect 285714 64046 285770 64102
rect 285838 64046 285894 64102
rect 285962 64046 286018 64102
rect 286086 64046 286142 64102
rect 285714 63922 285770 63978
rect 285838 63922 285894 63978
rect 285962 63922 286018 63978
rect 286086 63922 286142 63978
rect 285714 46294 285770 46350
rect 285838 46294 285894 46350
rect 285962 46294 286018 46350
rect 286086 46294 286142 46350
rect 285714 46170 285770 46226
rect 285838 46170 285894 46226
rect 285962 46170 286018 46226
rect 286086 46170 286142 46226
rect 285714 46046 285770 46102
rect 285838 46046 285894 46102
rect 285962 46046 286018 46102
rect 286086 46046 286142 46102
rect 285714 45922 285770 45978
rect 285838 45922 285894 45978
rect 285962 45922 286018 45978
rect 286086 45922 286142 45978
rect 285714 28294 285770 28350
rect 285838 28294 285894 28350
rect 285962 28294 286018 28350
rect 286086 28294 286142 28350
rect 285714 28170 285770 28226
rect 285838 28170 285894 28226
rect 285962 28170 286018 28226
rect 286086 28170 286142 28226
rect 285714 28046 285770 28102
rect 285838 28046 285894 28102
rect 285962 28046 286018 28102
rect 286086 28046 286142 28102
rect 285714 27922 285770 27978
rect 285838 27922 285894 27978
rect 285962 27922 286018 27978
rect 286086 27922 286142 27978
rect 285714 10294 285770 10350
rect 285838 10294 285894 10350
rect 285962 10294 286018 10350
rect 286086 10294 286142 10350
rect 285714 10170 285770 10226
rect 285838 10170 285894 10226
rect 285962 10170 286018 10226
rect 286086 10170 286142 10226
rect 285714 10046 285770 10102
rect 285838 10046 285894 10102
rect 285962 10046 286018 10102
rect 286086 10046 286142 10102
rect 285714 9922 285770 9978
rect 285838 9922 285894 9978
rect 285962 9922 286018 9978
rect 286086 9922 286142 9978
rect 312714 238294 312770 238350
rect 312838 238294 312894 238350
rect 312962 238294 313018 238350
rect 313086 238294 313142 238350
rect 312714 238170 312770 238226
rect 312838 238170 312894 238226
rect 312962 238170 313018 238226
rect 313086 238170 313142 238226
rect 312714 238046 312770 238102
rect 312838 238046 312894 238102
rect 312962 238046 313018 238102
rect 313086 238046 313142 238102
rect 312714 237922 312770 237978
rect 312838 237922 312894 237978
rect 312962 237922 313018 237978
rect 313086 237922 313142 237978
rect 312714 220294 312770 220350
rect 312838 220294 312894 220350
rect 312962 220294 313018 220350
rect 313086 220294 313142 220350
rect 312714 220170 312770 220226
rect 312838 220170 312894 220226
rect 312962 220170 313018 220226
rect 313086 220170 313142 220226
rect 312714 220046 312770 220102
rect 312838 220046 312894 220102
rect 312962 220046 313018 220102
rect 313086 220046 313142 220102
rect 312714 219922 312770 219978
rect 312838 219922 312894 219978
rect 312962 219922 313018 219978
rect 313086 219922 313142 219978
rect 291564 211022 291620 211078
rect 296492 210842 296548 210898
rect 299528 82091 299584 82147
rect 299632 82091 299688 82147
rect 299736 82091 299792 82147
rect 299528 81987 299584 82043
rect 299632 81987 299688 82043
rect 299736 81987 299792 82043
rect 299528 81883 299584 81939
rect 299632 81883 299688 81939
rect 299736 81883 299792 81939
rect 295412 76294 295468 76350
rect 295536 76294 295592 76350
rect 295412 76170 295468 76226
rect 295536 76170 295592 76226
rect 295412 76046 295468 76102
rect 295536 76046 295592 76102
rect 295412 75922 295468 75978
rect 295536 75922 295592 75978
rect 303728 76294 303784 76350
rect 303852 76294 303908 76350
rect 303728 76170 303784 76226
rect 303852 76170 303908 76226
rect 303728 76046 303784 76102
rect 303852 76046 303908 76102
rect 303728 75922 303784 75978
rect 303852 75922 303908 75978
rect 299570 64294 299626 64350
rect 299694 64294 299750 64350
rect 299570 64170 299626 64226
rect 299694 64170 299750 64226
rect 299570 64046 299626 64102
rect 299694 64046 299750 64102
rect 299570 63922 299626 63978
rect 299694 63922 299750 63978
rect 295412 58294 295468 58350
rect 295536 58294 295592 58350
rect 295412 58170 295468 58226
rect 295536 58170 295592 58226
rect 295412 58046 295468 58102
rect 295536 58046 295592 58102
rect 295412 57922 295468 57978
rect 295536 57922 295592 57978
rect 303728 58294 303784 58350
rect 303852 58294 303908 58350
rect 303728 58170 303784 58226
rect 303852 58170 303908 58226
rect 303728 58046 303784 58102
rect 303852 58046 303908 58102
rect 303728 57922 303784 57978
rect 303852 57922 303908 57978
rect 316434 244294 316490 244350
rect 316558 244294 316614 244350
rect 316682 244294 316738 244350
rect 316806 244294 316862 244350
rect 316434 244170 316490 244226
rect 316558 244170 316614 244226
rect 316682 244170 316738 244226
rect 316806 244170 316862 244226
rect 316434 244046 316490 244102
rect 316558 244046 316614 244102
rect 316682 244046 316738 244102
rect 316806 244046 316862 244102
rect 316434 243922 316490 243978
rect 316558 243922 316614 243978
rect 316682 243922 316738 243978
rect 316806 243922 316862 243978
rect 316434 226294 316490 226350
rect 316558 226294 316614 226350
rect 316682 226294 316738 226350
rect 316806 226294 316862 226350
rect 316434 226170 316490 226226
rect 316558 226170 316614 226226
rect 316682 226170 316738 226226
rect 316806 226170 316862 226226
rect 316434 226046 316490 226102
rect 316558 226046 316614 226102
rect 316682 226046 316738 226102
rect 316806 226046 316862 226102
rect 316434 225922 316490 225978
rect 316558 225922 316614 225978
rect 316682 225922 316738 225978
rect 316806 225922 316862 225978
rect 312714 202294 312770 202350
rect 312838 202294 312894 202350
rect 312962 202294 313018 202350
rect 313086 202294 313142 202350
rect 312714 202170 312770 202226
rect 312838 202170 312894 202226
rect 312962 202170 313018 202226
rect 313086 202170 313142 202226
rect 312714 202046 312770 202102
rect 312838 202046 312894 202102
rect 312962 202046 313018 202102
rect 313086 202046 313142 202102
rect 312714 201922 312770 201978
rect 312838 201922 312894 201978
rect 312962 201922 313018 201978
rect 313086 201922 313142 201978
rect 312714 184294 312770 184350
rect 312838 184294 312894 184350
rect 312962 184294 313018 184350
rect 313086 184294 313142 184350
rect 312714 184170 312770 184226
rect 312838 184170 312894 184226
rect 312962 184170 313018 184226
rect 313086 184170 313142 184226
rect 312714 184046 312770 184102
rect 312838 184046 312894 184102
rect 312962 184046 313018 184102
rect 313086 184046 313142 184102
rect 312714 183922 312770 183978
rect 312838 183922 312894 183978
rect 312962 183922 313018 183978
rect 313086 183922 313142 183978
rect 312714 166294 312770 166350
rect 312838 166294 312894 166350
rect 312962 166294 313018 166350
rect 313086 166294 313142 166350
rect 312714 166170 312770 166226
rect 312838 166170 312894 166226
rect 312962 166170 313018 166226
rect 313086 166170 313142 166226
rect 312714 166046 312770 166102
rect 312838 166046 312894 166102
rect 312962 166046 313018 166102
rect 313086 166046 313142 166102
rect 312714 165922 312770 165978
rect 312838 165922 312894 165978
rect 312962 165922 313018 165978
rect 313086 165922 313142 165978
rect 312714 148294 312770 148350
rect 312838 148294 312894 148350
rect 312962 148294 313018 148350
rect 313086 148294 313142 148350
rect 312714 148170 312770 148226
rect 312838 148170 312894 148226
rect 312962 148170 313018 148226
rect 313086 148170 313142 148226
rect 312714 148046 312770 148102
rect 312838 148046 312894 148102
rect 312962 148046 313018 148102
rect 313086 148046 313142 148102
rect 312714 147922 312770 147978
rect 312838 147922 312894 147978
rect 312962 147922 313018 147978
rect 313086 147922 313142 147978
rect 312714 130294 312770 130350
rect 312838 130294 312894 130350
rect 312962 130294 313018 130350
rect 313086 130294 313142 130350
rect 312714 130170 312770 130226
rect 312838 130170 312894 130226
rect 312962 130170 313018 130226
rect 313086 130170 313142 130226
rect 312714 130046 312770 130102
rect 312838 130046 312894 130102
rect 312962 130046 313018 130102
rect 313086 130046 313142 130102
rect 312714 129922 312770 129978
rect 312838 129922 312894 129978
rect 312962 129922 313018 129978
rect 313086 129922 313142 129978
rect 313404 153602 313460 153658
rect 312714 112294 312770 112350
rect 312838 112294 312894 112350
rect 312962 112294 313018 112350
rect 313086 112294 313142 112350
rect 312714 112170 312770 112226
rect 312838 112170 312894 112226
rect 312962 112170 313018 112226
rect 313086 112170 313142 112226
rect 312714 112046 312770 112102
rect 312838 112046 312894 112102
rect 312962 112046 313018 112102
rect 313086 112046 313142 112102
rect 312714 111922 312770 111978
rect 312838 111922 312894 111978
rect 312962 111922 313018 111978
rect 313086 111922 313142 111978
rect 312714 94294 312770 94350
rect 312838 94294 312894 94350
rect 312962 94294 313018 94350
rect 313086 94294 313142 94350
rect 312714 94170 312770 94226
rect 312838 94170 312894 94226
rect 312962 94170 313018 94226
rect 313086 94170 313142 94226
rect 312714 94046 312770 94102
rect 312838 94046 312894 94102
rect 312962 94046 313018 94102
rect 313086 94046 313142 94102
rect 312714 93922 312770 93978
rect 312838 93922 312894 93978
rect 312962 93922 313018 93978
rect 313086 93922 313142 93978
rect 307844 82091 307900 82147
rect 307948 82091 308004 82147
rect 308052 82091 308108 82147
rect 307844 81987 307900 82043
rect 307948 81987 308004 82043
rect 308052 81987 308108 82043
rect 307844 81883 307900 81939
rect 307948 81883 308004 81939
rect 308052 81883 308108 81939
rect 312044 76294 312100 76350
rect 312168 76294 312224 76350
rect 312044 76170 312100 76226
rect 312168 76170 312224 76226
rect 312044 76046 312100 76102
rect 312168 76046 312224 76102
rect 312044 75922 312100 75978
rect 312168 75922 312224 75978
rect 312714 76294 312770 76350
rect 312838 76294 312894 76350
rect 312962 76294 313018 76350
rect 313086 76294 313142 76350
rect 312714 76170 312770 76226
rect 312838 76170 312894 76226
rect 312962 76170 313018 76226
rect 313086 76170 313142 76226
rect 312714 76046 312770 76102
rect 312838 76046 312894 76102
rect 312962 76046 313018 76102
rect 313086 76046 313142 76102
rect 312714 75922 312770 75978
rect 312838 75922 312894 75978
rect 312962 75922 313018 75978
rect 313086 75922 313142 75978
rect 307886 64294 307942 64350
rect 308010 64294 308066 64350
rect 307886 64170 307942 64226
rect 308010 64170 308066 64226
rect 307886 64046 307942 64102
rect 308010 64046 308066 64102
rect 307886 63922 307942 63978
rect 308010 63922 308066 63978
rect 312044 58294 312100 58350
rect 312168 58294 312224 58350
rect 312044 58170 312100 58226
rect 312168 58170 312224 58226
rect 312044 58046 312100 58102
rect 312168 58046 312224 58102
rect 312044 57922 312100 57978
rect 312168 57922 312224 57978
rect 312714 58294 312770 58350
rect 312838 58294 312894 58350
rect 312962 58294 313018 58350
rect 313086 58294 313142 58350
rect 312714 58170 312770 58226
rect 312838 58170 312894 58226
rect 312962 58170 313018 58226
rect 313086 58170 313142 58226
rect 312714 58046 312770 58102
rect 312838 58046 312894 58102
rect 312962 58046 313018 58102
rect 313086 58046 313142 58102
rect 312714 57922 312770 57978
rect 312838 57922 312894 57978
rect 312962 57922 313018 57978
rect 313086 57922 313142 57978
rect 343434 256294 343490 256350
rect 343558 256294 343614 256350
rect 343682 256294 343738 256350
rect 343806 256294 343862 256350
rect 343434 256170 343490 256226
rect 343558 256170 343614 256226
rect 343682 256170 343738 256226
rect 343806 256170 343862 256226
rect 343434 256046 343490 256102
rect 343558 256046 343614 256102
rect 343682 256046 343738 256102
rect 343806 256046 343862 256102
rect 343434 255922 343490 255978
rect 343558 255922 343614 255978
rect 343682 255922 343738 255978
rect 343806 255922 343862 255978
rect 343434 238294 343490 238350
rect 343558 238294 343614 238350
rect 343682 238294 343738 238350
rect 343806 238294 343862 238350
rect 343434 238170 343490 238226
rect 343558 238170 343614 238226
rect 343682 238170 343738 238226
rect 343806 238170 343862 238226
rect 343434 238046 343490 238102
rect 343558 238046 343614 238102
rect 343682 238046 343738 238102
rect 343806 238046 343862 238102
rect 343434 237922 343490 237978
rect 343558 237922 343614 237978
rect 343682 237922 343738 237978
rect 343806 237922 343862 237978
rect 343434 220294 343490 220350
rect 343558 220294 343614 220350
rect 343682 220294 343738 220350
rect 343806 220294 343862 220350
rect 343434 220170 343490 220226
rect 343558 220170 343614 220226
rect 343682 220170 343738 220226
rect 343806 220170 343862 220226
rect 343434 220046 343490 220102
rect 343558 220046 343614 220102
rect 343682 220046 343738 220102
rect 343806 220046 343862 220102
rect 343434 219922 343490 219978
rect 343558 219922 343614 219978
rect 343682 219922 343738 219978
rect 343806 219922 343862 219978
rect 316434 208294 316490 208350
rect 316558 208294 316614 208350
rect 316682 208294 316738 208350
rect 316806 208294 316862 208350
rect 316434 208170 316490 208226
rect 316558 208170 316614 208226
rect 316682 208170 316738 208226
rect 316806 208170 316862 208226
rect 316434 208046 316490 208102
rect 316558 208046 316614 208102
rect 316682 208046 316738 208102
rect 316806 208046 316862 208102
rect 316434 207922 316490 207978
rect 316558 207922 316614 207978
rect 316682 207922 316738 207978
rect 316806 207922 316862 207978
rect 316434 190294 316490 190350
rect 316558 190294 316614 190350
rect 316682 190294 316738 190350
rect 316806 190294 316862 190350
rect 316434 190170 316490 190226
rect 316558 190170 316614 190226
rect 316682 190170 316738 190226
rect 316806 190170 316862 190226
rect 316434 190046 316490 190102
rect 316558 190046 316614 190102
rect 316682 190046 316738 190102
rect 316806 190046 316862 190102
rect 316434 189922 316490 189978
rect 316558 189922 316614 189978
rect 316682 189922 316738 189978
rect 316806 189922 316862 189978
rect 316434 172294 316490 172350
rect 316558 172294 316614 172350
rect 316682 172294 316738 172350
rect 316806 172294 316862 172350
rect 316434 172170 316490 172226
rect 316558 172170 316614 172226
rect 316682 172170 316738 172226
rect 316806 172170 316862 172226
rect 316434 172046 316490 172102
rect 316558 172046 316614 172102
rect 316682 172046 316738 172102
rect 316806 172046 316862 172102
rect 316434 171922 316490 171978
rect 316558 171922 316614 171978
rect 316682 171922 316738 171978
rect 316806 171922 316862 171978
rect 316434 154294 316490 154350
rect 316558 154294 316614 154350
rect 316682 154294 316738 154350
rect 316806 154294 316862 154350
rect 316434 154170 316490 154226
rect 316558 154170 316614 154226
rect 316682 154170 316738 154226
rect 316806 154170 316862 154226
rect 316434 154046 316490 154102
rect 316558 154046 316614 154102
rect 316682 154046 316738 154102
rect 316806 154046 316862 154102
rect 316434 153922 316490 153978
rect 316558 153922 316614 153978
rect 316682 153922 316738 153978
rect 316806 153922 316862 153978
rect 316434 136294 316490 136350
rect 316558 136294 316614 136350
rect 316682 136294 316738 136350
rect 316806 136294 316862 136350
rect 316434 136170 316490 136226
rect 316558 136170 316614 136226
rect 316682 136170 316738 136226
rect 316806 136170 316862 136226
rect 316434 136046 316490 136102
rect 316558 136046 316614 136102
rect 316682 136046 316738 136102
rect 316806 136046 316862 136102
rect 316434 135922 316490 135978
rect 316558 135922 316614 135978
rect 316682 135922 316738 135978
rect 316806 135922 316862 135978
rect 316434 118294 316490 118350
rect 316558 118294 316614 118350
rect 316682 118294 316738 118350
rect 316806 118294 316862 118350
rect 316434 118170 316490 118226
rect 316558 118170 316614 118226
rect 316682 118170 316738 118226
rect 316806 118170 316862 118226
rect 316434 118046 316490 118102
rect 316558 118046 316614 118102
rect 316682 118046 316738 118102
rect 316806 118046 316862 118102
rect 316434 117922 316490 117978
rect 316558 117922 316614 117978
rect 316682 117922 316738 117978
rect 316806 117922 316862 117978
rect 316434 100294 316490 100350
rect 316558 100294 316614 100350
rect 316682 100294 316738 100350
rect 316806 100294 316862 100350
rect 316434 100170 316490 100226
rect 316558 100170 316614 100226
rect 316682 100170 316738 100226
rect 316806 100170 316862 100226
rect 316434 100046 316490 100102
rect 316558 100046 316614 100102
rect 316682 100046 316738 100102
rect 316806 100046 316862 100102
rect 316434 99922 316490 99978
rect 316558 99922 316614 99978
rect 316682 99922 316738 99978
rect 316806 99922 316862 99978
rect 316160 82091 316216 82147
rect 316264 82091 316320 82147
rect 316368 82091 316424 82147
rect 316160 81987 316216 82043
rect 316264 81987 316320 82043
rect 316368 81987 316424 82043
rect 316160 81883 316216 81939
rect 316264 81883 316320 81939
rect 316368 81883 316424 81939
rect 320360 76294 320416 76350
rect 320484 76294 320540 76350
rect 320360 76170 320416 76226
rect 320484 76170 320540 76226
rect 320360 76046 320416 76102
rect 320484 76046 320540 76102
rect 320360 75922 320416 75978
rect 320484 75922 320540 75978
rect 316202 64294 316258 64350
rect 316326 64294 316382 64350
rect 316202 64170 316258 64226
rect 316326 64170 316382 64226
rect 316202 64046 316258 64102
rect 316326 64046 316382 64102
rect 316202 63922 316258 63978
rect 316326 63922 316382 63978
rect 320360 58294 320416 58350
rect 320484 58294 320540 58350
rect 320360 58170 320416 58226
rect 320484 58170 320540 58226
rect 320360 58046 320416 58102
rect 320484 58046 320540 58102
rect 320360 57922 320416 57978
rect 320484 57922 320540 57978
rect 312714 40294 312770 40350
rect 312838 40294 312894 40350
rect 312962 40294 313018 40350
rect 313086 40294 313142 40350
rect 312714 40170 312770 40226
rect 312838 40170 312894 40226
rect 312962 40170 313018 40226
rect 313086 40170 313142 40226
rect 312714 40046 312770 40102
rect 312838 40046 312894 40102
rect 312962 40046 313018 40102
rect 313086 40046 313142 40102
rect 312714 39922 312770 39978
rect 312838 39922 312894 39978
rect 312962 39922 313018 39978
rect 313086 39922 313142 39978
rect 312714 22294 312770 22350
rect 312838 22294 312894 22350
rect 312962 22294 313018 22350
rect 313086 22294 313142 22350
rect 312714 22170 312770 22226
rect 312838 22170 312894 22226
rect 312962 22170 313018 22226
rect 313086 22170 313142 22226
rect 312714 22046 312770 22102
rect 312838 22046 312894 22102
rect 312962 22046 313018 22102
rect 313086 22046 313142 22102
rect 312714 21922 312770 21978
rect 312838 21922 312894 21978
rect 312962 21922 313018 21978
rect 313086 21922 313142 21978
rect 285714 -1176 285770 -1120
rect 285838 -1176 285894 -1120
rect 285962 -1176 286018 -1120
rect 286086 -1176 286142 -1120
rect 285714 -1300 285770 -1244
rect 285838 -1300 285894 -1244
rect 285962 -1300 286018 -1244
rect 286086 -1300 286142 -1244
rect 285714 -1424 285770 -1368
rect 285838 -1424 285894 -1368
rect 285962 -1424 286018 -1368
rect 286086 -1424 286142 -1368
rect 285714 -1548 285770 -1492
rect 285838 -1548 285894 -1492
rect 285962 -1548 286018 -1492
rect 286086 -1548 286142 -1492
rect 312714 4294 312770 4350
rect 312838 4294 312894 4350
rect 312962 4294 313018 4350
rect 313086 4294 313142 4350
rect 312714 4170 312770 4226
rect 312838 4170 312894 4226
rect 312962 4170 313018 4226
rect 313086 4170 313142 4226
rect 312714 4046 312770 4102
rect 312838 4046 312894 4102
rect 312962 4046 313018 4102
rect 313086 4046 313142 4102
rect 312714 3922 312770 3978
rect 312838 3922 312894 3978
rect 312962 3922 313018 3978
rect 313086 3922 313142 3978
rect 312714 -216 312770 -160
rect 312838 -216 312894 -160
rect 312962 -216 313018 -160
rect 313086 -216 313142 -160
rect 312714 -340 312770 -284
rect 312838 -340 312894 -284
rect 312962 -340 313018 -284
rect 313086 -340 313142 -284
rect 312714 -464 312770 -408
rect 312838 -464 312894 -408
rect 312962 -464 313018 -408
rect 313086 -464 313142 -408
rect 312714 -588 312770 -532
rect 312838 -588 312894 -532
rect 312962 -588 313018 -532
rect 313086 -588 313142 -532
rect 343434 202294 343490 202350
rect 343558 202294 343614 202350
rect 343682 202294 343738 202350
rect 343806 202294 343862 202350
rect 343434 202170 343490 202226
rect 343558 202170 343614 202226
rect 343682 202170 343738 202226
rect 343806 202170 343862 202226
rect 343434 202046 343490 202102
rect 343558 202046 343614 202102
rect 343682 202046 343738 202102
rect 343806 202046 343862 202102
rect 343434 201922 343490 201978
rect 343558 201922 343614 201978
rect 343682 201922 343738 201978
rect 343806 201922 343862 201978
rect 343434 184294 343490 184350
rect 343558 184294 343614 184350
rect 343682 184294 343738 184350
rect 343806 184294 343862 184350
rect 343434 184170 343490 184226
rect 343558 184170 343614 184226
rect 343682 184170 343738 184226
rect 343806 184170 343862 184226
rect 343434 184046 343490 184102
rect 343558 184046 343614 184102
rect 343682 184046 343738 184102
rect 343806 184046 343862 184102
rect 343434 183922 343490 183978
rect 343558 183922 343614 183978
rect 343682 183922 343738 183978
rect 343806 183922 343862 183978
rect 343434 166294 343490 166350
rect 343558 166294 343614 166350
rect 343682 166294 343738 166350
rect 343806 166294 343862 166350
rect 343434 166170 343490 166226
rect 343558 166170 343614 166226
rect 343682 166170 343738 166226
rect 343806 166170 343862 166226
rect 343434 166046 343490 166102
rect 343558 166046 343614 166102
rect 343682 166046 343738 166102
rect 343806 166046 343862 166102
rect 343434 165922 343490 165978
rect 343558 165922 343614 165978
rect 343682 165922 343738 165978
rect 343806 165922 343862 165978
rect 343434 148294 343490 148350
rect 343558 148294 343614 148350
rect 343682 148294 343738 148350
rect 343806 148294 343862 148350
rect 343434 148170 343490 148226
rect 343558 148170 343614 148226
rect 343682 148170 343738 148226
rect 343806 148170 343862 148226
rect 343434 148046 343490 148102
rect 343558 148046 343614 148102
rect 343682 148046 343738 148102
rect 343806 148046 343862 148102
rect 343434 147922 343490 147978
rect 343558 147922 343614 147978
rect 343682 147922 343738 147978
rect 343806 147922 343862 147978
rect 343434 130294 343490 130350
rect 343558 130294 343614 130350
rect 343682 130294 343738 130350
rect 343806 130294 343862 130350
rect 343434 130170 343490 130226
rect 343558 130170 343614 130226
rect 343682 130170 343738 130226
rect 343806 130170 343862 130226
rect 343434 130046 343490 130102
rect 343558 130046 343614 130102
rect 343682 130046 343738 130102
rect 343806 130046 343862 130102
rect 343434 129922 343490 129978
rect 343558 129922 343614 129978
rect 343682 129922 343738 129978
rect 343806 129922 343862 129978
rect 343434 112294 343490 112350
rect 343558 112294 343614 112350
rect 343682 112294 343738 112350
rect 343806 112294 343862 112350
rect 343434 112170 343490 112226
rect 343558 112170 343614 112226
rect 343682 112170 343738 112226
rect 343806 112170 343862 112226
rect 343434 112046 343490 112102
rect 343558 112046 343614 112102
rect 343682 112046 343738 112102
rect 343806 112046 343862 112102
rect 343434 111922 343490 111978
rect 343558 111922 343614 111978
rect 343682 111922 343738 111978
rect 343806 111922 343862 111978
rect 343434 94294 343490 94350
rect 343558 94294 343614 94350
rect 343682 94294 343738 94350
rect 343806 94294 343862 94350
rect 343434 94170 343490 94226
rect 343558 94170 343614 94226
rect 343682 94170 343738 94226
rect 343806 94170 343862 94226
rect 343434 94046 343490 94102
rect 343558 94046 343614 94102
rect 343682 94046 343738 94102
rect 343806 94046 343862 94102
rect 343434 93922 343490 93978
rect 343558 93922 343614 93978
rect 343682 93922 343738 93978
rect 343806 93922 343862 93978
rect 324476 82091 324532 82147
rect 324580 82091 324636 82147
rect 324684 82091 324740 82147
rect 324476 81987 324532 82043
rect 324580 81987 324636 82043
rect 324684 81987 324740 82043
rect 324476 81883 324532 81939
rect 324580 81883 324636 81939
rect 324684 81883 324740 81939
rect 343434 76294 343490 76350
rect 343558 76294 343614 76350
rect 343682 76294 343738 76350
rect 343806 76294 343862 76350
rect 343434 76170 343490 76226
rect 343558 76170 343614 76226
rect 343682 76170 343738 76226
rect 343806 76170 343862 76226
rect 343434 76046 343490 76102
rect 343558 76046 343614 76102
rect 343682 76046 343738 76102
rect 343806 76046 343862 76102
rect 343434 75922 343490 75978
rect 343558 75922 343614 75978
rect 343682 75922 343738 75978
rect 343806 75922 343862 75978
rect 324518 64294 324574 64350
rect 324642 64294 324698 64350
rect 324518 64170 324574 64226
rect 324642 64170 324698 64226
rect 324518 64046 324574 64102
rect 324642 64046 324698 64102
rect 324518 63922 324574 63978
rect 324642 63922 324698 63978
rect 343434 58294 343490 58350
rect 343558 58294 343614 58350
rect 343682 58294 343738 58350
rect 343806 58294 343862 58350
rect 343434 58170 343490 58226
rect 343558 58170 343614 58226
rect 343682 58170 343738 58226
rect 343806 58170 343862 58226
rect 343434 58046 343490 58102
rect 343558 58046 343614 58102
rect 343682 58046 343738 58102
rect 343806 58046 343862 58102
rect 343434 57922 343490 57978
rect 343558 57922 343614 57978
rect 343682 57922 343738 57978
rect 343806 57922 343862 57978
rect 316434 46294 316490 46350
rect 316558 46294 316614 46350
rect 316682 46294 316738 46350
rect 316806 46294 316862 46350
rect 316434 46170 316490 46226
rect 316558 46170 316614 46226
rect 316682 46170 316738 46226
rect 316806 46170 316862 46226
rect 316434 46046 316490 46102
rect 316558 46046 316614 46102
rect 316682 46046 316738 46102
rect 316806 46046 316862 46102
rect 316434 45922 316490 45978
rect 316558 45922 316614 45978
rect 316682 45922 316738 45978
rect 316806 45922 316862 45978
rect 316434 28294 316490 28350
rect 316558 28294 316614 28350
rect 316682 28294 316738 28350
rect 316806 28294 316862 28350
rect 316434 28170 316490 28226
rect 316558 28170 316614 28226
rect 316682 28170 316738 28226
rect 316806 28170 316862 28226
rect 316434 28046 316490 28102
rect 316558 28046 316614 28102
rect 316682 28046 316738 28102
rect 316806 28046 316862 28102
rect 316434 27922 316490 27978
rect 316558 27922 316614 27978
rect 316682 27922 316738 27978
rect 316806 27922 316862 27978
rect 316434 10294 316490 10350
rect 316558 10294 316614 10350
rect 316682 10294 316738 10350
rect 316806 10294 316862 10350
rect 316434 10170 316490 10226
rect 316558 10170 316614 10226
rect 316682 10170 316738 10226
rect 316806 10170 316862 10226
rect 316434 10046 316490 10102
rect 316558 10046 316614 10102
rect 316682 10046 316738 10102
rect 316806 10046 316862 10102
rect 316434 9922 316490 9978
rect 316558 9922 316614 9978
rect 316682 9922 316738 9978
rect 316806 9922 316862 9978
rect 316434 -1176 316490 -1120
rect 316558 -1176 316614 -1120
rect 316682 -1176 316738 -1120
rect 316806 -1176 316862 -1120
rect 316434 -1300 316490 -1244
rect 316558 -1300 316614 -1244
rect 316682 -1300 316738 -1244
rect 316806 -1300 316862 -1244
rect 316434 -1424 316490 -1368
rect 316558 -1424 316614 -1368
rect 316682 -1424 316738 -1368
rect 316806 -1424 316862 -1368
rect 316434 -1548 316490 -1492
rect 316558 -1548 316614 -1492
rect 316682 -1548 316738 -1492
rect 316806 -1548 316862 -1492
rect 343434 40294 343490 40350
rect 343558 40294 343614 40350
rect 343682 40294 343738 40350
rect 343806 40294 343862 40350
rect 343434 40170 343490 40226
rect 343558 40170 343614 40226
rect 343682 40170 343738 40226
rect 343806 40170 343862 40226
rect 343434 40046 343490 40102
rect 343558 40046 343614 40102
rect 343682 40046 343738 40102
rect 343806 40046 343862 40102
rect 343434 39922 343490 39978
rect 343558 39922 343614 39978
rect 343682 39922 343738 39978
rect 343806 39922 343862 39978
rect 343434 22294 343490 22350
rect 343558 22294 343614 22350
rect 343682 22294 343738 22350
rect 343806 22294 343862 22350
rect 343434 22170 343490 22226
rect 343558 22170 343614 22226
rect 343682 22170 343738 22226
rect 343806 22170 343862 22226
rect 343434 22046 343490 22102
rect 343558 22046 343614 22102
rect 343682 22046 343738 22102
rect 343806 22046 343862 22102
rect 343434 21922 343490 21978
rect 343558 21922 343614 21978
rect 343682 21922 343738 21978
rect 343806 21922 343862 21978
rect 343434 4294 343490 4350
rect 343558 4294 343614 4350
rect 343682 4294 343738 4350
rect 343806 4294 343862 4350
rect 343434 4170 343490 4226
rect 343558 4170 343614 4226
rect 343682 4170 343738 4226
rect 343806 4170 343862 4226
rect 343434 4046 343490 4102
rect 343558 4046 343614 4102
rect 343682 4046 343738 4102
rect 343806 4046 343862 4102
rect 343434 3922 343490 3978
rect 343558 3922 343614 3978
rect 343682 3922 343738 3978
rect 343806 3922 343862 3978
rect 343434 -216 343490 -160
rect 343558 -216 343614 -160
rect 343682 -216 343738 -160
rect 343806 -216 343862 -160
rect 343434 -340 343490 -284
rect 343558 -340 343614 -284
rect 343682 -340 343738 -284
rect 343806 -340 343862 -284
rect 343434 -464 343490 -408
rect 343558 -464 343614 -408
rect 343682 -464 343738 -408
rect 343806 -464 343862 -408
rect 343434 -588 343490 -532
rect 343558 -588 343614 -532
rect 343682 -588 343738 -532
rect 343806 -588 343862 -532
rect 347154 244294 347210 244350
rect 347278 244294 347334 244350
rect 347402 244294 347458 244350
rect 347526 244294 347582 244350
rect 347154 244170 347210 244226
rect 347278 244170 347334 244226
rect 347402 244170 347458 244226
rect 347526 244170 347582 244226
rect 347154 244046 347210 244102
rect 347278 244046 347334 244102
rect 347402 244046 347458 244102
rect 347526 244046 347582 244102
rect 347154 243922 347210 243978
rect 347278 243922 347334 243978
rect 347402 243922 347458 243978
rect 347526 243922 347582 243978
rect 347154 226294 347210 226350
rect 347278 226294 347334 226350
rect 347402 226294 347458 226350
rect 347526 226294 347582 226350
rect 347154 226170 347210 226226
rect 347278 226170 347334 226226
rect 347402 226170 347458 226226
rect 347526 226170 347582 226226
rect 347154 226046 347210 226102
rect 347278 226046 347334 226102
rect 347402 226046 347458 226102
rect 347526 226046 347582 226102
rect 347154 225922 347210 225978
rect 347278 225922 347334 225978
rect 347402 225922 347458 225978
rect 347526 225922 347582 225978
rect 347154 208294 347210 208350
rect 347278 208294 347334 208350
rect 347402 208294 347458 208350
rect 347526 208294 347582 208350
rect 347154 208170 347210 208226
rect 347278 208170 347334 208226
rect 347402 208170 347458 208226
rect 347526 208170 347582 208226
rect 347154 208046 347210 208102
rect 347278 208046 347334 208102
rect 347402 208046 347458 208102
rect 347526 208046 347582 208102
rect 347154 207922 347210 207978
rect 347278 207922 347334 207978
rect 347402 207922 347458 207978
rect 347526 207922 347582 207978
rect 347154 190294 347210 190350
rect 347278 190294 347334 190350
rect 347402 190294 347458 190350
rect 347526 190294 347582 190350
rect 347154 190170 347210 190226
rect 347278 190170 347334 190226
rect 347402 190170 347458 190226
rect 347526 190170 347582 190226
rect 347154 190046 347210 190102
rect 347278 190046 347334 190102
rect 347402 190046 347458 190102
rect 347526 190046 347582 190102
rect 347154 189922 347210 189978
rect 347278 189922 347334 189978
rect 347402 189922 347458 189978
rect 347526 189922 347582 189978
rect 347154 172294 347210 172350
rect 347278 172294 347334 172350
rect 347402 172294 347458 172350
rect 347526 172294 347582 172350
rect 347154 172170 347210 172226
rect 347278 172170 347334 172226
rect 347402 172170 347458 172226
rect 347526 172170 347582 172226
rect 347154 172046 347210 172102
rect 347278 172046 347334 172102
rect 347402 172046 347458 172102
rect 347526 172046 347582 172102
rect 347154 171922 347210 171978
rect 347278 171922 347334 171978
rect 347402 171922 347458 171978
rect 347526 171922 347582 171978
rect 347154 154294 347210 154350
rect 347278 154294 347334 154350
rect 347402 154294 347458 154350
rect 347526 154294 347582 154350
rect 347154 154170 347210 154226
rect 347278 154170 347334 154226
rect 347402 154170 347458 154226
rect 347526 154170 347582 154226
rect 347154 154046 347210 154102
rect 347278 154046 347334 154102
rect 347402 154046 347458 154102
rect 347526 154046 347582 154102
rect 347154 153922 347210 153978
rect 347278 153922 347334 153978
rect 347402 153922 347458 153978
rect 347526 153922 347582 153978
rect 347154 136294 347210 136350
rect 347278 136294 347334 136350
rect 347402 136294 347458 136350
rect 347526 136294 347582 136350
rect 347154 136170 347210 136226
rect 347278 136170 347334 136226
rect 347402 136170 347458 136226
rect 347526 136170 347582 136226
rect 347154 136046 347210 136102
rect 347278 136046 347334 136102
rect 347402 136046 347458 136102
rect 347526 136046 347582 136102
rect 347154 135922 347210 135978
rect 347278 135922 347334 135978
rect 347402 135922 347458 135978
rect 347526 135922 347582 135978
rect 347154 118294 347210 118350
rect 347278 118294 347334 118350
rect 347402 118294 347458 118350
rect 347526 118294 347582 118350
rect 347154 118170 347210 118226
rect 347278 118170 347334 118226
rect 347402 118170 347458 118226
rect 347526 118170 347582 118226
rect 347154 118046 347210 118102
rect 347278 118046 347334 118102
rect 347402 118046 347458 118102
rect 347526 118046 347582 118102
rect 347154 117922 347210 117978
rect 347278 117922 347334 117978
rect 347402 117922 347458 117978
rect 347526 117922 347582 117978
rect 347154 100294 347210 100350
rect 347278 100294 347334 100350
rect 347402 100294 347458 100350
rect 347526 100294 347582 100350
rect 347154 100170 347210 100226
rect 347278 100170 347334 100226
rect 347402 100170 347458 100226
rect 347526 100170 347582 100226
rect 347154 100046 347210 100102
rect 347278 100046 347334 100102
rect 347402 100046 347458 100102
rect 347526 100046 347582 100102
rect 347154 99922 347210 99978
rect 347278 99922 347334 99978
rect 347402 99922 347458 99978
rect 347526 99922 347582 99978
rect 347154 82294 347210 82350
rect 347278 82294 347334 82350
rect 347402 82294 347458 82350
rect 347526 82294 347582 82350
rect 347154 82170 347210 82226
rect 347278 82170 347334 82226
rect 347402 82170 347458 82226
rect 347526 82170 347582 82226
rect 347154 82046 347210 82102
rect 347278 82046 347334 82102
rect 347402 82046 347458 82102
rect 347526 82046 347582 82102
rect 347154 81922 347210 81978
rect 347278 81922 347334 81978
rect 347402 81922 347458 81978
rect 347526 81922 347582 81978
rect 347154 64294 347210 64350
rect 347278 64294 347334 64350
rect 347402 64294 347458 64350
rect 347526 64294 347582 64350
rect 347154 64170 347210 64226
rect 347278 64170 347334 64226
rect 347402 64170 347458 64226
rect 347526 64170 347582 64226
rect 347154 64046 347210 64102
rect 347278 64046 347334 64102
rect 347402 64046 347458 64102
rect 347526 64046 347582 64102
rect 347154 63922 347210 63978
rect 347278 63922 347334 63978
rect 347402 63922 347458 63978
rect 347526 63922 347582 63978
rect 347154 46294 347210 46350
rect 347278 46294 347334 46350
rect 347402 46294 347458 46350
rect 347526 46294 347582 46350
rect 347154 46170 347210 46226
rect 347278 46170 347334 46226
rect 347402 46170 347458 46226
rect 347526 46170 347582 46226
rect 347154 46046 347210 46102
rect 347278 46046 347334 46102
rect 347402 46046 347458 46102
rect 347526 46046 347582 46102
rect 347154 45922 347210 45978
rect 347278 45922 347334 45978
rect 347402 45922 347458 45978
rect 347526 45922 347582 45978
rect 347154 28294 347210 28350
rect 347278 28294 347334 28350
rect 347402 28294 347458 28350
rect 347526 28294 347582 28350
rect 347154 28170 347210 28226
rect 347278 28170 347334 28226
rect 347402 28170 347458 28226
rect 347526 28170 347582 28226
rect 347154 28046 347210 28102
rect 347278 28046 347334 28102
rect 347402 28046 347458 28102
rect 347526 28046 347582 28102
rect 347154 27922 347210 27978
rect 347278 27922 347334 27978
rect 347402 27922 347458 27978
rect 347526 27922 347582 27978
rect 347154 10294 347210 10350
rect 347278 10294 347334 10350
rect 347402 10294 347458 10350
rect 347526 10294 347582 10350
rect 347154 10170 347210 10226
rect 347278 10170 347334 10226
rect 347402 10170 347458 10226
rect 347526 10170 347582 10226
rect 347154 10046 347210 10102
rect 347278 10046 347334 10102
rect 347402 10046 347458 10102
rect 347526 10046 347582 10102
rect 347154 9922 347210 9978
rect 347278 9922 347334 9978
rect 347402 9922 347458 9978
rect 347526 9922 347582 9978
rect 358764 253142 358820 253198
rect 358988 252962 359044 253018
rect 359212 252782 359268 252838
rect 373100 385622 373156 385678
rect 373772 288242 373828 288298
rect 375228 288242 375284 288298
rect 373884 286082 373940 286138
rect 375228 286132 375284 286138
rect 375228 286082 375284 286132
rect 375228 257822 375284 257878
rect 373884 253142 373940 253198
rect 374154 256294 374210 256350
rect 374278 256294 374334 256350
rect 374402 256294 374458 256350
rect 374526 256294 374582 256350
rect 374154 256170 374210 256226
rect 374278 256170 374334 256226
rect 374402 256170 374458 256226
rect 374526 256170 374582 256226
rect 374154 256046 374210 256102
rect 374278 256046 374334 256102
rect 374402 256046 374458 256102
rect 374526 256046 374582 256102
rect 374154 255922 374210 255978
rect 374278 255922 374334 255978
rect 374402 255922 374458 255978
rect 374526 255922 374582 255978
rect 374154 238294 374210 238350
rect 374278 238294 374334 238350
rect 374402 238294 374458 238350
rect 374526 238294 374582 238350
rect 374154 238170 374210 238226
rect 374278 238170 374334 238226
rect 374402 238170 374458 238226
rect 374526 238170 374582 238226
rect 374154 238046 374210 238102
rect 374278 238046 374334 238102
rect 374402 238046 374458 238102
rect 374526 238046 374582 238102
rect 374154 237922 374210 237978
rect 374278 237922 374334 237978
rect 374402 237922 374458 237978
rect 374526 237922 374582 237978
rect 374154 220294 374210 220350
rect 374278 220294 374334 220350
rect 374402 220294 374458 220350
rect 374526 220294 374582 220350
rect 374154 220170 374210 220226
rect 374278 220170 374334 220226
rect 374402 220170 374458 220226
rect 374526 220170 374582 220226
rect 374154 220046 374210 220102
rect 374278 220046 374334 220102
rect 374402 220046 374458 220102
rect 374526 220046 374582 220102
rect 374154 219922 374210 219978
rect 374278 219922 374334 219978
rect 374402 219922 374458 219978
rect 374526 219922 374582 219978
rect 374154 202294 374210 202350
rect 374278 202294 374334 202350
rect 374402 202294 374458 202350
rect 374526 202294 374582 202350
rect 374154 202170 374210 202226
rect 374278 202170 374334 202226
rect 374402 202170 374458 202226
rect 374526 202170 374582 202226
rect 374154 202046 374210 202102
rect 374278 202046 374334 202102
rect 374402 202046 374458 202102
rect 374526 202046 374582 202102
rect 374154 201922 374210 201978
rect 374278 201922 374334 201978
rect 374402 201922 374458 201978
rect 374526 201922 374582 201978
rect 374154 184294 374210 184350
rect 374278 184294 374334 184350
rect 374402 184294 374458 184350
rect 374526 184294 374582 184350
rect 374154 184170 374210 184226
rect 374278 184170 374334 184226
rect 374402 184170 374458 184226
rect 374526 184170 374582 184226
rect 374154 184046 374210 184102
rect 374278 184046 374334 184102
rect 374402 184046 374458 184102
rect 374526 184046 374582 184102
rect 374154 183922 374210 183978
rect 374278 183922 374334 183978
rect 374402 183922 374458 183978
rect 374526 183922 374582 183978
rect 374154 166294 374210 166350
rect 374278 166294 374334 166350
rect 374402 166294 374458 166350
rect 374526 166294 374582 166350
rect 374154 166170 374210 166226
rect 374278 166170 374334 166226
rect 374402 166170 374458 166226
rect 374526 166170 374582 166226
rect 374154 166046 374210 166102
rect 374278 166046 374334 166102
rect 374402 166046 374458 166102
rect 374526 166046 374582 166102
rect 374154 165922 374210 165978
rect 374278 165922 374334 165978
rect 374402 165922 374458 165978
rect 374526 165922 374582 165978
rect 372428 153602 372484 153658
rect 377874 406294 377930 406350
rect 377998 406294 378054 406350
rect 378122 406294 378178 406350
rect 378246 406294 378302 406350
rect 377874 406170 377930 406226
rect 377998 406170 378054 406226
rect 378122 406170 378178 406226
rect 378246 406170 378302 406226
rect 377874 406046 377930 406102
rect 377998 406046 378054 406102
rect 378122 406046 378178 406102
rect 378246 406046 378302 406102
rect 377874 405922 377930 405978
rect 377998 405922 378054 405978
rect 378122 405922 378178 405978
rect 378246 405922 378302 405978
rect 377874 388294 377930 388350
rect 377998 388294 378054 388350
rect 378122 388294 378178 388350
rect 378246 388294 378302 388350
rect 377874 388170 377930 388226
rect 377998 388170 378054 388226
rect 378122 388170 378178 388226
rect 378246 388170 378302 388226
rect 377874 388046 377930 388102
rect 377998 388046 378054 388102
rect 378122 388046 378178 388102
rect 378246 388046 378302 388102
rect 377874 387922 377930 387978
rect 377998 387922 378054 387978
rect 378122 387922 378178 387978
rect 378246 387922 378302 387978
rect 377874 370294 377930 370350
rect 377998 370294 378054 370350
rect 378122 370294 378178 370350
rect 378246 370294 378302 370350
rect 377874 370170 377930 370226
rect 377998 370170 378054 370226
rect 378122 370170 378178 370226
rect 378246 370170 378302 370226
rect 377874 370046 377930 370102
rect 377998 370046 378054 370102
rect 378122 370046 378178 370102
rect 378246 370046 378302 370102
rect 377874 369922 377930 369978
rect 377998 369922 378054 369978
rect 378122 369922 378178 369978
rect 378246 369922 378302 369978
rect 377874 352294 377930 352350
rect 377998 352294 378054 352350
rect 378122 352294 378178 352350
rect 378246 352294 378302 352350
rect 377874 352170 377930 352226
rect 377998 352170 378054 352226
rect 378122 352170 378178 352226
rect 378246 352170 378302 352226
rect 377874 352046 377930 352102
rect 377998 352046 378054 352102
rect 378122 352046 378178 352102
rect 378246 352046 378302 352102
rect 377874 351922 377930 351978
rect 377998 351922 378054 351978
rect 378122 351922 378178 351978
rect 378246 351922 378302 351978
rect 377874 334294 377930 334350
rect 377998 334294 378054 334350
rect 378122 334294 378178 334350
rect 378246 334294 378302 334350
rect 377874 334170 377930 334226
rect 377998 334170 378054 334226
rect 378122 334170 378178 334226
rect 378246 334170 378302 334226
rect 377874 334046 377930 334102
rect 377998 334046 378054 334102
rect 378122 334046 378178 334102
rect 378246 334046 378302 334102
rect 377874 333922 377930 333978
rect 377998 333922 378054 333978
rect 378122 333922 378178 333978
rect 378246 333922 378302 333978
rect 404874 400294 404930 400350
rect 404998 400294 405054 400350
rect 405122 400294 405178 400350
rect 405246 400294 405302 400350
rect 404874 400170 404930 400226
rect 404998 400170 405054 400226
rect 405122 400170 405178 400226
rect 405246 400170 405302 400226
rect 404874 400046 404930 400102
rect 404998 400046 405054 400102
rect 405122 400046 405178 400102
rect 405246 400046 405302 400102
rect 404874 399922 404930 399978
rect 404998 399922 405054 399978
rect 405122 399922 405178 399978
rect 405246 399922 405302 399978
rect 377874 316294 377930 316350
rect 377998 316294 378054 316350
rect 378122 316294 378178 316350
rect 378246 316294 378302 316350
rect 377874 316170 377930 316226
rect 377998 316170 378054 316226
rect 378122 316170 378178 316226
rect 378246 316170 378302 316226
rect 377874 316046 377930 316102
rect 377998 316046 378054 316102
rect 378122 316046 378178 316102
rect 378246 316046 378302 316102
rect 377874 315922 377930 315978
rect 377998 315922 378054 315978
rect 378122 315922 378178 315978
rect 378246 315922 378302 315978
rect 375676 252962 375732 253018
rect 383964 388682 384020 388738
rect 377874 298294 377930 298350
rect 377998 298294 378054 298350
rect 378122 298294 378178 298350
rect 378246 298294 378302 298350
rect 377874 298170 377930 298226
rect 377998 298170 378054 298226
rect 378122 298170 378178 298226
rect 378246 298170 378302 298226
rect 377874 298046 377930 298102
rect 377998 298046 378054 298102
rect 378122 298046 378178 298102
rect 378246 298046 378302 298102
rect 377874 297922 377930 297978
rect 377998 297922 378054 297978
rect 378122 297922 378178 297978
rect 378246 297922 378302 297978
rect 376460 252782 376516 252838
rect 377874 280294 377930 280350
rect 377998 280294 378054 280350
rect 378122 280294 378178 280350
rect 378246 280294 378302 280350
rect 377874 280170 377930 280226
rect 377998 280170 378054 280226
rect 378122 280170 378178 280226
rect 378246 280170 378302 280226
rect 377874 280046 377930 280102
rect 377998 280046 378054 280102
rect 378122 280046 378178 280102
rect 378246 280046 378302 280102
rect 377874 279922 377930 279978
rect 377998 279922 378054 279978
rect 378122 279922 378178 279978
rect 378246 279922 378302 279978
rect 377874 262294 377930 262350
rect 377998 262294 378054 262350
rect 378122 262294 378178 262350
rect 378246 262294 378302 262350
rect 377874 262170 377930 262226
rect 377998 262170 378054 262226
rect 378122 262170 378178 262226
rect 378246 262170 378302 262226
rect 377874 262046 377930 262102
rect 377998 262046 378054 262102
rect 378122 262046 378178 262102
rect 378246 262046 378302 262102
rect 377874 261922 377930 261978
rect 377998 261922 378054 261978
rect 378122 261922 378178 261978
rect 378246 261922 378302 261978
rect 377874 244294 377930 244350
rect 377998 244294 378054 244350
rect 378122 244294 378178 244350
rect 378246 244294 378302 244350
rect 377874 244170 377930 244226
rect 377998 244170 378054 244226
rect 378122 244170 378178 244226
rect 378246 244170 378302 244226
rect 377874 244046 377930 244102
rect 377998 244046 378054 244102
rect 378122 244046 378178 244102
rect 378246 244046 378302 244102
rect 377874 243922 377930 243978
rect 377998 243922 378054 243978
rect 378122 243922 378178 243978
rect 378246 243922 378302 243978
rect 377874 226294 377930 226350
rect 377998 226294 378054 226350
rect 378122 226294 378178 226350
rect 378246 226294 378302 226350
rect 377874 226170 377930 226226
rect 377998 226170 378054 226226
rect 378122 226170 378178 226226
rect 378246 226170 378302 226226
rect 377874 226046 377930 226102
rect 377998 226046 378054 226102
rect 378122 226046 378178 226102
rect 378246 226046 378302 226102
rect 377874 225922 377930 225978
rect 377998 225922 378054 225978
rect 378122 225922 378178 225978
rect 378246 225922 378302 225978
rect 377874 208294 377930 208350
rect 377998 208294 378054 208350
rect 378122 208294 378178 208350
rect 378246 208294 378302 208350
rect 377874 208170 377930 208226
rect 377998 208170 378054 208226
rect 378122 208170 378178 208226
rect 378246 208170 378302 208226
rect 377874 208046 377930 208102
rect 377998 208046 378054 208102
rect 378122 208046 378178 208102
rect 378246 208046 378302 208102
rect 377874 207922 377930 207978
rect 377998 207922 378054 207978
rect 378122 207922 378178 207978
rect 378246 207922 378302 207978
rect 377874 190294 377930 190350
rect 377998 190294 378054 190350
rect 378122 190294 378178 190350
rect 378246 190294 378302 190350
rect 377874 190170 377930 190226
rect 377998 190170 378054 190226
rect 378122 190170 378178 190226
rect 378246 190170 378302 190226
rect 377874 190046 377930 190102
rect 377998 190046 378054 190102
rect 378122 190046 378178 190102
rect 378246 190046 378302 190102
rect 377874 189922 377930 189978
rect 377998 189922 378054 189978
rect 378122 189922 378178 189978
rect 378246 189922 378302 189978
rect 377874 172294 377930 172350
rect 377998 172294 378054 172350
rect 378122 172294 378178 172350
rect 378246 172294 378302 172350
rect 377874 172170 377930 172226
rect 377998 172170 378054 172226
rect 378122 172170 378178 172226
rect 378246 172170 378302 172226
rect 377874 172046 377930 172102
rect 377998 172046 378054 172102
rect 378122 172046 378178 172102
rect 378246 172046 378302 172102
rect 377874 171922 377930 171978
rect 377998 171922 378054 171978
rect 378122 171922 378178 171978
rect 378246 171922 378302 171978
rect 377874 154294 377930 154350
rect 377998 154294 378054 154350
rect 378122 154294 378178 154350
rect 378246 154294 378302 154350
rect 377874 154170 377930 154226
rect 377998 154170 378054 154226
rect 378122 154170 378178 154226
rect 378246 154170 378302 154226
rect 377874 154046 377930 154102
rect 377998 154046 378054 154102
rect 378122 154046 378178 154102
rect 378246 154046 378302 154102
rect 377874 153922 377930 153978
rect 377998 153922 378054 153978
rect 378122 153922 378178 153978
rect 378246 153922 378302 153978
rect 374154 148294 374210 148350
rect 374278 148294 374334 148350
rect 374402 148294 374458 148350
rect 374526 148294 374582 148350
rect 374154 148170 374210 148226
rect 374278 148170 374334 148226
rect 374402 148170 374458 148226
rect 374526 148170 374582 148226
rect 374154 148046 374210 148102
rect 374278 148046 374334 148102
rect 374402 148046 374458 148102
rect 374526 148046 374582 148102
rect 374154 147922 374210 147978
rect 374278 147922 374334 147978
rect 374402 147922 374458 147978
rect 374526 147922 374582 147978
rect 374154 130294 374210 130350
rect 374278 130294 374334 130350
rect 374402 130294 374458 130350
rect 374526 130294 374582 130350
rect 374154 130170 374210 130226
rect 374278 130170 374334 130226
rect 374402 130170 374458 130226
rect 374526 130170 374582 130226
rect 374154 130046 374210 130102
rect 374278 130046 374334 130102
rect 374402 130046 374458 130102
rect 374526 130046 374582 130102
rect 374154 129922 374210 129978
rect 374278 129922 374334 129978
rect 374402 129922 374458 129978
rect 374526 129922 374582 129978
rect 377874 136294 377930 136350
rect 377998 136294 378054 136350
rect 378122 136294 378178 136350
rect 378246 136294 378302 136350
rect 377874 136170 377930 136226
rect 377998 136170 378054 136226
rect 378122 136170 378178 136226
rect 378246 136170 378302 136226
rect 377874 136046 377930 136102
rect 377998 136046 378054 136102
rect 378122 136046 378178 136102
rect 378246 136046 378302 136102
rect 377874 135922 377930 135978
rect 377998 135922 378054 135978
rect 378122 135922 378178 135978
rect 378246 135922 378302 135978
rect 404874 382294 404930 382350
rect 404998 382294 405054 382350
rect 405122 382294 405178 382350
rect 405246 382294 405302 382350
rect 404874 382170 404930 382226
rect 404998 382170 405054 382226
rect 405122 382170 405178 382226
rect 405246 382170 405302 382226
rect 404874 382046 404930 382102
rect 404998 382046 405054 382102
rect 405122 382046 405178 382102
rect 405246 382046 405302 382102
rect 404874 381922 404930 381978
rect 404998 381922 405054 381978
rect 405122 381922 405178 381978
rect 405246 381922 405302 381978
rect 404874 364294 404930 364350
rect 404998 364294 405054 364350
rect 405122 364294 405178 364350
rect 405246 364294 405302 364350
rect 404874 364170 404930 364226
rect 404998 364170 405054 364226
rect 405122 364170 405178 364226
rect 405246 364170 405302 364226
rect 404874 364046 404930 364102
rect 404998 364046 405054 364102
rect 405122 364046 405178 364102
rect 405246 364046 405302 364102
rect 404874 363922 404930 363978
rect 404998 363922 405054 363978
rect 405122 363922 405178 363978
rect 405246 363922 405302 363978
rect 404874 346294 404930 346350
rect 404998 346294 405054 346350
rect 405122 346294 405178 346350
rect 405246 346294 405302 346350
rect 404874 346170 404930 346226
rect 404998 346170 405054 346226
rect 405122 346170 405178 346226
rect 405246 346170 405302 346226
rect 404874 346046 404930 346102
rect 404998 346046 405054 346102
rect 405122 346046 405178 346102
rect 405246 346046 405302 346102
rect 404874 345922 404930 345978
rect 404998 345922 405054 345978
rect 405122 345922 405178 345978
rect 405246 345922 405302 345978
rect 404874 328294 404930 328350
rect 404998 328294 405054 328350
rect 405122 328294 405178 328350
rect 405246 328294 405302 328350
rect 404874 328170 404930 328226
rect 404998 328170 405054 328226
rect 405122 328170 405178 328226
rect 405246 328170 405302 328226
rect 404874 328046 404930 328102
rect 404998 328046 405054 328102
rect 405122 328046 405178 328102
rect 405246 328046 405302 328102
rect 404874 327922 404930 327978
rect 404998 327922 405054 327978
rect 405122 327922 405178 327978
rect 405246 327922 405302 327978
rect 404874 310294 404930 310350
rect 404998 310294 405054 310350
rect 405122 310294 405178 310350
rect 405246 310294 405302 310350
rect 404874 310170 404930 310226
rect 404998 310170 405054 310226
rect 405122 310170 405178 310226
rect 405246 310170 405302 310226
rect 404874 310046 404930 310102
rect 404998 310046 405054 310102
rect 405122 310046 405178 310102
rect 405246 310046 405302 310102
rect 404874 309922 404930 309978
rect 404998 309922 405054 309978
rect 405122 309922 405178 309978
rect 405246 309922 405302 309978
rect 404874 292294 404930 292350
rect 404998 292294 405054 292350
rect 405122 292294 405178 292350
rect 405246 292294 405302 292350
rect 404874 292170 404930 292226
rect 404998 292170 405054 292226
rect 405122 292170 405178 292226
rect 405246 292170 405302 292226
rect 404874 292046 404930 292102
rect 404998 292046 405054 292102
rect 405122 292046 405178 292102
rect 405246 292046 405302 292102
rect 404874 291922 404930 291978
rect 404998 291922 405054 291978
rect 405122 291922 405178 291978
rect 405246 291922 405302 291978
rect 404874 274294 404930 274350
rect 404998 274294 405054 274350
rect 405122 274294 405178 274350
rect 405246 274294 405302 274350
rect 404874 274170 404930 274226
rect 404998 274170 405054 274226
rect 405122 274170 405178 274226
rect 405246 274170 405302 274226
rect 404874 274046 404930 274102
rect 404998 274046 405054 274102
rect 405122 274046 405178 274102
rect 405246 274046 405302 274102
rect 404874 273922 404930 273978
rect 404998 273922 405054 273978
rect 405122 273922 405178 273978
rect 405246 273922 405302 273978
rect 404874 256294 404930 256350
rect 404998 256294 405054 256350
rect 405122 256294 405178 256350
rect 405246 256294 405302 256350
rect 404874 256170 404930 256226
rect 404998 256170 405054 256226
rect 405122 256170 405178 256226
rect 405246 256170 405302 256226
rect 404874 256046 404930 256102
rect 404998 256046 405054 256102
rect 405122 256046 405178 256102
rect 405246 256046 405302 256102
rect 404874 255922 404930 255978
rect 404998 255922 405054 255978
rect 405122 255922 405178 255978
rect 405246 255922 405302 255978
rect 404874 238294 404930 238350
rect 404998 238294 405054 238350
rect 405122 238294 405178 238350
rect 405246 238294 405302 238350
rect 404874 238170 404930 238226
rect 404998 238170 405054 238226
rect 405122 238170 405178 238226
rect 405246 238170 405302 238226
rect 404874 238046 404930 238102
rect 404998 238046 405054 238102
rect 405122 238046 405178 238102
rect 405246 238046 405302 238102
rect 404874 237922 404930 237978
rect 404998 237922 405054 237978
rect 405122 237922 405178 237978
rect 405246 237922 405302 237978
rect 404874 220294 404930 220350
rect 404998 220294 405054 220350
rect 405122 220294 405178 220350
rect 405246 220294 405302 220350
rect 404874 220170 404930 220226
rect 404998 220170 405054 220226
rect 405122 220170 405178 220226
rect 405246 220170 405302 220226
rect 404874 220046 404930 220102
rect 404998 220046 405054 220102
rect 405122 220046 405178 220102
rect 405246 220046 405302 220102
rect 404874 219922 404930 219978
rect 404998 219922 405054 219978
rect 405122 219922 405178 219978
rect 405246 219922 405302 219978
rect 404874 202294 404930 202350
rect 404998 202294 405054 202350
rect 405122 202294 405178 202350
rect 405246 202294 405302 202350
rect 404874 202170 404930 202226
rect 404998 202170 405054 202226
rect 405122 202170 405178 202226
rect 405246 202170 405302 202226
rect 404874 202046 404930 202102
rect 404998 202046 405054 202102
rect 405122 202046 405178 202102
rect 405246 202046 405302 202102
rect 404874 201922 404930 201978
rect 404998 201922 405054 201978
rect 405122 201922 405178 201978
rect 405246 201922 405302 201978
rect 404874 184294 404930 184350
rect 404998 184294 405054 184350
rect 405122 184294 405178 184350
rect 405246 184294 405302 184350
rect 404874 184170 404930 184226
rect 404998 184170 405054 184226
rect 405122 184170 405178 184226
rect 405246 184170 405302 184226
rect 404874 184046 404930 184102
rect 404998 184046 405054 184102
rect 405122 184046 405178 184102
rect 405246 184046 405302 184102
rect 404874 183922 404930 183978
rect 404998 183922 405054 183978
rect 405122 183922 405178 183978
rect 405246 183922 405302 183978
rect 404874 166294 404930 166350
rect 404998 166294 405054 166350
rect 405122 166294 405178 166350
rect 405246 166294 405302 166350
rect 404874 166170 404930 166226
rect 404998 166170 405054 166226
rect 405122 166170 405178 166226
rect 405246 166170 405302 166226
rect 404874 166046 404930 166102
rect 404998 166046 405054 166102
rect 405122 166046 405178 166102
rect 405246 166046 405302 166102
rect 404874 165922 404930 165978
rect 404998 165922 405054 165978
rect 405122 165922 405178 165978
rect 405246 165922 405302 165978
rect 404874 148294 404930 148350
rect 404998 148294 405054 148350
rect 405122 148294 405178 148350
rect 405246 148294 405302 148350
rect 404874 148170 404930 148226
rect 404998 148170 405054 148226
rect 405122 148170 405178 148226
rect 405246 148170 405302 148226
rect 404874 148046 404930 148102
rect 404998 148046 405054 148102
rect 405122 148046 405178 148102
rect 405246 148046 405302 148102
rect 404874 147922 404930 147978
rect 404998 147922 405054 147978
rect 405122 147922 405178 147978
rect 405246 147922 405302 147978
rect 404874 130294 404930 130350
rect 404998 130294 405054 130350
rect 405122 130294 405178 130350
rect 405246 130294 405302 130350
rect 404874 130170 404930 130226
rect 404998 130170 405054 130226
rect 405122 130170 405178 130226
rect 405246 130170 405302 130226
rect 404874 130046 404930 130102
rect 404998 130046 405054 130102
rect 405122 130046 405178 130102
rect 405246 130046 405302 130102
rect 404874 129922 404930 129978
rect 404998 129922 405054 129978
rect 405122 129922 405178 129978
rect 405246 129922 405302 129978
rect 377874 118294 377930 118350
rect 377998 118294 378054 118350
rect 378122 118294 378178 118350
rect 378246 118294 378302 118350
rect 377874 118170 377930 118226
rect 377998 118170 378054 118226
rect 378122 118170 378178 118226
rect 378246 118170 378302 118226
rect 377874 118046 377930 118102
rect 377998 118046 378054 118102
rect 378122 118046 378178 118102
rect 378246 118046 378302 118102
rect 377874 117922 377930 117978
rect 377998 117922 378054 117978
rect 378122 117922 378178 117978
rect 378246 117922 378302 117978
rect 408594 406294 408650 406350
rect 408718 406294 408774 406350
rect 408842 406294 408898 406350
rect 408966 406294 409022 406350
rect 408594 406170 408650 406226
rect 408718 406170 408774 406226
rect 408842 406170 408898 406226
rect 408966 406170 409022 406226
rect 408594 406046 408650 406102
rect 408718 406046 408774 406102
rect 408842 406046 408898 406102
rect 408966 406046 409022 406102
rect 408594 405922 408650 405978
rect 408718 405922 408774 405978
rect 408842 405922 408898 405978
rect 408966 405922 409022 405978
rect 408594 388294 408650 388350
rect 408718 388294 408774 388350
rect 408842 388294 408898 388350
rect 408966 388294 409022 388350
rect 408594 388170 408650 388226
rect 408718 388170 408774 388226
rect 408842 388170 408898 388226
rect 408966 388170 409022 388226
rect 408594 388046 408650 388102
rect 408718 388046 408774 388102
rect 408842 388046 408898 388102
rect 408966 388046 409022 388102
rect 408594 387922 408650 387978
rect 408718 387922 408774 387978
rect 408842 387922 408898 387978
rect 408966 387922 409022 387978
rect 408594 370294 408650 370350
rect 408718 370294 408774 370350
rect 408842 370294 408898 370350
rect 408966 370294 409022 370350
rect 408594 370170 408650 370226
rect 408718 370170 408774 370226
rect 408842 370170 408898 370226
rect 408966 370170 409022 370226
rect 408594 370046 408650 370102
rect 408718 370046 408774 370102
rect 408842 370046 408898 370102
rect 408966 370046 409022 370102
rect 408594 369922 408650 369978
rect 408718 369922 408774 369978
rect 408842 369922 408898 369978
rect 408966 369922 409022 369978
rect 408594 352294 408650 352350
rect 408718 352294 408774 352350
rect 408842 352294 408898 352350
rect 408966 352294 409022 352350
rect 408594 352170 408650 352226
rect 408718 352170 408774 352226
rect 408842 352170 408898 352226
rect 408966 352170 409022 352226
rect 408594 352046 408650 352102
rect 408718 352046 408774 352102
rect 408842 352046 408898 352102
rect 408966 352046 409022 352102
rect 408594 351922 408650 351978
rect 408718 351922 408774 351978
rect 408842 351922 408898 351978
rect 408966 351922 409022 351978
rect 435594 400294 435650 400350
rect 435718 400294 435774 400350
rect 435842 400294 435898 400350
rect 435966 400294 436022 400350
rect 435594 400170 435650 400226
rect 435718 400170 435774 400226
rect 435842 400170 435898 400226
rect 435966 400170 436022 400226
rect 435594 400046 435650 400102
rect 435718 400046 435774 400102
rect 435842 400046 435898 400102
rect 435966 400046 436022 400102
rect 435594 399922 435650 399978
rect 435718 399922 435774 399978
rect 435842 399922 435898 399978
rect 435966 399922 436022 399978
rect 435594 382294 435650 382350
rect 435718 382294 435774 382350
rect 435842 382294 435898 382350
rect 435966 382294 436022 382350
rect 435594 382170 435650 382226
rect 435718 382170 435774 382226
rect 435842 382170 435898 382226
rect 435966 382170 436022 382226
rect 435594 382046 435650 382102
rect 435718 382046 435774 382102
rect 435842 382046 435898 382102
rect 435966 382046 436022 382102
rect 435594 381922 435650 381978
rect 435718 381922 435774 381978
rect 435842 381922 435898 381978
rect 435966 381922 436022 381978
rect 435594 364294 435650 364350
rect 435718 364294 435774 364350
rect 435842 364294 435898 364350
rect 435966 364294 436022 364350
rect 435594 364170 435650 364226
rect 435718 364170 435774 364226
rect 435842 364170 435898 364226
rect 435966 364170 436022 364226
rect 435594 364046 435650 364102
rect 435718 364046 435774 364102
rect 435842 364046 435898 364102
rect 435966 364046 436022 364102
rect 435594 363922 435650 363978
rect 435718 363922 435774 363978
rect 435842 363922 435898 363978
rect 435966 363922 436022 363978
rect 435594 346294 435650 346350
rect 435718 346294 435774 346350
rect 435842 346294 435898 346350
rect 435966 346294 436022 346350
rect 435594 346170 435650 346226
rect 435718 346170 435774 346226
rect 435842 346170 435898 346226
rect 435966 346170 436022 346226
rect 435594 346046 435650 346102
rect 435718 346046 435774 346102
rect 435842 346046 435898 346102
rect 435966 346046 436022 346102
rect 435594 345922 435650 345978
rect 435718 345922 435774 345978
rect 435842 345922 435898 345978
rect 435966 345922 436022 345978
rect 408594 334294 408650 334350
rect 408718 334294 408774 334350
rect 408842 334294 408898 334350
rect 408966 334294 409022 334350
rect 408594 334170 408650 334226
rect 408718 334170 408774 334226
rect 408842 334170 408898 334226
rect 408966 334170 409022 334226
rect 408594 334046 408650 334102
rect 408718 334046 408774 334102
rect 408842 334046 408898 334102
rect 408966 334046 409022 334102
rect 408594 333922 408650 333978
rect 408718 333922 408774 333978
rect 408842 333922 408898 333978
rect 408966 333922 409022 333978
rect 408594 316294 408650 316350
rect 408718 316294 408774 316350
rect 408842 316294 408898 316350
rect 408966 316294 409022 316350
rect 408594 316170 408650 316226
rect 408718 316170 408774 316226
rect 408842 316170 408898 316226
rect 408966 316170 409022 316226
rect 408594 316046 408650 316102
rect 408718 316046 408774 316102
rect 408842 316046 408898 316102
rect 408966 316046 409022 316102
rect 408594 315922 408650 315978
rect 408718 315922 408774 315978
rect 408842 315922 408898 315978
rect 408966 315922 409022 315978
rect 408594 298294 408650 298350
rect 408718 298294 408774 298350
rect 408842 298294 408898 298350
rect 408966 298294 409022 298350
rect 408594 298170 408650 298226
rect 408718 298170 408774 298226
rect 408842 298170 408898 298226
rect 408966 298170 409022 298226
rect 408594 298046 408650 298102
rect 408718 298046 408774 298102
rect 408842 298046 408898 298102
rect 408966 298046 409022 298102
rect 408594 297922 408650 297978
rect 408718 297922 408774 297978
rect 408842 297922 408898 297978
rect 408966 297922 409022 297978
rect 408594 280294 408650 280350
rect 408718 280294 408774 280350
rect 408842 280294 408898 280350
rect 408966 280294 409022 280350
rect 408594 280170 408650 280226
rect 408718 280170 408774 280226
rect 408842 280170 408898 280226
rect 408966 280170 409022 280226
rect 408594 280046 408650 280102
rect 408718 280046 408774 280102
rect 408842 280046 408898 280102
rect 408966 280046 409022 280102
rect 408594 279922 408650 279978
rect 408718 279922 408774 279978
rect 408842 279922 408898 279978
rect 408966 279922 409022 279978
rect 408594 262294 408650 262350
rect 408718 262294 408774 262350
rect 408842 262294 408898 262350
rect 408966 262294 409022 262350
rect 408594 262170 408650 262226
rect 408718 262170 408774 262226
rect 408842 262170 408898 262226
rect 408966 262170 409022 262226
rect 408594 262046 408650 262102
rect 408718 262046 408774 262102
rect 408842 262046 408898 262102
rect 408966 262046 409022 262102
rect 408594 261922 408650 261978
rect 408718 261922 408774 261978
rect 408842 261922 408898 261978
rect 408966 261922 409022 261978
rect 408594 244294 408650 244350
rect 408718 244294 408774 244350
rect 408842 244294 408898 244350
rect 408966 244294 409022 244350
rect 408594 244170 408650 244226
rect 408718 244170 408774 244226
rect 408842 244170 408898 244226
rect 408966 244170 409022 244226
rect 408594 244046 408650 244102
rect 408718 244046 408774 244102
rect 408842 244046 408898 244102
rect 408966 244046 409022 244102
rect 408594 243922 408650 243978
rect 408718 243922 408774 243978
rect 408842 243922 408898 243978
rect 408966 243922 409022 243978
rect 408594 226294 408650 226350
rect 408718 226294 408774 226350
rect 408842 226294 408898 226350
rect 408966 226294 409022 226350
rect 408594 226170 408650 226226
rect 408718 226170 408774 226226
rect 408842 226170 408898 226226
rect 408966 226170 409022 226226
rect 408594 226046 408650 226102
rect 408718 226046 408774 226102
rect 408842 226046 408898 226102
rect 408966 226046 409022 226102
rect 408594 225922 408650 225978
rect 408718 225922 408774 225978
rect 408842 225922 408898 225978
rect 408966 225922 409022 225978
rect 408594 208294 408650 208350
rect 408718 208294 408774 208350
rect 408842 208294 408898 208350
rect 408966 208294 409022 208350
rect 408594 208170 408650 208226
rect 408718 208170 408774 208226
rect 408842 208170 408898 208226
rect 408966 208170 409022 208226
rect 408594 208046 408650 208102
rect 408718 208046 408774 208102
rect 408842 208046 408898 208102
rect 408966 208046 409022 208102
rect 408594 207922 408650 207978
rect 408718 207922 408774 207978
rect 408842 207922 408898 207978
rect 408966 207922 409022 207978
rect 408594 190294 408650 190350
rect 408718 190294 408774 190350
rect 408842 190294 408898 190350
rect 408966 190294 409022 190350
rect 408594 190170 408650 190226
rect 408718 190170 408774 190226
rect 408842 190170 408898 190226
rect 408966 190170 409022 190226
rect 408594 190046 408650 190102
rect 408718 190046 408774 190102
rect 408842 190046 408898 190102
rect 408966 190046 409022 190102
rect 408594 189922 408650 189978
rect 408718 189922 408774 189978
rect 408842 189922 408898 189978
rect 408966 189922 409022 189978
rect 408594 172294 408650 172350
rect 408718 172294 408774 172350
rect 408842 172294 408898 172350
rect 408966 172294 409022 172350
rect 408594 172170 408650 172226
rect 408718 172170 408774 172226
rect 408842 172170 408898 172226
rect 408966 172170 409022 172226
rect 408594 172046 408650 172102
rect 408718 172046 408774 172102
rect 408842 172046 408898 172102
rect 408966 172046 409022 172102
rect 408594 171922 408650 171978
rect 408718 171922 408774 171978
rect 408842 171922 408898 171978
rect 408966 171922 409022 171978
rect 408594 154294 408650 154350
rect 408718 154294 408774 154350
rect 408842 154294 408898 154350
rect 408966 154294 409022 154350
rect 408594 154170 408650 154226
rect 408718 154170 408774 154226
rect 408842 154170 408898 154226
rect 408966 154170 409022 154226
rect 408594 154046 408650 154102
rect 408718 154046 408774 154102
rect 408842 154046 408898 154102
rect 408966 154046 409022 154102
rect 408594 153922 408650 153978
rect 408718 153922 408774 153978
rect 408842 153922 408898 153978
rect 408966 153922 409022 153978
rect 408594 136294 408650 136350
rect 408718 136294 408774 136350
rect 408842 136294 408898 136350
rect 408966 136294 409022 136350
rect 408594 136170 408650 136226
rect 408718 136170 408774 136226
rect 408842 136170 408898 136226
rect 408966 136170 409022 136226
rect 408594 136046 408650 136102
rect 408718 136046 408774 136102
rect 408842 136046 408898 136102
rect 408966 136046 409022 136102
rect 408594 135922 408650 135978
rect 408718 135922 408774 135978
rect 408842 135922 408898 135978
rect 408966 135922 409022 135978
rect 408594 118294 408650 118350
rect 408718 118294 408774 118350
rect 408842 118294 408898 118350
rect 408966 118294 409022 118350
rect 408594 118170 408650 118226
rect 408718 118170 408774 118226
rect 408842 118170 408898 118226
rect 408966 118170 409022 118226
rect 408594 118046 408650 118102
rect 408718 118046 408774 118102
rect 408842 118046 408898 118102
rect 408966 118046 409022 118102
rect 408594 117922 408650 117978
rect 408718 117922 408774 117978
rect 408842 117922 408898 117978
rect 408966 117922 409022 117978
rect 364518 112294 364574 112350
rect 364642 112294 364698 112350
rect 364518 112170 364574 112226
rect 364642 112170 364698 112226
rect 364518 112046 364574 112102
rect 364642 112046 364698 112102
rect 364518 111922 364574 111978
rect 364642 111922 364698 111978
rect 395238 112294 395294 112350
rect 395362 112294 395418 112350
rect 395238 112170 395294 112226
rect 395362 112170 395418 112226
rect 395238 112046 395294 112102
rect 395362 112046 395418 112102
rect 395238 111922 395294 111978
rect 395362 111922 395418 111978
rect 379878 100294 379934 100350
rect 380002 100294 380058 100350
rect 379878 100170 379934 100226
rect 380002 100170 380058 100226
rect 379878 100046 379934 100102
rect 380002 100046 380058 100102
rect 379878 99922 379934 99978
rect 380002 99922 380058 99978
rect 410598 100294 410654 100350
rect 410722 100294 410778 100350
rect 410598 100170 410654 100226
rect 410722 100170 410778 100226
rect 410598 100046 410654 100102
rect 410722 100046 410778 100102
rect 410598 99922 410654 99978
rect 410722 99922 410778 99978
rect 364518 94294 364574 94350
rect 364642 94294 364698 94350
rect 364518 94170 364574 94226
rect 364642 94170 364698 94226
rect 364518 94046 364574 94102
rect 364642 94046 364698 94102
rect 364518 93922 364574 93978
rect 364642 93922 364698 93978
rect 395238 94294 395294 94350
rect 395362 94294 395418 94350
rect 395238 94170 395294 94226
rect 395362 94170 395418 94226
rect 395238 94046 395294 94102
rect 395362 94046 395418 94102
rect 395238 93922 395294 93978
rect 395362 93922 395418 93978
rect 379878 82294 379934 82350
rect 380002 82294 380058 82350
rect 379878 82170 379934 82226
rect 380002 82170 380058 82226
rect 379878 82046 379934 82102
rect 380002 82046 380058 82102
rect 379878 81922 379934 81978
rect 380002 81922 380058 81978
rect 410598 82294 410654 82350
rect 410722 82294 410778 82350
rect 410598 82170 410654 82226
rect 410722 82170 410778 82226
rect 410598 82046 410654 82102
rect 410722 82046 410778 82102
rect 410598 81922 410654 81978
rect 410722 81922 410778 81978
rect 364518 76294 364574 76350
rect 364642 76294 364698 76350
rect 364518 76170 364574 76226
rect 364642 76170 364698 76226
rect 364518 76046 364574 76102
rect 364642 76046 364698 76102
rect 364518 75922 364574 75978
rect 364642 75922 364698 75978
rect 395238 76294 395294 76350
rect 395362 76294 395418 76350
rect 395238 76170 395294 76226
rect 395362 76170 395418 76226
rect 395238 76046 395294 76102
rect 395362 76046 395418 76102
rect 395238 75922 395294 75978
rect 395362 75922 395418 75978
rect 379878 64294 379934 64350
rect 380002 64294 380058 64350
rect 379878 64170 379934 64226
rect 380002 64170 380058 64226
rect 379878 64046 379934 64102
rect 380002 64046 380058 64102
rect 379878 63922 379934 63978
rect 380002 63922 380058 63978
rect 410598 64294 410654 64350
rect 410722 64294 410778 64350
rect 410598 64170 410654 64226
rect 410722 64170 410778 64226
rect 410598 64046 410654 64102
rect 410722 64046 410778 64102
rect 410598 63922 410654 63978
rect 410722 63922 410778 63978
rect 364518 58294 364574 58350
rect 364642 58294 364698 58350
rect 364518 58170 364574 58226
rect 364642 58170 364698 58226
rect 364518 58046 364574 58102
rect 364642 58046 364698 58102
rect 364518 57922 364574 57978
rect 364642 57922 364698 57978
rect 395238 58294 395294 58350
rect 395362 58294 395418 58350
rect 395238 58170 395294 58226
rect 395362 58170 395418 58226
rect 395238 58046 395294 58102
rect 395362 58046 395418 58102
rect 395238 57922 395294 57978
rect 395362 57922 395418 57978
rect 374154 40294 374210 40350
rect 374278 40294 374334 40350
rect 374402 40294 374458 40350
rect 374526 40294 374582 40350
rect 374154 40170 374210 40226
rect 374278 40170 374334 40226
rect 374402 40170 374458 40226
rect 374526 40170 374582 40226
rect 374154 40046 374210 40102
rect 374278 40046 374334 40102
rect 374402 40046 374458 40102
rect 374526 40046 374582 40102
rect 374154 39922 374210 39978
rect 374278 39922 374334 39978
rect 374402 39922 374458 39978
rect 374526 39922 374582 39978
rect 374154 22294 374210 22350
rect 374278 22294 374334 22350
rect 374402 22294 374458 22350
rect 374526 22294 374582 22350
rect 374154 22170 374210 22226
rect 374278 22170 374334 22226
rect 374402 22170 374458 22226
rect 374526 22170 374582 22226
rect 374154 22046 374210 22102
rect 374278 22046 374334 22102
rect 374402 22046 374458 22102
rect 374526 22046 374582 22102
rect 374154 21922 374210 21978
rect 374278 21922 374334 21978
rect 374402 21922 374458 21978
rect 374526 21922 374582 21978
rect 347154 -1176 347210 -1120
rect 347278 -1176 347334 -1120
rect 347402 -1176 347458 -1120
rect 347526 -1176 347582 -1120
rect 347154 -1300 347210 -1244
rect 347278 -1300 347334 -1244
rect 347402 -1300 347458 -1244
rect 347526 -1300 347582 -1244
rect 347154 -1424 347210 -1368
rect 347278 -1424 347334 -1368
rect 347402 -1424 347458 -1368
rect 347526 -1424 347582 -1368
rect 347154 -1548 347210 -1492
rect 347278 -1548 347334 -1492
rect 347402 -1548 347458 -1492
rect 347526 -1548 347582 -1492
rect 374154 4294 374210 4350
rect 374278 4294 374334 4350
rect 374402 4294 374458 4350
rect 374526 4294 374582 4350
rect 374154 4170 374210 4226
rect 374278 4170 374334 4226
rect 374402 4170 374458 4226
rect 374526 4170 374582 4226
rect 374154 4046 374210 4102
rect 374278 4046 374334 4102
rect 374402 4046 374458 4102
rect 374526 4046 374582 4102
rect 374154 3922 374210 3978
rect 374278 3922 374334 3978
rect 374402 3922 374458 3978
rect 374526 3922 374582 3978
rect 374154 -216 374210 -160
rect 374278 -216 374334 -160
rect 374402 -216 374458 -160
rect 374526 -216 374582 -160
rect 374154 -340 374210 -284
rect 374278 -340 374334 -284
rect 374402 -340 374458 -284
rect 374526 -340 374582 -284
rect 374154 -464 374210 -408
rect 374278 -464 374334 -408
rect 374402 -464 374458 -408
rect 374526 -464 374582 -408
rect 374154 -588 374210 -532
rect 374278 -588 374334 -532
rect 374402 -588 374458 -532
rect 374526 -588 374582 -532
rect 377874 46294 377930 46350
rect 377998 46294 378054 46350
rect 378122 46294 378178 46350
rect 378246 46294 378302 46350
rect 377874 46170 377930 46226
rect 377998 46170 378054 46226
rect 378122 46170 378178 46226
rect 378246 46170 378302 46226
rect 377874 46046 377930 46102
rect 377998 46046 378054 46102
rect 378122 46046 378178 46102
rect 378246 46046 378302 46102
rect 377874 45922 377930 45978
rect 377998 45922 378054 45978
rect 378122 45922 378178 45978
rect 378246 45922 378302 45978
rect 377874 28294 377930 28350
rect 377998 28294 378054 28350
rect 378122 28294 378178 28350
rect 378246 28294 378302 28350
rect 377874 28170 377930 28226
rect 377998 28170 378054 28226
rect 378122 28170 378178 28226
rect 378246 28170 378302 28226
rect 377874 28046 377930 28102
rect 377998 28046 378054 28102
rect 378122 28046 378178 28102
rect 378246 28046 378302 28102
rect 377874 27922 377930 27978
rect 377998 27922 378054 27978
rect 378122 27922 378178 27978
rect 378246 27922 378302 27978
rect 377874 10294 377930 10350
rect 377998 10294 378054 10350
rect 378122 10294 378178 10350
rect 378246 10294 378302 10350
rect 377874 10170 377930 10226
rect 377998 10170 378054 10226
rect 378122 10170 378178 10226
rect 378246 10170 378302 10226
rect 377874 10046 377930 10102
rect 377998 10046 378054 10102
rect 378122 10046 378178 10102
rect 378246 10046 378302 10102
rect 377874 9922 377930 9978
rect 377998 9922 378054 9978
rect 378122 9922 378178 9978
rect 378246 9922 378302 9978
rect 377874 -1176 377930 -1120
rect 377998 -1176 378054 -1120
rect 378122 -1176 378178 -1120
rect 378246 -1176 378302 -1120
rect 377874 -1300 377930 -1244
rect 377998 -1300 378054 -1244
rect 378122 -1300 378178 -1244
rect 378246 -1300 378302 -1244
rect 377874 -1424 377930 -1368
rect 377998 -1424 378054 -1368
rect 378122 -1424 378178 -1368
rect 378246 -1424 378302 -1368
rect 377874 -1548 377930 -1492
rect 377998 -1548 378054 -1492
rect 378122 -1548 378178 -1492
rect 378246 -1548 378302 -1492
rect 404874 40294 404930 40350
rect 404998 40294 405054 40350
rect 405122 40294 405178 40350
rect 405246 40294 405302 40350
rect 404874 40170 404930 40226
rect 404998 40170 405054 40226
rect 405122 40170 405178 40226
rect 405246 40170 405302 40226
rect 404874 40046 404930 40102
rect 404998 40046 405054 40102
rect 405122 40046 405178 40102
rect 405246 40046 405302 40102
rect 404874 39922 404930 39978
rect 404998 39922 405054 39978
rect 405122 39922 405178 39978
rect 405246 39922 405302 39978
rect 404874 22294 404930 22350
rect 404998 22294 405054 22350
rect 405122 22294 405178 22350
rect 405246 22294 405302 22350
rect 404874 22170 404930 22226
rect 404998 22170 405054 22226
rect 405122 22170 405178 22226
rect 405246 22170 405302 22226
rect 404874 22046 404930 22102
rect 404998 22046 405054 22102
rect 405122 22046 405178 22102
rect 405246 22046 405302 22102
rect 404874 21922 404930 21978
rect 404998 21922 405054 21978
rect 405122 21922 405178 21978
rect 405246 21922 405302 21978
rect 404874 4294 404930 4350
rect 404998 4294 405054 4350
rect 405122 4294 405178 4350
rect 405246 4294 405302 4350
rect 404874 4170 404930 4226
rect 404998 4170 405054 4226
rect 405122 4170 405178 4226
rect 405246 4170 405302 4226
rect 404874 4046 404930 4102
rect 404998 4046 405054 4102
rect 405122 4046 405178 4102
rect 405246 4046 405302 4102
rect 404874 3922 404930 3978
rect 404998 3922 405054 3978
rect 405122 3922 405178 3978
rect 405246 3922 405302 3978
rect 404874 -216 404930 -160
rect 404998 -216 405054 -160
rect 405122 -216 405178 -160
rect 405246 -216 405302 -160
rect 404874 -340 404930 -284
rect 404998 -340 405054 -284
rect 405122 -340 405178 -284
rect 405246 -340 405302 -284
rect 404874 -464 404930 -408
rect 404998 -464 405054 -408
rect 405122 -464 405178 -408
rect 405246 -464 405302 -408
rect 404874 -588 404930 -532
rect 404998 -588 405054 -532
rect 405122 -588 405178 -532
rect 405246 -588 405302 -532
rect 408594 46294 408650 46350
rect 408718 46294 408774 46350
rect 408842 46294 408898 46350
rect 408966 46294 409022 46350
rect 408594 46170 408650 46226
rect 408718 46170 408774 46226
rect 408842 46170 408898 46226
rect 408966 46170 409022 46226
rect 408594 46046 408650 46102
rect 408718 46046 408774 46102
rect 408842 46046 408898 46102
rect 408966 46046 409022 46102
rect 408594 45922 408650 45978
rect 408718 45922 408774 45978
rect 408842 45922 408898 45978
rect 408966 45922 409022 45978
rect 408594 28294 408650 28350
rect 408718 28294 408774 28350
rect 408842 28294 408898 28350
rect 408966 28294 409022 28350
rect 408594 28170 408650 28226
rect 408718 28170 408774 28226
rect 408842 28170 408898 28226
rect 408966 28170 409022 28226
rect 408594 28046 408650 28102
rect 408718 28046 408774 28102
rect 408842 28046 408898 28102
rect 408966 28046 409022 28102
rect 408594 27922 408650 27978
rect 408718 27922 408774 27978
rect 408842 27922 408898 27978
rect 408966 27922 409022 27978
rect 408594 10294 408650 10350
rect 408718 10294 408774 10350
rect 408842 10294 408898 10350
rect 408966 10294 409022 10350
rect 408594 10170 408650 10226
rect 408718 10170 408774 10226
rect 408842 10170 408898 10226
rect 408966 10170 409022 10226
rect 408594 10046 408650 10102
rect 408718 10046 408774 10102
rect 408842 10046 408898 10102
rect 408966 10046 409022 10102
rect 408594 9922 408650 9978
rect 408718 9922 408774 9978
rect 408842 9922 408898 9978
rect 408966 9922 409022 9978
rect 435594 328294 435650 328350
rect 435718 328294 435774 328350
rect 435842 328294 435898 328350
rect 435966 328294 436022 328350
rect 435594 328170 435650 328226
rect 435718 328170 435774 328226
rect 435842 328170 435898 328226
rect 435966 328170 436022 328226
rect 435594 328046 435650 328102
rect 435718 328046 435774 328102
rect 435842 328046 435898 328102
rect 435966 328046 436022 328102
rect 435594 327922 435650 327978
rect 435718 327922 435774 327978
rect 435842 327922 435898 327978
rect 435966 327922 436022 327978
rect 439314 406294 439370 406350
rect 439438 406294 439494 406350
rect 439562 406294 439618 406350
rect 439686 406294 439742 406350
rect 439314 406170 439370 406226
rect 439438 406170 439494 406226
rect 439562 406170 439618 406226
rect 439686 406170 439742 406226
rect 439314 406046 439370 406102
rect 439438 406046 439494 406102
rect 439562 406046 439618 406102
rect 439686 406046 439742 406102
rect 439314 405922 439370 405978
rect 439438 405922 439494 405978
rect 439562 405922 439618 405978
rect 439686 405922 439742 405978
rect 439314 388294 439370 388350
rect 439438 388294 439494 388350
rect 439562 388294 439618 388350
rect 439686 388294 439742 388350
rect 439314 388170 439370 388226
rect 439438 388170 439494 388226
rect 439562 388170 439618 388226
rect 439686 388170 439742 388226
rect 439314 388046 439370 388102
rect 439438 388046 439494 388102
rect 439562 388046 439618 388102
rect 439686 388046 439742 388102
rect 439314 387922 439370 387978
rect 439438 387922 439494 387978
rect 439562 387922 439618 387978
rect 439686 387922 439742 387978
rect 466314 400294 466370 400350
rect 466438 400294 466494 400350
rect 466562 400294 466618 400350
rect 466686 400294 466742 400350
rect 466314 400170 466370 400226
rect 466438 400170 466494 400226
rect 466562 400170 466618 400226
rect 466686 400170 466742 400226
rect 466314 400046 466370 400102
rect 466438 400046 466494 400102
rect 466562 400046 466618 400102
rect 466686 400046 466742 400102
rect 466314 399922 466370 399978
rect 466438 399922 466494 399978
rect 466562 399922 466618 399978
rect 466686 399922 466742 399978
rect 439314 370294 439370 370350
rect 439438 370294 439494 370350
rect 439562 370294 439618 370350
rect 439686 370294 439742 370350
rect 439314 370170 439370 370226
rect 439438 370170 439494 370226
rect 439562 370170 439618 370226
rect 439686 370170 439742 370226
rect 439314 370046 439370 370102
rect 439438 370046 439494 370102
rect 439562 370046 439618 370102
rect 439686 370046 439742 370102
rect 439314 369922 439370 369978
rect 439438 369922 439494 369978
rect 439562 369922 439618 369978
rect 439686 369922 439742 369978
rect 439314 352294 439370 352350
rect 439438 352294 439494 352350
rect 439562 352294 439618 352350
rect 439686 352294 439742 352350
rect 439314 352170 439370 352226
rect 439438 352170 439494 352226
rect 439562 352170 439618 352226
rect 439686 352170 439742 352226
rect 439314 352046 439370 352102
rect 439438 352046 439494 352102
rect 439562 352046 439618 352102
rect 439686 352046 439742 352102
rect 439314 351922 439370 351978
rect 439438 351922 439494 351978
rect 439562 351922 439618 351978
rect 439686 351922 439742 351978
rect 439314 334294 439370 334350
rect 439438 334294 439494 334350
rect 439562 334294 439618 334350
rect 439686 334294 439742 334350
rect 439314 334170 439370 334226
rect 439438 334170 439494 334226
rect 439562 334170 439618 334226
rect 439686 334170 439742 334226
rect 439314 334046 439370 334102
rect 439438 334046 439494 334102
rect 439562 334046 439618 334102
rect 439686 334046 439742 334102
rect 439314 333922 439370 333978
rect 439438 333922 439494 333978
rect 439562 333922 439618 333978
rect 439686 333922 439742 333978
rect 435594 310294 435650 310350
rect 435718 310294 435774 310350
rect 435842 310294 435898 310350
rect 435966 310294 436022 310350
rect 435594 310170 435650 310226
rect 435718 310170 435774 310226
rect 435842 310170 435898 310226
rect 435966 310170 436022 310226
rect 435594 310046 435650 310102
rect 435718 310046 435774 310102
rect 435842 310046 435898 310102
rect 435966 310046 436022 310102
rect 435594 309922 435650 309978
rect 435718 309922 435774 309978
rect 435842 309922 435898 309978
rect 435966 309922 436022 309978
rect 435594 292294 435650 292350
rect 435718 292294 435774 292350
rect 435842 292294 435898 292350
rect 435966 292294 436022 292350
rect 435594 292170 435650 292226
rect 435718 292170 435774 292226
rect 435842 292170 435898 292226
rect 435966 292170 436022 292226
rect 435594 292046 435650 292102
rect 435718 292046 435774 292102
rect 435842 292046 435898 292102
rect 435966 292046 436022 292102
rect 435594 291922 435650 291978
rect 435718 291922 435774 291978
rect 435842 291922 435898 291978
rect 435966 291922 436022 291978
rect 435594 274294 435650 274350
rect 435718 274294 435774 274350
rect 435842 274294 435898 274350
rect 435966 274294 436022 274350
rect 435594 274170 435650 274226
rect 435718 274170 435774 274226
rect 435842 274170 435898 274226
rect 435966 274170 436022 274226
rect 435594 274046 435650 274102
rect 435718 274046 435774 274102
rect 435842 274046 435898 274102
rect 435966 274046 436022 274102
rect 435594 273922 435650 273978
rect 435718 273922 435774 273978
rect 435842 273922 435898 273978
rect 435966 273922 436022 273978
rect 435594 256294 435650 256350
rect 435718 256294 435774 256350
rect 435842 256294 435898 256350
rect 435966 256294 436022 256350
rect 435594 256170 435650 256226
rect 435718 256170 435774 256226
rect 435842 256170 435898 256226
rect 435966 256170 436022 256226
rect 435594 256046 435650 256102
rect 435718 256046 435774 256102
rect 435842 256046 435898 256102
rect 435966 256046 436022 256102
rect 435594 255922 435650 255978
rect 435718 255922 435774 255978
rect 435842 255922 435898 255978
rect 435966 255922 436022 255978
rect 435594 238294 435650 238350
rect 435718 238294 435774 238350
rect 435842 238294 435898 238350
rect 435966 238294 436022 238350
rect 435594 238170 435650 238226
rect 435718 238170 435774 238226
rect 435842 238170 435898 238226
rect 435966 238170 436022 238226
rect 435594 238046 435650 238102
rect 435718 238046 435774 238102
rect 435842 238046 435898 238102
rect 435966 238046 436022 238102
rect 435594 237922 435650 237978
rect 435718 237922 435774 237978
rect 435842 237922 435898 237978
rect 435966 237922 436022 237978
rect 435594 220294 435650 220350
rect 435718 220294 435774 220350
rect 435842 220294 435898 220350
rect 435966 220294 436022 220350
rect 435594 220170 435650 220226
rect 435718 220170 435774 220226
rect 435842 220170 435898 220226
rect 435966 220170 436022 220226
rect 435594 220046 435650 220102
rect 435718 220046 435774 220102
rect 435842 220046 435898 220102
rect 435966 220046 436022 220102
rect 435594 219922 435650 219978
rect 435718 219922 435774 219978
rect 435842 219922 435898 219978
rect 435966 219922 436022 219978
rect 435594 202294 435650 202350
rect 435718 202294 435774 202350
rect 435842 202294 435898 202350
rect 435966 202294 436022 202350
rect 435594 202170 435650 202226
rect 435718 202170 435774 202226
rect 435842 202170 435898 202226
rect 435966 202170 436022 202226
rect 435594 202046 435650 202102
rect 435718 202046 435774 202102
rect 435842 202046 435898 202102
rect 435966 202046 436022 202102
rect 435594 201922 435650 201978
rect 435718 201922 435774 201978
rect 435842 201922 435898 201978
rect 435966 201922 436022 201978
rect 435594 184294 435650 184350
rect 435718 184294 435774 184350
rect 435842 184294 435898 184350
rect 435966 184294 436022 184350
rect 435594 184170 435650 184226
rect 435718 184170 435774 184226
rect 435842 184170 435898 184226
rect 435966 184170 436022 184226
rect 435594 184046 435650 184102
rect 435718 184046 435774 184102
rect 435842 184046 435898 184102
rect 435966 184046 436022 184102
rect 435594 183922 435650 183978
rect 435718 183922 435774 183978
rect 435842 183922 435898 183978
rect 435966 183922 436022 183978
rect 435594 166294 435650 166350
rect 435718 166294 435774 166350
rect 435842 166294 435898 166350
rect 435966 166294 436022 166350
rect 435594 166170 435650 166226
rect 435718 166170 435774 166226
rect 435842 166170 435898 166226
rect 435966 166170 436022 166226
rect 435594 166046 435650 166102
rect 435718 166046 435774 166102
rect 435842 166046 435898 166102
rect 435966 166046 436022 166102
rect 435594 165922 435650 165978
rect 435718 165922 435774 165978
rect 435842 165922 435898 165978
rect 435966 165922 436022 165978
rect 435594 148294 435650 148350
rect 435718 148294 435774 148350
rect 435842 148294 435898 148350
rect 435966 148294 436022 148350
rect 435594 148170 435650 148226
rect 435718 148170 435774 148226
rect 435842 148170 435898 148226
rect 435966 148170 436022 148226
rect 435594 148046 435650 148102
rect 435718 148046 435774 148102
rect 435842 148046 435898 148102
rect 435966 148046 436022 148102
rect 435594 147922 435650 147978
rect 435718 147922 435774 147978
rect 435842 147922 435898 147978
rect 435966 147922 436022 147978
rect 435594 130294 435650 130350
rect 435718 130294 435774 130350
rect 435842 130294 435898 130350
rect 435966 130294 436022 130350
rect 435594 130170 435650 130226
rect 435718 130170 435774 130226
rect 435842 130170 435898 130226
rect 435966 130170 436022 130226
rect 435594 130046 435650 130102
rect 435718 130046 435774 130102
rect 435842 130046 435898 130102
rect 435966 130046 436022 130102
rect 435594 129922 435650 129978
rect 435718 129922 435774 129978
rect 435842 129922 435898 129978
rect 435966 129922 436022 129978
rect 464492 384362 464548 384418
rect 439314 316294 439370 316350
rect 439438 316294 439494 316350
rect 439562 316294 439618 316350
rect 439686 316294 439742 316350
rect 439314 316170 439370 316226
rect 439438 316170 439494 316226
rect 439562 316170 439618 316226
rect 439686 316170 439742 316226
rect 439314 316046 439370 316102
rect 439438 316046 439494 316102
rect 439562 316046 439618 316102
rect 439686 316046 439742 316102
rect 439314 315922 439370 315978
rect 439438 315922 439494 315978
rect 439562 315922 439618 315978
rect 439686 315922 439742 315978
rect 439314 298294 439370 298350
rect 439438 298294 439494 298350
rect 439562 298294 439618 298350
rect 439686 298294 439742 298350
rect 439314 298170 439370 298226
rect 439438 298170 439494 298226
rect 439562 298170 439618 298226
rect 439686 298170 439742 298226
rect 439314 298046 439370 298102
rect 439438 298046 439494 298102
rect 439562 298046 439618 298102
rect 439686 298046 439742 298102
rect 439314 297922 439370 297978
rect 439438 297922 439494 297978
rect 439562 297922 439618 297978
rect 439686 297922 439742 297978
rect 439314 280294 439370 280350
rect 439438 280294 439494 280350
rect 439562 280294 439618 280350
rect 439686 280294 439742 280350
rect 439314 280170 439370 280226
rect 439438 280170 439494 280226
rect 439562 280170 439618 280226
rect 439686 280170 439742 280226
rect 439314 280046 439370 280102
rect 439438 280046 439494 280102
rect 439562 280046 439618 280102
rect 439686 280046 439742 280102
rect 439314 279922 439370 279978
rect 439438 279922 439494 279978
rect 439562 279922 439618 279978
rect 439686 279922 439742 279978
rect 439314 262294 439370 262350
rect 439438 262294 439494 262350
rect 439562 262294 439618 262350
rect 439686 262294 439742 262350
rect 439314 262170 439370 262226
rect 439438 262170 439494 262226
rect 439562 262170 439618 262226
rect 439686 262170 439742 262226
rect 439314 262046 439370 262102
rect 439438 262046 439494 262102
rect 439562 262046 439618 262102
rect 439686 262046 439742 262102
rect 439314 261922 439370 261978
rect 439438 261922 439494 261978
rect 439562 261922 439618 261978
rect 439686 261922 439742 261978
rect 439314 244294 439370 244350
rect 439438 244294 439494 244350
rect 439562 244294 439618 244350
rect 439686 244294 439742 244350
rect 439314 244170 439370 244226
rect 439438 244170 439494 244226
rect 439562 244170 439618 244226
rect 439686 244170 439742 244226
rect 439314 244046 439370 244102
rect 439438 244046 439494 244102
rect 439562 244046 439618 244102
rect 439686 244046 439742 244102
rect 439314 243922 439370 243978
rect 439438 243922 439494 243978
rect 439562 243922 439618 243978
rect 439686 243922 439742 243978
rect 439314 226294 439370 226350
rect 439438 226294 439494 226350
rect 439562 226294 439618 226350
rect 439686 226294 439742 226350
rect 439314 226170 439370 226226
rect 439438 226170 439494 226226
rect 439562 226170 439618 226226
rect 439686 226170 439742 226226
rect 439314 226046 439370 226102
rect 439438 226046 439494 226102
rect 439562 226046 439618 226102
rect 439686 226046 439742 226102
rect 439314 225922 439370 225978
rect 439438 225922 439494 225978
rect 439562 225922 439618 225978
rect 439686 225922 439742 225978
rect 439314 208294 439370 208350
rect 439438 208294 439494 208350
rect 439562 208294 439618 208350
rect 439686 208294 439742 208350
rect 439314 208170 439370 208226
rect 439438 208170 439494 208226
rect 439562 208170 439618 208226
rect 439686 208170 439742 208226
rect 439314 208046 439370 208102
rect 439438 208046 439494 208102
rect 439562 208046 439618 208102
rect 439686 208046 439742 208102
rect 439314 207922 439370 207978
rect 439438 207922 439494 207978
rect 439562 207922 439618 207978
rect 439686 207922 439742 207978
rect 439314 190294 439370 190350
rect 439438 190294 439494 190350
rect 439562 190294 439618 190350
rect 439686 190294 439742 190350
rect 439314 190170 439370 190226
rect 439438 190170 439494 190226
rect 439562 190170 439618 190226
rect 439686 190170 439742 190226
rect 439314 190046 439370 190102
rect 439438 190046 439494 190102
rect 439562 190046 439618 190102
rect 439686 190046 439742 190102
rect 439314 189922 439370 189978
rect 439438 189922 439494 189978
rect 439562 189922 439618 189978
rect 439686 189922 439742 189978
rect 439314 172294 439370 172350
rect 439438 172294 439494 172350
rect 439562 172294 439618 172350
rect 439686 172294 439742 172350
rect 439314 172170 439370 172226
rect 439438 172170 439494 172226
rect 439562 172170 439618 172226
rect 439686 172170 439742 172226
rect 439314 172046 439370 172102
rect 439438 172046 439494 172102
rect 439562 172046 439618 172102
rect 439686 172046 439742 172102
rect 439314 171922 439370 171978
rect 439438 171922 439494 171978
rect 439562 171922 439618 171978
rect 439686 171922 439742 171978
rect 439314 154294 439370 154350
rect 439438 154294 439494 154350
rect 439562 154294 439618 154350
rect 439686 154294 439742 154350
rect 439314 154170 439370 154226
rect 439438 154170 439494 154226
rect 439562 154170 439618 154226
rect 439686 154170 439742 154226
rect 439314 154046 439370 154102
rect 439438 154046 439494 154102
rect 439562 154046 439618 154102
rect 439686 154046 439742 154102
rect 439314 153922 439370 153978
rect 439438 153922 439494 153978
rect 439562 153922 439618 153978
rect 439686 153922 439742 153978
rect 439314 136294 439370 136350
rect 439438 136294 439494 136350
rect 439562 136294 439618 136350
rect 439686 136294 439742 136350
rect 439314 136170 439370 136226
rect 439438 136170 439494 136226
rect 439562 136170 439618 136226
rect 439686 136170 439742 136226
rect 439314 136046 439370 136102
rect 439438 136046 439494 136102
rect 439562 136046 439618 136102
rect 439686 136046 439742 136102
rect 439314 135922 439370 135978
rect 439438 135922 439494 135978
rect 439562 135922 439618 135978
rect 439686 135922 439742 135978
rect 439314 118294 439370 118350
rect 439438 118294 439494 118350
rect 439562 118294 439618 118350
rect 439686 118294 439742 118350
rect 439314 118170 439370 118226
rect 439438 118170 439494 118226
rect 439562 118170 439618 118226
rect 439686 118170 439742 118226
rect 439314 118046 439370 118102
rect 439438 118046 439494 118102
rect 439562 118046 439618 118102
rect 439686 118046 439742 118102
rect 439314 117922 439370 117978
rect 439438 117922 439494 117978
rect 439562 117922 439618 117978
rect 439686 117922 439742 117978
rect 435594 112294 435650 112350
rect 435718 112294 435774 112350
rect 435842 112294 435898 112350
rect 435966 112294 436022 112350
rect 435594 112170 435650 112226
rect 435718 112170 435774 112226
rect 435842 112170 435898 112226
rect 435966 112170 436022 112226
rect 435594 112046 435650 112102
rect 435718 112046 435774 112102
rect 435842 112046 435898 112102
rect 435966 112046 436022 112102
rect 435594 111922 435650 111978
rect 435718 111922 435774 111978
rect 435842 111922 435898 111978
rect 435966 111922 436022 111978
rect 435594 94294 435650 94350
rect 435718 94294 435774 94350
rect 435842 94294 435898 94350
rect 435966 94294 436022 94350
rect 435594 94170 435650 94226
rect 435718 94170 435774 94226
rect 435842 94170 435898 94226
rect 435966 94170 436022 94226
rect 435594 94046 435650 94102
rect 435718 94046 435774 94102
rect 435842 94046 435898 94102
rect 435966 94046 436022 94102
rect 435594 93922 435650 93978
rect 435718 93922 435774 93978
rect 435842 93922 435898 93978
rect 435966 93922 436022 93978
rect 435594 76294 435650 76350
rect 435718 76294 435774 76350
rect 435842 76294 435898 76350
rect 435966 76294 436022 76350
rect 435594 76170 435650 76226
rect 435718 76170 435774 76226
rect 435842 76170 435898 76226
rect 435966 76170 436022 76226
rect 435594 76046 435650 76102
rect 435718 76046 435774 76102
rect 435842 76046 435898 76102
rect 435966 76046 436022 76102
rect 435594 75922 435650 75978
rect 435718 75922 435774 75978
rect 435842 75922 435898 75978
rect 435966 75922 436022 75978
rect 435594 58294 435650 58350
rect 435718 58294 435774 58350
rect 435842 58294 435898 58350
rect 435966 58294 436022 58350
rect 435594 58170 435650 58226
rect 435718 58170 435774 58226
rect 435842 58170 435898 58226
rect 435966 58170 436022 58226
rect 435594 58046 435650 58102
rect 435718 58046 435774 58102
rect 435842 58046 435898 58102
rect 435966 58046 436022 58102
rect 435594 57922 435650 57978
rect 435718 57922 435774 57978
rect 435842 57922 435898 57978
rect 435966 57922 436022 57978
rect 435594 40294 435650 40350
rect 435718 40294 435774 40350
rect 435842 40294 435898 40350
rect 435966 40294 436022 40350
rect 435594 40170 435650 40226
rect 435718 40170 435774 40226
rect 435842 40170 435898 40226
rect 435966 40170 436022 40226
rect 435594 40046 435650 40102
rect 435718 40046 435774 40102
rect 435842 40046 435898 40102
rect 435966 40046 436022 40102
rect 435594 39922 435650 39978
rect 435718 39922 435774 39978
rect 435842 39922 435898 39978
rect 435966 39922 436022 39978
rect 435594 22294 435650 22350
rect 435718 22294 435774 22350
rect 435842 22294 435898 22350
rect 435966 22294 436022 22350
rect 435594 22170 435650 22226
rect 435718 22170 435774 22226
rect 435842 22170 435898 22226
rect 435966 22170 436022 22226
rect 435594 22046 435650 22102
rect 435718 22046 435774 22102
rect 435842 22046 435898 22102
rect 435966 22046 436022 22102
rect 435594 21922 435650 21978
rect 435718 21922 435774 21978
rect 435842 21922 435898 21978
rect 435966 21922 436022 21978
rect 408594 -1176 408650 -1120
rect 408718 -1176 408774 -1120
rect 408842 -1176 408898 -1120
rect 408966 -1176 409022 -1120
rect 408594 -1300 408650 -1244
rect 408718 -1300 408774 -1244
rect 408842 -1300 408898 -1244
rect 408966 -1300 409022 -1244
rect 408594 -1424 408650 -1368
rect 408718 -1424 408774 -1368
rect 408842 -1424 408898 -1368
rect 408966 -1424 409022 -1368
rect 408594 -1548 408650 -1492
rect 408718 -1548 408774 -1492
rect 408842 -1548 408898 -1492
rect 408966 -1548 409022 -1492
rect 435594 4294 435650 4350
rect 435718 4294 435774 4350
rect 435842 4294 435898 4350
rect 435966 4294 436022 4350
rect 435594 4170 435650 4226
rect 435718 4170 435774 4226
rect 435842 4170 435898 4226
rect 435966 4170 436022 4226
rect 435594 4046 435650 4102
rect 435718 4046 435774 4102
rect 435842 4046 435898 4102
rect 435966 4046 436022 4102
rect 435594 3922 435650 3978
rect 435718 3922 435774 3978
rect 435842 3922 435898 3978
rect 435966 3922 436022 3978
rect 435594 -216 435650 -160
rect 435718 -216 435774 -160
rect 435842 -216 435898 -160
rect 435966 -216 436022 -160
rect 435594 -340 435650 -284
rect 435718 -340 435774 -284
rect 435842 -340 435898 -284
rect 435966 -340 436022 -284
rect 435594 -464 435650 -408
rect 435718 -464 435774 -408
rect 435842 -464 435898 -408
rect 435966 -464 436022 -408
rect 435594 -588 435650 -532
rect 435718 -588 435774 -532
rect 435842 -588 435898 -532
rect 435966 -588 436022 -532
rect 439314 100294 439370 100350
rect 439438 100294 439494 100350
rect 439562 100294 439618 100350
rect 439686 100294 439742 100350
rect 439314 100170 439370 100226
rect 439438 100170 439494 100226
rect 439562 100170 439618 100226
rect 439686 100170 439742 100226
rect 439314 100046 439370 100102
rect 439438 100046 439494 100102
rect 439562 100046 439618 100102
rect 439686 100046 439742 100102
rect 439314 99922 439370 99978
rect 439438 99922 439494 99978
rect 439562 99922 439618 99978
rect 439686 99922 439742 99978
rect 439314 82294 439370 82350
rect 439438 82294 439494 82350
rect 439562 82294 439618 82350
rect 439686 82294 439742 82350
rect 439314 82170 439370 82226
rect 439438 82170 439494 82226
rect 439562 82170 439618 82226
rect 439686 82170 439742 82226
rect 439314 82046 439370 82102
rect 439438 82046 439494 82102
rect 439562 82046 439618 82102
rect 439686 82046 439742 82102
rect 439314 81922 439370 81978
rect 439438 81922 439494 81978
rect 439562 81922 439618 81978
rect 439686 81922 439742 81978
rect 439314 64294 439370 64350
rect 439438 64294 439494 64350
rect 439562 64294 439618 64350
rect 439686 64294 439742 64350
rect 439314 64170 439370 64226
rect 439438 64170 439494 64226
rect 439562 64170 439618 64226
rect 439686 64170 439742 64226
rect 439314 64046 439370 64102
rect 439438 64046 439494 64102
rect 439562 64046 439618 64102
rect 439686 64046 439742 64102
rect 439314 63922 439370 63978
rect 439438 63922 439494 63978
rect 439562 63922 439618 63978
rect 439686 63922 439742 63978
rect 464492 198062 464548 198118
rect 466314 382294 466370 382350
rect 466438 382294 466494 382350
rect 466562 382294 466618 382350
rect 466686 382294 466742 382350
rect 466314 382170 466370 382226
rect 466438 382170 466494 382226
rect 466562 382170 466618 382226
rect 466686 382170 466742 382226
rect 466314 382046 466370 382102
rect 466438 382046 466494 382102
rect 466562 382046 466618 382102
rect 466686 382046 466742 382102
rect 466314 381922 466370 381978
rect 466438 381922 466494 381978
rect 466562 381922 466618 381978
rect 466686 381922 466742 381978
rect 466314 364294 466370 364350
rect 466438 364294 466494 364350
rect 466562 364294 466618 364350
rect 466686 364294 466742 364350
rect 466314 364170 466370 364226
rect 466438 364170 466494 364226
rect 466562 364170 466618 364226
rect 466686 364170 466742 364226
rect 466314 364046 466370 364102
rect 466438 364046 466494 364102
rect 466562 364046 466618 364102
rect 466686 364046 466742 364102
rect 466314 363922 466370 363978
rect 466438 363922 466494 363978
rect 466562 363922 466618 363978
rect 466686 363922 466742 363978
rect 466314 346294 466370 346350
rect 466438 346294 466494 346350
rect 466562 346294 466618 346350
rect 466686 346294 466742 346350
rect 466314 346170 466370 346226
rect 466438 346170 466494 346226
rect 466562 346170 466618 346226
rect 466686 346170 466742 346226
rect 466314 346046 466370 346102
rect 466438 346046 466494 346102
rect 466562 346046 466618 346102
rect 466686 346046 466742 346102
rect 466314 345922 466370 345978
rect 466438 345922 466494 345978
rect 466562 345922 466618 345978
rect 466686 345922 466742 345978
rect 466314 328294 466370 328350
rect 466438 328294 466494 328350
rect 466562 328294 466618 328350
rect 466686 328294 466742 328350
rect 466314 328170 466370 328226
rect 466438 328170 466494 328226
rect 466562 328170 466618 328226
rect 466686 328170 466742 328226
rect 466314 328046 466370 328102
rect 466438 328046 466494 328102
rect 466562 328046 466618 328102
rect 466686 328046 466742 328102
rect 466314 327922 466370 327978
rect 466438 327922 466494 327978
rect 466562 327922 466618 327978
rect 466686 327922 466742 327978
rect 466314 310294 466370 310350
rect 466438 310294 466494 310350
rect 466562 310294 466618 310350
rect 466686 310294 466742 310350
rect 466314 310170 466370 310226
rect 466438 310170 466494 310226
rect 466562 310170 466618 310226
rect 466686 310170 466742 310226
rect 466314 310046 466370 310102
rect 466438 310046 466494 310102
rect 466562 310046 466618 310102
rect 466686 310046 466742 310102
rect 466314 309922 466370 309978
rect 466438 309922 466494 309978
rect 466562 309922 466618 309978
rect 466686 309922 466742 309978
rect 466314 292294 466370 292350
rect 466438 292294 466494 292350
rect 466562 292294 466618 292350
rect 466686 292294 466742 292350
rect 466314 292170 466370 292226
rect 466438 292170 466494 292226
rect 466562 292170 466618 292226
rect 466686 292170 466742 292226
rect 466314 292046 466370 292102
rect 466438 292046 466494 292102
rect 466562 292046 466618 292102
rect 466686 292046 466742 292102
rect 466314 291922 466370 291978
rect 466438 291922 466494 291978
rect 466562 291922 466618 291978
rect 466686 291922 466742 291978
rect 466314 274294 466370 274350
rect 466438 274294 466494 274350
rect 466562 274294 466618 274350
rect 466686 274294 466742 274350
rect 466314 274170 466370 274226
rect 466438 274170 466494 274226
rect 466562 274170 466618 274226
rect 466686 274170 466742 274226
rect 466314 274046 466370 274102
rect 466438 274046 466494 274102
rect 466562 274046 466618 274102
rect 466686 274046 466742 274102
rect 466314 273922 466370 273978
rect 466438 273922 466494 273978
rect 466562 273922 466618 273978
rect 466686 273922 466742 273978
rect 466314 256294 466370 256350
rect 466438 256294 466494 256350
rect 466562 256294 466618 256350
rect 466686 256294 466742 256350
rect 466314 256170 466370 256226
rect 466438 256170 466494 256226
rect 466562 256170 466618 256226
rect 466686 256170 466742 256226
rect 466314 256046 466370 256102
rect 466438 256046 466494 256102
rect 466562 256046 466618 256102
rect 466686 256046 466742 256102
rect 466314 255922 466370 255978
rect 466438 255922 466494 255978
rect 466562 255922 466618 255978
rect 466686 255922 466742 255978
rect 466314 238294 466370 238350
rect 466438 238294 466494 238350
rect 466562 238294 466618 238350
rect 466686 238294 466742 238350
rect 466314 238170 466370 238226
rect 466438 238170 466494 238226
rect 466562 238170 466618 238226
rect 466686 238170 466742 238226
rect 466314 238046 466370 238102
rect 466438 238046 466494 238102
rect 466562 238046 466618 238102
rect 466686 238046 466742 238102
rect 466314 237922 466370 237978
rect 466438 237922 466494 237978
rect 466562 237922 466618 237978
rect 466686 237922 466742 237978
rect 466314 220294 466370 220350
rect 466438 220294 466494 220350
rect 466562 220294 466618 220350
rect 466686 220294 466742 220350
rect 466314 220170 466370 220226
rect 466438 220170 466494 220226
rect 466562 220170 466618 220226
rect 466686 220170 466742 220226
rect 466314 220046 466370 220102
rect 466438 220046 466494 220102
rect 466562 220046 466618 220102
rect 466686 220046 466742 220102
rect 466314 219922 466370 219978
rect 466438 219922 466494 219978
rect 466562 219922 466618 219978
rect 466686 219922 466742 219978
rect 466314 202294 466370 202350
rect 466438 202294 466494 202350
rect 466562 202294 466618 202350
rect 466686 202294 466742 202350
rect 466314 202170 466370 202226
rect 466438 202170 466494 202226
rect 466562 202170 466618 202226
rect 466686 202170 466742 202226
rect 466314 202046 466370 202102
rect 466438 202046 466494 202102
rect 466562 202046 466618 202102
rect 466686 202046 466742 202102
rect 466314 201922 466370 201978
rect 466438 201922 466494 201978
rect 466562 201922 466618 201978
rect 466686 201922 466742 201978
rect 466314 184294 466370 184350
rect 466438 184294 466494 184350
rect 466562 184294 466618 184350
rect 466686 184294 466742 184350
rect 466314 184170 466370 184226
rect 466438 184170 466494 184226
rect 466562 184170 466618 184226
rect 466686 184170 466742 184226
rect 466314 184046 466370 184102
rect 466438 184046 466494 184102
rect 466562 184046 466618 184102
rect 466686 184046 466742 184102
rect 466314 183922 466370 183978
rect 466438 183922 466494 183978
rect 466562 183922 466618 183978
rect 466686 183922 466742 183978
rect 466314 166294 466370 166350
rect 466438 166294 466494 166350
rect 466562 166294 466618 166350
rect 466686 166294 466742 166350
rect 466314 166170 466370 166226
rect 466438 166170 466494 166226
rect 466562 166170 466618 166226
rect 466686 166170 466742 166226
rect 466314 166046 466370 166102
rect 466438 166046 466494 166102
rect 466562 166046 466618 166102
rect 466686 166046 466742 166102
rect 466314 165922 466370 165978
rect 466438 165922 466494 165978
rect 466562 165922 466618 165978
rect 466686 165922 466742 165978
rect 477148 407582 477204 407638
rect 475468 407402 475524 407458
rect 470034 406294 470090 406350
rect 470158 406294 470214 406350
rect 470282 406294 470338 406350
rect 470406 406294 470462 406350
rect 470034 406170 470090 406226
rect 470158 406170 470214 406226
rect 470282 406170 470338 406226
rect 470406 406170 470462 406226
rect 470034 406046 470090 406102
rect 470158 406046 470214 406102
rect 470282 406046 470338 406102
rect 470406 406046 470462 406102
rect 470034 405922 470090 405978
rect 470158 405922 470214 405978
rect 470282 405922 470338 405978
rect 470406 405922 470462 405978
rect 470034 388294 470090 388350
rect 470158 388294 470214 388350
rect 470282 388294 470338 388350
rect 470406 388294 470462 388350
rect 470034 388170 470090 388226
rect 470158 388170 470214 388226
rect 470282 388170 470338 388226
rect 470406 388170 470462 388226
rect 470034 388046 470090 388102
rect 470158 388046 470214 388102
rect 470282 388046 470338 388102
rect 470406 388046 470462 388102
rect 470034 387922 470090 387978
rect 470158 387922 470214 387978
rect 470282 387922 470338 387978
rect 470406 387922 470462 387978
rect 497034 400294 497090 400350
rect 497158 400294 497214 400350
rect 497282 400294 497338 400350
rect 497406 400294 497462 400350
rect 497034 400170 497090 400226
rect 497158 400170 497214 400226
rect 497282 400170 497338 400226
rect 497406 400170 497462 400226
rect 497034 400046 497090 400102
rect 497158 400046 497214 400102
rect 497282 400046 497338 400102
rect 497406 400046 497462 400102
rect 497034 399922 497090 399978
rect 497158 399922 497214 399978
rect 497282 399922 497338 399978
rect 497406 399922 497462 399978
rect 470034 370294 470090 370350
rect 470158 370294 470214 370350
rect 470282 370294 470338 370350
rect 470406 370294 470462 370350
rect 470034 370170 470090 370226
rect 470158 370170 470214 370226
rect 470282 370170 470338 370226
rect 470406 370170 470462 370226
rect 470034 370046 470090 370102
rect 470158 370046 470214 370102
rect 470282 370046 470338 370102
rect 470406 370046 470462 370102
rect 470034 369922 470090 369978
rect 470158 369922 470214 369978
rect 470282 369922 470338 369978
rect 470406 369922 470462 369978
rect 470034 352294 470090 352350
rect 470158 352294 470214 352350
rect 470282 352294 470338 352350
rect 470406 352294 470462 352350
rect 470034 352170 470090 352226
rect 470158 352170 470214 352226
rect 470282 352170 470338 352226
rect 470406 352170 470462 352226
rect 470034 352046 470090 352102
rect 470158 352046 470214 352102
rect 470282 352046 470338 352102
rect 470406 352046 470462 352102
rect 470034 351922 470090 351978
rect 470158 351922 470214 351978
rect 470282 351922 470338 351978
rect 470406 351922 470462 351978
rect 470034 334294 470090 334350
rect 470158 334294 470214 334350
rect 470282 334294 470338 334350
rect 470406 334294 470462 334350
rect 470034 334170 470090 334226
rect 470158 334170 470214 334226
rect 470282 334170 470338 334226
rect 470406 334170 470462 334226
rect 470034 334046 470090 334102
rect 470158 334046 470214 334102
rect 470282 334046 470338 334102
rect 470406 334046 470462 334102
rect 470034 333922 470090 333978
rect 470158 333922 470214 333978
rect 470282 333922 470338 333978
rect 470406 333922 470462 333978
rect 470034 316294 470090 316350
rect 470158 316294 470214 316350
rect 470282 316294 470338 316350
rect 470406 316294 470462 316350
rect 470034 316170 470090 316226
rect 470158 316170 470214 316226
rect 470282 316170 470338 316226
rect 470406 316170 470462 316226
rect 470034 316046 470090 316102
rect 470158 316046 470214 316102
rect 470282 316046 470338 316102
rect 470406 316046 470462 316102
rect 470034 315922 470090 315978
rect 470158 315922 470214 315978
rect 470282 315922 470338 315978
rect 470406 315922 470462 315978
rect 470034 298294 470090 298350
rect 470158 298294 470214 298350
rect 470282 298294 470338 298350
rect 470406 298294 470462 298350
rect 470034 298170 470090 298226
rect 470158 298170 470214 298226
rect 470282 298170 470338 298226
rect 470406 298170 470462 298226
rect 470034 298046 470090 298102
rect 470158 298046 470214 298102
rect 470282 298046 470338 298102
rect 470406 298046 470462 298102
rect 470034 297922 470090 297978
rect 470158 297922 470214 297978
rect 470282 297922 470338 297978
rect 470406 297922 470462 297978
rect 470034 280294 470090 280350
rect 470158 280294 470214 280350
rect 470282 280294 470338 280350
rect 470406 280294 470462 280350
rect 470034 280170 470090 280226
rect 470158 280170 470214 280226
rect 470282 280170 470338 280226
rect 470406 280170 470462 280226
rect 470034 280046 470090 280102
rect 470158 280046 470214 280102
rect 470282 280046 470338 280102
rect 470406 280046 470462 280102
rect 470034 279922 470090 279978
rect 470158 279922 470214 279978
rect 470282 279922 470338 279978
rect 470406 279922 470462 279978
rect 470034 262294 470090 262350
rect 470158 262294 470214 262350
rect 470282 262294 470338 262350
rect 470406 262294 470462 262350
rect 470034 262170 470090 262226
rect 470158 262170 470214 262226
rect 470282 262170 470338 262226
rect 470406 262170 470462 262226
rect 470034 262046 470090 262102
rect 470158 262046 470214 262102
rect 470282 262046 470338 262102
rect 470406 262046 470462 262102
rect 470034 261922 470090 261978
rect 470158 261922 470214 261978
rect 470282 261922 470338 261978
rect 470406 261922 470462 261978
rect 470034 244294 470090 244350
rect 470158 244294 470214 244350
rect 470282 244294 470338 244350
rect 470406 244294 470462 244350
rect 470034 244170 470090 244226
rect 470158 244170 470214 244226
rect 470282 244170 470338 244226
rect 470406 244170 470462 244226
rect 470034 244046 470090 244102
rect 470158 244046 470214 244102
rect 470282 244046 470338 244102
rect 470406 244046 470462 244102
rect 470034 243922 470090 243978
rect 470158 243922 470214 243978
rect 470282 243922 470338 243978
rect 470406 243922 470462 243978
rect 470034 226294 470090 226350
rect 470158 226294 470214 226350
rect 470282 226294 470338 226350
rect 470406 226294 470462 226350
rect 470034 226170 470090 226226
rect 470158 226170 470214 226226
rect 470282 226170 470338 226226
rect 470406 226170 470462 226226
rect 470034 226046 470090 226102
rect 470158 226046 470214 226102
rect 470282 226046 470338 226102
rect 470406 226046 470462 226102
rect 470034 225922 470090 225978
rect 470158 225922 470214 225978
rect 470282 225922 470338 225978
rect 470406 225922 470462 225978
rect 470034 208294 470090 208350
rect 470158 208294 470214 208350
rect 470282 208294 470338 208350
rect 470406 208294 470462 208350
rect 470034 208170 470090 208226
rect 470158 208170 470214 208226
rect 470282 208170 470338 208226
rect 470406 208170 470462 208226
rect 470034 208046 470090 208102
rect 470158 208046 470214 208102
rect 470282 208046 470338 208102
rect 470406 208046 470462 208102
rect 470034 207922 470090 207978
rect 470158 207922 470214 207978
rect 470282 207922 470338 207978
rect 470406 207922 470462 207978
rect 476252 384182 476308 384238
rect 476252 197882 476308 197938
rect 479612 384002 479668 384058
rect 481292 383822 481348 383878
rect 497034 382294 497090 382350
rect 497158 382294 497214 382350
rect 497282 382294 497338 382350
rect 497406 382294 497462 382350
rect 497034 382170 497090 382226
rect 497158 382170 497214 382226
rect 497282 382170 497338 382226
rect 497406 382170 497462 382226
rect 497034 382046 497090 382102
rect 497158 382046 497214 382102
rect 497282 382046 497338 382102
rect 497406 382046 497462 382102
rect 497034 381922 497090 381978
rect 497158 381922 497214 381978
rect 497282 381922 497338 381978
rect 497406 381922 497462 381978
rect 497034 364294 497090 364350
rect 497158 364294 497214 364350
rect 497282 364294 497338 364350
rect 497406 364294 497462 364350
rect 497034 364170 497090 364226
rect 497158 364170 497214 364226
rect 497282 364170 497338 364226
rect 497406 364170 497462 364226
rect 497034 364046 497090 364102
rect 497158 364046 497214 364102
rect 497282 364046 497338 364102
rect 497406 364046 497462 364102
rect 497034 363922 497090 363978
rect 497158 363922 497214 363978
rect 497282 363922 497338 363978
rect 497406 363922 497462 363978
rect 497034 346294 497090 346350
rect 497158 346294 497214 346350
rect 497282 346294 497338 346350
rect 497406 346294 497462 346350
rect 497034 346170 497090 346226
rect 497158 346170 497214 346226
rect 497282 346170 497338 346226
rect 497406 346170 497462 346226
rect 497034 346046 497090 346102
rect 497158 346046 497214 346102
rect 497282 346046 497338 346102
rect 497406 346046 497462 346102
rect 497034 345922 497090 345978
rect 497158 345922 497214 345978
rect 497282 345922 497338 345978
rect 497406 345922 497462 345978
rect 497034 328294 497090 328350
rect 497158 328294 497214 328350
rect 497282 328294 497338 328350
rect 497406 328294 497462 328350
rect 497034 328170 497090 328226
rect 497158 328170 497214 328226
rect 497282 328170 497338 328226
rect 497406 328170 497462 328226
rect 497034 328046 497090 328102
rect 497158 328046 497214 328102
rect 497282 328046 497338 328102
rect 497406 328046 497462 328102
rect 497034 327922 497090 327978
rect 497158 327922 497214 327978
rect 497282 327922 497338 327978
rect 497406 327922 497462 327978
rect 497034 310294 497090 310350
rect 497158 310294 497214 310350
rect 497282 310294 497338 310350
rect 497406 310294 497462 310350
rect 497034 310170 497090 310226
rect 497158 310170 497214 310226
rect 497282 310170 497338 310226
rect 497406 310170 497462 310226
rect 497034 310046 497090 310102
rect 497158 310046 497214 310102
rect 497282 310046 497338 310102
rect 497406 310046 497462 310102
rect 497034 309922 497090 309978
rect 497158 309922 497214 309978
rect 497282 309922 497338 309978
rect 497406 309922 497462 309978
rect 497034 292294 497090 292350
rect 497158 292294 497214 292350
rect 497282 292294 497338 292350
rect 497406 292294 497462 292350
rect 497034 292170 497090 292226
rect 497158 292170 497214 292226
rect 497282 292170 497338 292226
rect 497406 292170 497462 292226
rect 497034 292046 497090 292102
rect 497158 292046 497214 292102
rect 497282 292046 497338 292102
rect 497406 292046 497462 292102
rect 497034 291922 497090 291978
rect 497158 291922 497214 291978
rect 497282 291922 497338 291978
rect 497406 291922 497462 291978
rect 497034 274294 497090 274350
rect 497158 274294 497214 274350
rect 497282 274294 497338 274350
rect 497406 274294 497462 274350
rect 497034 274170 497090 274226
rect 497158 274170 497214 274226
rect 497282 274170 497338 274226
rect 497406 274170 497462 274226
rect 497034 274046 497090 274102
rect 497158 274046 497214 274102
rect 497282 274046 497338 274102
rect 497406 274046 497462 274102
rect 497034 273922 497090 273978
rect 497158 273922 497214 273978
rect 497282 273922 497338 273978
rect 497406 273922 497462 273978
rect 497034 256294 497090 256350
rect 497158 256294 497214 256350
rect 497282 256294 497338 256350
rect 497406 256294 497462 256350
rect 497034 256170 497090 256226
rect 497158 256170 497214 256226
rect 497282 256170 497338 256226
rect 497406 256170 497462 256226
rect 497034 256046 497090 256102
rect 497158 256046 497214 256102
rect 497282 256046 497338 256102
rect 497406 256046 497462 256102
rect 497034 255922 497090 255978
rect 497158 255922 497214 255978
rect 497282 255922 497338 255978
rect 497406 255922 497462 255978
rect 497034 238294 497090 238350
rect 497158 238294 497214 238350
rect 497282 238294 497338 238350
rect 497406 238294 497462 238350
rect 497034 238170 497090 238226
rect 497158 238170 497214 238226
rect 497282 238170 497338 238226
rect 497406 238170 497462 238226
rect 497034 238046 497090 238102
rect 497158 238046 497214 238102
rect 497282 238046 497338 238102
rect 497406 238046 497462 238102
rect 497034 237922 497090 237978
rect 497158 237922 497214 237978
rect 497282 237922 497338 237978
rect 497406 237922 497462 237978
rect 500754 406294 500810 406350
rect 500878 406294 500934 406350
rect 501002 406294 501058 406350
rect 501126 406294 501182 406350
rect 500754 406170 500810 406226
rect 500878 406170 500934 406226
rect 501002 406170 501058 406226
rect 501126 406170 501182 406226
rect 500754 406046 500810 406102
rect 500878 406046 500934 406102
rect 501002 406046 501058 406102
rect 501126 406046 501182 406102
rect 500754 405922 500810 405978
rect 500878 405922 500934 405978
rect 501002 405922 501058 405978
rect 501126 405922 501182 405978
rect 500754 388294 500810 388350
rect 500878 388294 500934 388350
rect 501002 388294 501058 388350
rect 501126 388294 501182 388350
rect 500754 388170 500810 388226
rect 500878 388170 500934 388226
rect 501002 388170 501058 388226
rect 501126 388170 501182 388226
rect 500754 388046 500810 388102
rect 500878 388046 500934 388102
rect 501002 388046 501058 388102
rect 501126 388046 501182 388102
rect 500754 387922 500810 387978
rect 500878 387922 500934 387978
rect 501002 387922 501058 387978
rect 501126 387922 501182 387978
rect 527754 400294 527810 400350
rect 527878 400294 527934 400350
rect 528002 400294 528058 400350
rect 528126 400294 528182 400350
rect 527754 400170 527810 400226
rect 527878 400170 527934 400226
rect 528002 400170 528058 400226
rect 528126 400170 528182 400226
rect 527754 400046 527810 400102
rect 527878 400046 527934 400102
rect 528002 400046 528058 400102
rect 528126 400046 528182 400102
rect 527754 399922 527810 399978
rect 527878 399922 527934 399978
rect 528002 399922 528058 399978
rect 528126 399922 528182 399978
rect 500754 370294 500810 370350
rect 500878 370294 500934 370350
rect 501002 370294 501058 370350
rect 501126 370294 501182 370350
rect 500754 370170 500810 370226
rect 500878 370170 500934 370226
rect 501002 370170 501058 370226
rect 501126 370170 501182 370226
rect 500754 370046 500810 370102
rect 500878 370046 500934 370102
rect 501002 370046 501058 370102
rect 501126 370046 501182 370102
rect 500754 369922 500810 369978
rect 500878 369922 500934 369978
rect 501002 369922 501058 369978
rect 501126 369922 501182 369978
rect 500754 352294 500810 352350
rect 500878 352294 500934 352350
rect 501002 352294 501058 352350
rect 501126 352294 501182 352350
rect 500754 352170 500810 352226
rect 500878 352170 500934 352226
rect 501002 352170 501058 352226
rect 501126 352170 501182 352226
rect 500754 352046 500810 352102
rect 500878 352046 500934 352102
rect 501002 352046 501058 352102
rect 501126 352046 501182 352102
rect 500754 351922 500810 351978
rect 500878 351922 500934 351978
rect 501002 351922 501058 351978
rect 501126 351922 501182 351978
rect 519932 382562 519988 382618
rect 527754 382294 527810 382350
rect 527878 382294 527934 382350
rect 528002 382294 528058 382350
rect 528126 382294 528182 382350
rect 527754 382170 527810 382226
rect 527878 382170 527934 382226
rect 528002 382170 528058 382226
rect 528126 382170 528182 382226
rect 527754 382046 527810 382102
rect 527878 382046 527934 382102
rect 528002 382046 528058 382102
rect 528126 382046 528182 382102
rect 527754 381922 527810 381978
rect 527878 381922 527934 381978
rect 528002 381922 528058 381978
rect 528126 381922 528182 381978
rect 527754 364294 527810 364350
rect 527878 364294 527934 364350
rect 528002 364294 528058 364350
rect 528126 364294 528182 364350
rect 527754 364170 527810 364226
rect 527878 364170 527934 364226
rect 528002 364170 528058 364226
rect 528126 364170 528182 364226
rect 527754 364046 527810 364102
rect 527878 364046 527934 364102
rect 528002 364046 528058 364102
rect 528126 364046 528182 364102
rect 527754 363922 527810 363978
rect 527878 363922 527934 363978
rect 528002 363922 528058 363978
rect 528126 363922 528182 363978
rect 500754 334294 500810 334350
rect 500878 334294 500934 334350
rect 501002 334294 501058 334350
rect 501126 334294 501182 334350
rect 500754 334170 500810 334226
rect 500878 334170 500934 334226
rect 501002 334170 501058 334226
rect 501126 334170 501182 334226
rect 500754 334046 500810 334102
rect 500878 334046 500934 334102
rect 501002 334046 501058 334102
rect 501126 334046 501182 334102
rect 500754 333922 500810 333978
rect 500878 333922 500934 333978
rect 501002 333922 501058 333978
rect 501126 333922 501182 333978
rect 527754 346294 527810 346350
rect 527878 346294 527934 346350
rect 528002 346294 528058 346350
rect 528126 346294 528182 346350
rect 527754 346170 527810 346226
rect 527878 346170 527934 346226
rect 528002 346170 528058 346226
rect 528126 346170 528182 346226
rect 527754 346046 527810 346102
rect 527878 346046 527934 346102
rect 528002 346046 528058 346102
rect 528126 346046 528182 346102
rect 527754 345922 527810 345978
rect 527878 345922 527934 345978
rect 528002 345922 528058 345978
rect 528126 345922 528182 345978
rect 527754 328294 527810 328350
rect 527878 328294 527934 328350
rect 528002 328294 528058 328350
rect 528126 328294 528182 328350
rect 527754 328170 527810 328226
rect 527878 328170 527934 328226
rect 528002 328170 528058 328226
rect 528126 328170 528182 328226
rect 527754 328046 527810 328102
rect 527878 328046 527934 328102
rect 528002 328046 528058 328102
rect 528126 328046 528182 328102
rect 527754 327922 527810 327978
rect 527878 327922 527934 327978
rect 528002 327922 528058 327978
rect 528126 327922 528182 327978
rect 500754 316294 500810 316350
rect 500878 316294 500934 316350
rect 501002 316294 501058 316350
rect 501126 316294 501182 316350
rect 500754 316170 500810 316226
rect 500878 316170 500934 316226
rect 501002 316170 501058 316226
rect 501126 316170 501182 316226
rect 500754 316046 500810 316102
rect 500878 316046 500934 316102
rect 501002 316046 501058 316102
rect 501126 316046 501182 316102
rect 500754 315922 500810 315978
rect 500878 315922 500934 315978
rect 501002 315922 501058 315978
rect 501126 315922 501182 315978
rect 500754 298294 500810 298350
rect 500878 298294 500934 298350
rect 501002 298294 501058 298350
rect 501126 298294 501182 298350
rect 500754 298170 500810 298226
rect 500878 298170 500934 298226
rect 501002 298170 501058 298226
rect 501126 298170 501182 298226
rect 500754 298046 500810 298102
rect 500878 298046 500934 298102
rect 501002 298046 501058 298102
rect 501126 298046 501182 298102
rect 500754 297922 500810 297978
rect 500878 297922 500934 297978
rect 501002 297922 501058 297978
rect 501126 297922 501182 297978
rect 500754 280294 500810 280350
rect 500878 280294 500934 280350
rect 501002 280294 501058 280350
rect 501126 280294 501182 280350
rect 500754 280170 500810 280226
rect 500878 280170 500934 280226
rect 501002 280170 501058 280226
rect 501126 280170 501182 280226
rect 500754 280046 500810 280102
rect 500878 280046 500934 280102
rect 501002 280046 501058 280102
rect 501126 280046 501182 280102
rect 500754 279922 500810 279978
rect 500878 279922 500934 279978
rect 501002 279922 501058 279978
rect 501126 279922 501182 279978
rect 500754 262294 500810 262350
rect 500878 262294 500934 262350
rect 501002 262294 501058 262350
rect 501126 262294 501182 262350
rect 500754 262170 500810 262226
rect 500878 262170 500934 262226
rect 501002 262170 501058 262226
rect 501126 262170 501182 262226
rect 500754 262046 500810 262102
rect 500878 262046 500934 262102
rect 501002 262046 501058 262102
rect 501126 262046 501182 262102
rect 500754 261922 500810 261978
rect 500878 261922 500934 261978
rect 501002 261922 501058 261978
rect 501126 261922 501182 261978
rect 500754 244294 500810 244350
rect 500878 244294 500934 244350
rect 501002 244294 501058 244350
rect 501126 244294 501182 244350
rect 500754 244170 500810 244226
rect 500878 244170 500934 244226
rect 501002 244170 501058 244226
rect 501126 244170 501182 244226
rect 500754 244046 500810 244102
rect 500878 244046 500934 244102
rect 501002 244046 501058 244102
rect 501126 244046 501182 244102
rect 500754 243922 500810 243978
rect 500878 243922 500934 243978
rect 501002 243922 501058 243978
rect 501126 243922 501182 243978
rect 527754 310294 527810 310350
rect 527878 310294 527934 310350
rect 528002 310294 528058 310350
rect 528126 310294 528182 310350
rect 527754 310170 527810 310226
rect 527878 310170 527934 310226
rect 528002 310170 528058 310226
rect 528126 310170 528182 310226
rect 527754 310046 527810 310102
rect 527878 310046 527934 310102
rect 528002 310046 528058 310102
rect 528126 310046 528182 310102
rect 527754 309922 527810 309978
rect 527878 309922 527934 309978
rect 528002 309922 528058 309978
rect 528126 309922 528182 309978
rect 527754 292294 527810 292350
rect 527878 292294 527934 292350
rect 528002 292294 528058 292350
rect 528126 292294 528182 292350
rect 527754 292170 527810 292226
rect 527878 292170 527934 292226
rect 528002 292170 528058 292226
rect 528126 292170 528182 292226
rect 527754 292046 527810 292102
rect 527878 292046 527934 292102
rect 528002 292046 528058 292102
rect 528126 292046 528182 292102
rect 527754 291922 527810 291978
rect 527878 291922 527934 291978
rect 528002 291922 528058 291978
rect 528126 291922 528182 291978
rect 527754 274294 527810 274350
rect 527878 274294 527934 274350
rect 528002 274294 528058 274350
rect 528126 274294 528182 274350
rect 527754 274170 527810 274226
rect 527878 274170 527934 274226
rect 528002 274170 528058 274226
rect 528126 274170 528182 274226
rect 527754 274046 527810 274102
rect 527878 274046 527934 274102
rect 528002 274046 528058 274102
rect 528126 274046 528182 274102
rect 527754 273922 527810 273978
rect 527878 273922 527934 273978
rect 528002 273922 528058 273978
rect 528126 273922 528182 273978
rect 527754 256294 527810 256350
rect 527878 256294 527934 256350
rect 528002 256294 528058 256350
rect 528126 256294 528182 256350
rect 527754 256170 527810 256226
rect 527878 256170 527934 256226
rect 528002 256170 528058 256226
rect 528126 256170 528182 256226
rect 527754 256046 527810 256102
rect 527878 256046 527934 256102
rect 528002 256046 528058 256102
rect 528126 256046 528182 256102
rect 527754 255922 527810 255978
rect 527878 255922 527934 255978
rect 528002 255922 528058 255978
rect 528126 255922 528182 255978
rect 527754 238294 527810 238350
rect 527878 238294 527934 238350
rect 528002 238294 528058 238350
rect 528126 238294 528182 238350
rect 527754 238170 527810 238226
rect 527878 238170 527934 238226
rect 528002 238170 528058 238226
rect 528126 238170 528182 238226
rect 527754 238046 527810 238102
rect 527878 238046 527934 238102
rect 528002 238046 528058 238102
rect 528126 238046 528182 238102
rect 527754 237922 527810 237978
rect 527878 237922 527934 237978
rect 528002 237922 528058 237978
rect 528126 237922 528182 237978
rect 489822 226294 489878 226350
rect 489946 226294 490002 226350
rect 489822 226170 489878 226226
rect 489946 226170 490002 226226
rect 489822 226046 489878 226102
rect 489946 226046 490002 226102
rect 489822 225922 489878 225978
rect 489946 225922 490002 225978
rect 498390 226294 498446 226350
rect 498514 226294 498570 226350
rect 498390 226170 498446 226226
rect 498514 226170 498570 226226
rect 498390 226046 498446 226102
rect 498514 226046 498570 226102
rect 498390 225922 498446 225978
rect 498514 225922 498570 225978
rect 506958 226294 507014 226350
rect 507082 226294 507138 226350
rect 506958 226170 507014 226226
rect 507082 226170 507138 226226
rect 506958 226046 507014 226102
rect 507082 226046 507138 226102
rect 506958 225922 507014 225978
rect 507082 225922 507138 225978
rect 515526 226294 515582 226350
rect 515650 226294 515706 226350
rect 515526 226170 515582 226226
rect 515650 226170 515706 226226
rect 515526 226046 515582 226102
rect 515650 226046 515706 226102
rect 515526 225922 515582 225978
rect 515650 225922 515706 225978
rect 485538 220294 485594 220350
rect 485662 220294 485718 220350
rect 485538 220170 485594 220226
rect 485662 220170 485718 220226
rect 485538 220046 485594 220102
rect 485662 220046 485718 220102
rect 485538 219922 485594 219978
rect 485662 219922 485718 219978
rect 494106 220294 494162 220350
rect 494230 220294 494286 220350
rect 494106 220170 494162 220226
rect 494230 220170 494286 220226
rect 494106 220046 494162 220102
rect 494230 220046 494286 220102
rect 494106 219922 494162 219978
rect 494230 219922 494286 219978
rect 502674 220294 502730 220350
rect 502798 220294 502854 220350
rect 502674 220170 502730 220226
rect 502798 220170 502854 220226
rect 502674 220046 502730 220102
rect 502798 220046 502854 220102
rect 502674 219922 502730 219978
rect 502798 219922 502854 219978
rect 511242 220294 511298 220350
rect 511366 220294 511422 220350
rect 511242 220170 511298 220226
rect 511366 220170 511422 220226
rect 511242 220046 511298 220102
rect 511366 220046 511422 220102
rect 511242 219922 511298 219978
rect 511366 219922 511422 219978
rect 489822 208294 489878 208350
rect 489946 208294 490002 208350
rect 489822 208170 489878 208226
rect 489946 208170 490002 208226
rect 489822 208046 489878 208102
rect 489946 208046 490002 208102
rect 489822 207922 489878 207978
rect 489946 207922 490002 207978
rect 498390 208294 498446 208350
rect 498514 208294 498570 208350
rect 498390 208170 498446 208226
rect 498514 208170 498570 208226
rect 498390 208046 498446 208102
rect 498514 208046 498570 208102
rect 498390 207922 498446 207978
rect 498514 207922 498570 207978
rect 506958 208294 507014 208350
rect 507082 208294 507138 208350
rect 506958 208170 507014 208226
rect 507082 208170 507138 208226
rect 506958 208046 507014 208102
rect 507082 208046 507138 208102
rect 506958 207922 507014 207978
rect 507082 207922 507138 207978
rect 515526 208294 515582 208350
rect 515650 208294 515706 208350
rect 515526 208170 515582 208226
rect 515650 208170 515706 208226
rect 515526 208046 515582 208102
rect 515650 208046 515706 208102
rect 515526 207922 515582 207978
rect 515650 207922 515706 207978
rect 527754 220294 527810 220350
rect 527878 220294 527934 220350
rect 528002 220294 528058 220350
rect 528126 220294 528182 220350
rect 527754 220170 527810 220226
rect 527878 220170 527934 220226
rect 528002 220170 528058 220226
rect 528126 220170 528182 220226
rect 527754 220046 527810 220102
rect 527878 220046 527934 220102
rect 528002 220046 528058 220102
rect 528126 220046 528182 220102
rect 527754 219922 527810 219978
rect 527878 219922 527934 219978
rect 528002 219922 528058 219978
rect 528126 219922 528182 219978
rect 497034 202294 497090 202350
rect 497158 202294 497214 202350
rect 497282 202294 497338 202350
rect 497406 202294 497462 202350
rect 497034 202170 497090 202226
rect 497158 202170 497214 202226
rect 497282 202170 497338 202226
rect 497406 202170 497462 202226
rect 497034 202046 497090 202102
rect 497158 202046 497214 202102
rect 497282 202046 497338 202102
rect 497406 202046 497462 202102
rect 497034 201922 497090 201978
rect 497158 201922 497214 201978
rect 497282 201922 497338 201978
rect 497406 201922 497462 201978
rect 479612 197702 479668 197758
rect 470034 190294 470090 190350
rect 470158 190294 470214 190350
rect 470282 190294 470338 190350
rect 470406 190294 470462 190350
rect 470034 190170 470090 190226
rect 470158 190170 470214 190226
rect 470282 190170 470338 190226
rect 470406 190170 470462 190226
rect 470034 190046 470090 190102
rect 470158 190046 470214 190102
rect 470282 190046 470338 190102
rect 470406 190046 470462 190102
rect 470034 189922 470090 189978
rect 470158 189922 470214 189978
rect 470282 189922 470338 189978
rect 470406 189922 470462 189978
rect 470034 172294 470090 172350
rect 470158 172294 470214 172350
rect 470282 172294 470338 172350
rect 470406 172294 470462 172350
rect 470034 172170 470090 172226
rect 470158 172170 470214 172226
rect 470282 172170 470338 172226
rect 470406 172170 470462 172226
rect 470034 172046 470090 172102
rect 470158 172046 470214 172102
rect 470282 172046 470338 172102
rect 470406 172046 470462 172102
rect 470034 171922 470090 171978
rect 470158 171922 470214 171978
rect 470282 171922 470338 171978
rect 470406 171922 470462 171978
rect 470034 154294 470090 154350
rect 470158 154294 470214 154350
rect 470282 154294 470338 154350
rect 470406 154294 470462 154350
rect 470034 154170 470090 154226
rect 470158 154170 470214 154226
rect 470282 154170 470338 154226
rect 470406 154170 470462 154226
rect 470034 154046 470090 154102
rect 470158 154046 470214 154102
rect 470282 154046 470338 154102
rect 470406 154046 470462 154102
rect 470034 153922 470090 153978
rect 470158 153922 470214 153978
rect 470282 153922 470338 153978
rect 470406 153922 470462 153978
rect 497644 198062 497700 198118
rect 499100 197882 499156 197938
rect 497034 184294 497090 184350
rect 497158 184294 497214 184350
rect 497282 184294 497338 184350
rect 497406 184294 497462 184350
rect 497034 184170 497090 184226
rect 497158 184170 497214 184226
rect 497282 184170 497338 184226
rect 497406 184170 497462 184226
rect 497034 184046 497090 184102
rect 497158 184046 497214 184102
rect 497282 184046 497338 184102
rect 497406 184046 497462 184102
rect 497034 183922 497090 183978
rect 497158 183922 497214 183978
rect 497282 183922 497338 183978
rect 497406 183922 497462 183978
rect 497034 166294 497090 166350
rect 497158 166294 497214 166350
rect 497282 166294 497338 166350
rect 497406 166294 497462 166350
rect 497034 166170 497090 166226
rect 497158 166170 497214 166226
rect 497282 166170 497338 166226
rect 497406 166170 497462 166226
rect 497034 166046 497090 166102
rect 497158 166046 497214 166102
rect 497282 166046 497338 166102
rect 497406 166046 497462 166102
rect 497034 165922 497090 165978
rect 497158 165922 497214 165978
rect 497282 165922 497338 165978
rect 497406 165922 497462 165978
rect 495852 153602 495908 153658
rect 527754 202294 527810 202350
rect 527878 202294 527934 202350
rect 528002 202294 528058 202350
rect 528126 202294 528182 202350
rect 527754 202170 527810 202226
rect 527878 202170 527934 202226
rect 528002 202170 528058 202226
rect 528126 202170 528182 202226
rect 527754 202046 527810 202102
rect 527878 202046 527934 202102
rect 528002 202046 528058 202102
rect 528126 202046 528182 202102
rect 527754 201922 527810 201978
rect 527878 201922 527934 201978
rect 528002 201922 528058 201978
rect 528126 201922 528182 201978
rect 502236 197702 502292 197758
rect 500754 190294 500810 190350
rect 500878 190294 500934 190350
rect 501002 190294 501058 190350
rect 501126 190294 501182 190350
rect 500754 190170 500810 190226
rect 500878 190170 500934 190226
rect 501002 190170 501058 190226
rect 501126 190170 501182 190226
rect 500754 190046 500810 190102
rect 500878 190046 500934 190102
rect 501002 190046 501058 190102
rect 501126 190046 501182 190102
rect 500754 189922 500810 189978
rect 500878 189922 500934 189978
rect 501002 189922 501058 189978
rect 501126 189922 501182 189978
rect 500754 172294 500810 172350
rect 500878 172294 500934 172350
rect 501002 172294 501058 172350
rect 501126 172294 501182 172350
rect 500754 172170 500810 172226
rect 500878 172170 500934 172226
rect 501002 172170 501058 172226
rect 501126 172170 501182 172226
rect 500754 172046 500810 172102
rect 500878 172046 500934 172102
rect 501002 172046 501058 172102
rect 501126 172046 501182 172102
rect 500754 171922 500810 171978
rect 500878 171922 500934 171978
rect 501002 171922 501058 171978
rect 501126 171922 501182 171978
rect 500754 154294 500810 154350
rect 500878 154294 500934 154350
rect 501002 154294 501058 154350
rect 501126 154294 501182 154350
rect 500754 154170 500810 154226
rect 500878 154170 500934 154226
rect 501002 154170 501058 154226
rect 501126 154170 501182 154226
rect 500754 154046 500810 154102
rect 500878 154046 500934 154102
rect 501002 154046 501058 154102
rect 501126 154046 501182 154102
rect 500754 153922 500810 153978
rect 500878 153922 500934 153978
rect 501002 153922 501058 153978
rect 501126 153922 501182 153978
rect 527754 184294 527810 184350
rect 527878 184294 527934 184350
rect 528002 184294 528058 184350
rect 528126 184294 528182 184350
rect 527754 184170 527810 184226
rect 527878 184170 527934 184226
rect 528002 184170 528058 184226
rect 528126 184170 528182 184226
rect 527754 184046 527810 184102
rect 527878 184046 527934 184102
rect 528002 184046 528058 184102
rect 528126 184046 528182 184102
rect 527754 183922 527810 183978
rect 527878 183922 527934 183978
rect 528002 183922 528058 183978
rect 528126 183922 528182 183978
rect 527754 166294 527810 166350
rect 527878 166294 527934 166350
rect 528002 166294 528058 166350
rect 528126 166294 528182 166350
rect 527754 166170 527810 166226
rect 527878 166170 527934 166226
rect 528002 166170 528058 166226
rect 528126 166170 528182 166226
rect 527754 166046 527810 166102
rect 527878 166046 527934 166102
rect 528002 166046 528058 166102
rect 528126 166046 528182 166102
rect 527754 165922 527810 165978
rect 527878 165922 527934 165978
rect 528002 165922 528058 165978
rect 528126 165922 528182 165978
rect 501340 152908 501396 152938
rect 501340 152882 501396 152908
rect 558474 580294 558530 580350
rect 558598 580294 558654 580350
rect 558722 580294 558778 580350
rect 558846 580294 558902 580350
rect 558474 580170 558530 580226
rect 558598 580170 558654 580226
rect 558722 580170 558778 580226
rect 558846 580170 558902 580226
rect 558474 580046 558530 580102
rect 558598 580046 558654 580102
rect 558722 580046 558778 580102
rect 558846 580046 558902 580102
rect 558474 579922 558530 579978
rect 558598 579922 558654 579978
rect 558722 579922 558778 579978
rect 558846 579922 558902 579978
rect 558474 562294 558530 562350
rect 558598 562294 558654 562350
rect 558722 562294 558778 562350
rect 558846 562294 558902 562350
rect 558474 562170 558530 562226
rect 558598 562170 558654 562226
rect 558722 562170 558778 562226
rect 558846 562170 558902 562226
rect 558474 562046 558530 562102
rect 558598 562046 558654 562102
rect 558722 562046 558778 562102
rect 558846 562046 558902 562102
rect 558474 561922 558530 561978
rect 558598 561922 558654 561978
rect 558722 561922 558778 561978
rect 558846 561922 558902 561978
rect 547798 550294 547854 550350
rect 547922 550294 547978 550350
rect 547798 550170 547854 550226
rect 547922 550170 547978 550226
rect 547798 550046 547854 550102
rect 547922 550046 547978 550102
rect 547798 549922 547854 549978
rect 547922 549922 547978 549978
rect 558474 544294 558530 544350
rect 558598 544294 558654 544350
rect 558722 544294 558778 544350
rect 558846 544294 558902 544350
rect 558474 544170 558530 544226
rect 558598 544170 558654 544226
rect 558722 544170 558778 544226
rect 558846 544170 558902 544226
rect 558474 544046 558530 544102
rect 558598 544046 558654 544102
rect 558722 544046 558778 544102
rect 558846 544046 558902 544102
rect 558474 543922 558530 543978
rect 558598 543922 558654 543978
rect 558722 543922 558778 543978
rect 558846 543922 558902 543978
rect 547798 532294 547854 532350
rect 547922 532294 547978 532350
rect 547798 532170 547854 532226
rect 547922 532170 547978 532226
rect 547798 532046 547854 532102
rect 547922 532046 547978 532102
rect 547798 531922 547854 531978
rect 547922 531922 547978 531978
rect 558474 526294 558530 526350
rect 558598 526294 558654 526350
rect 558722 526294 558778 526350
rect 558846 526294 558902 526350
rect 558474 526170 558530 526226
rect 558598 526170 558654 526226
rect 558722 526170 558778 526226
rect 558846 526170 558902 526226
rect 558474 526046 558530 526102
rect 558598 526046 558654 526102
rect 558722 526046 558778 526102
rect 558846 526046 558902 526102
rect 558474 525922 558530 525978
rect 558598 525922 558654 525978
rect 558722 525922 558778 525978
rect 558846 525922 558902 525978
rect 547798 514294 547854 514350
rect 547922 514294 547978 514350
rect 547798 514170 547854 514226
rect 547922 514170 547978 514226
rect 547798 514046 547854 514102
rect 547922 514046 547978 514102
rect 547798 513922 547854 513978
rect 547922 513922 547978 513978
rect 558474 508294 558530 508350
rect 558598 508294 558654 508350
rect 558722 508294 558778 508350
rect 558846 508294 558902 508350
rect 558474 508170 558530 508226
rect 558598 508170 558654 508226
rect 558722 508170 558778 508226
rect 558846 508170 558902 508226
rect 558474 508046 558530 508102
rect 558598 508046 558654 508102
rect 558722 508046 558778 508102
rect 558846 508046 558902 508102
rect 558474 507922 558530 507978
rect 558598 507922 558654 507978
rect 558722 507922 558778 507978
rect 558846 507922 558902 507978
rect 547798 496294 547854 496350
rect 547922 496294 547978 496350
rect 547798 496170 547854 496226
rect 547922 496170 547978 496226
rect 547798 496046 547854 496102
rect 547922 496046 547978 496102
rect 547798 495922 547854 495978
rect 547922 495922 547978 495978
rect 558474 490294 558530 490350
rect 558598 490294 558654 490350
rect 558722 490294 558778 490350
rect 558846 490294 558902 490350
rect 558474 490170 558530 490226
rect 558598 490170 558654 490226
rect 558722 490170 558778 490226
rect 558846 490170 558902 490226
rect 558474 490046 558530 490102
rect 558598 490046 558654 490102
rect 558722 490046 558778 490102
rect 558846 490046 558902 490102
rect 558474 489922 558530 489978
rect 558598 489922 558654 489978
rect 558722 489922 558778 489978
rect 558846 489922 558902 489978
rect 547798 478294 547854 478350
rect 547922 478294 547978 478350
rect 547798 478170 547854 478226
rect 547922 478170 547978 478226
rect 547798 478046 547854 478102
rect 547922 478046 547978 478102
rect 547798 477922 547854 477978
rect 547922 477922 547978 477978
rect 558474 472294 558530 472350
rect 558598 472294 558654 472350
rect 558722 472294 558778 472350
rect 558846 472294 558902 472350
rect 558474 472170 558530 472226
rect 558598 472170 558654 472226
rect 558722 472170 558778 472226
rect 558846 472170 558902 472226
rect 558474 472046 558530 472102
rect 558598 472046 558654 472102
rect 558722 472046 558778 472102
rect 558846 472046 558902 472102
rect 558474 471922 558530 471978
rect 558598 471922 558654 471978
rect 558722 471922 558778 471978
rect 558846 471922 558902 471978
rect 547798 460294 547854 460350
rect 547922 460294 547978 460350
rect 547798 460170 547854 460226
rect 547922 460170 547978 460226
rect 547798 460046 547854 460102
rect 547922 460046 547978 460102
rect 547798 459922 547854 459978
rect 547922 459922 547978 459978
rect 558474 454294 558530 454350
rect 558598 454294 558654 454350
rect 558722 454294 558778 454350
rect 558846 454294 558902 454350
rect 558474 454170 558530 454226
rect 558598 454170 558654 454226
rect 558722 454170 558778 454226
rect 558846 454170 558902 454226
rect 558474 454046 558530 454102
rect 558598 454046 558654 454102
rect 558722 454046 558778 454102
rect 558846 454046 558902 454102
rect 558474 453922 558530 453978
rect 558598 453922 558654 453978
rect 558722 453922 558778 453978
rect 558846 453922 558902 453978
rect 547798 442294 547854 442350
rect 547922 442294 547978 442350
rect 547798 442170 547854 442226
rect 547922 442170 547978 442226
rect 547798 442046 547854 442102
rect 547922 442046 547978 442102
rect 547798 441922 547854 441978
rect 547922 441922 547978 441978
rect 558474 436294 558530 436350
rect 558598 436294 558654 436350
rect 558722 436294 558778 436350
rect 558846 436294 558902 436350
rect 558474 436170 558530 436226
rect 558598 436170 558654 436226
rect 558722 436170 558778 436226
rect 558846 436170 558902 436226
rect 558474 436046 558530 436102
rect 558598 436046 558654 436102
rect 558722 436046 558778 436102
rect 558846 436046 558902 436102
rect 558474 435922 558530 435978
rect 558598 435922 558654 435978
rect 558722 435922 558778 435978
rect 558846 435922 558902 435978
rect 547798 424294 547854 424350
rect 547922 424294 547978 424350
rect 547798 424170 547854 424226
rect 547922 424170 547978 424226
rect 547798 424046 547854 424102
rect 547922 424046 547978 424102
rect 547798 423922 547854 423978
rect 547922 423922 547978 423978
rect 558474 418294 558530 418350
rect 558598 418294 558654 418350
rect 558722 418294 558778 418350
rect 558846 418294 558902 418350
rect 558474 418170 558530 418226
rect 558598 418170 558654 418226
rect 558722 418170 558778 418226
rect 558846 418170 558902 418226
rect 558474 418046 558530 418102
rect 558598 418046 558654 418102
rect 558722 418046 558778 418102
rect 558846 418046 558902 418102
rect 558474 417922 558530 417978
rect 558598 417922 558654 417978
rect 558722 417922 558778 417978
rect 558846 417922 558902 417978
rect 531474 406294 531530 406350
rect 531598 406294 531654 406350
rect 531722 406294 531778 406350
rect 531846 406294 531902 406350
rect 531474 406170 531530 406226
rect 531598 406170 531654 406226
rect 531722 406170 531778 406226
rect 531846 406170 531902 406226
rect 531474 406046 531530 406102
rect 531598 406046 531654 406102
rect 531722 406046 531778 406102
rect 531846 406046 531902 406102
rect 531474 405922 531530 405978
rect 531598 405922 531654 405978
rect 531722 405922 531778 405978
rect 531846 405922 531902 405978
rect 531474 388294 531530 388350
rect 531598 388294 531654 388350
rect 531722 388294 531778 388350
rect 531846 388294 531902 388350
rect 531474 388170 531530 388226
rect 531598 388170 531654 388226
rect 531722 388170 531778 388226
rect 531846 388170 531902 388226
rect 531474 388046 531530 388102
rect 531598 388046 531654 388102
rect 531722 388046 531778 388102
rect 531846 388046 531902 388102
rect 531474 387922 531530 387978
rect 531598 387922 531654 387978
rect 531722 387922 531778 387978
rect 531846 387922 531902 387978
rect 531474 370294 531530 370350
rect 531598 370294 531654 370350
rect 531722 370294 531778 370350
rect 531846 370294 531902 370350
rect 531474 370170 531530 370226
rect 531598 370170 531654 370226
rect 531722 370170 531778 370226
rect 531846 370170 531902 370226
rect 531474 370046 531530 370102
rect 531598 370046 531654 370102
rect 531722 370046 531778 370102
rect 531846 370046 531902 370102
rect 531474 369922 531530 369978
rect 531598 369922 531654 369978
rect 531722 369922 531778 369978
rect 531846 369922 531902 369978
rect 531474 352294 531530 352350
rect 531598 352294 531654 352350
rect 531722 352294 531778 352350
rect 531846 352294 531902 352350
rect 531474 352170 531530 352226
rect 531598 352170 531654 352226
rect 531722 352170 531778 352226
rect 531846 352170 531902 352226
rect 531474 352046 531530 352102
rect 531598 352046 531654 352102
rect 531722 352046 531778 352102
rect 531846 352046 531902 352102
rect 531474 351922 531530 351978
rect 531598 351922 531654 351978
rect 531722 351922 531778 351978
rect 531846 351922 531902 351978
rect 558474 400294 558530 400350
rect 558598 400294 558654 400350
rect 558722 400294 558778 400350
rect 558846 400294 558902 400350
rect 558474 400170 558530 400226
rect 558598 400170 558654 400226
rect 558722 400170 558778 400226
rect 558846 400170 558902 400226
rect 558474 400046 558530 400102
rect 558598 400046 558654 400102
rect 558722 400046 558778 400102
rect 558846 400046 558902 400102
rect 558474 399922 558530 399978
rect 558598 399922 558654 399978
rect 558722 399922 558778 399978
rect 558846 399922 558902 399978
rect 558474 382294 558530 382350
rect 558598 382294 558654 382350
rect 558722 382294 558778 382350
rect 558846 382294 558902 382350
rect 558474 382170 558530 382226
rect 558598 382170 558654 382226
rect 558722 382170 558778 382226
rect 558846 382170 558902 382226
rect 558474 382046 558530 382102
rect 558598 382046 558654 382102
rect 558722 382046 558778 382102
rect 558846 382046 558902 382102
rect 558474 381922 558530 381978
rect 558598 381922 558654 381978
rect 558722 381922 558778 381978
rect 558846 381922 558902 381978
rect 562194 598116 562250 598172
rect 562318 598116 562374 598172
rect 562442 598116 562498 598172
rect 562566 598116 562622 598172
rect 562194 597992 562250 598048
rect 562318 597992 562374 598048
rect 562442 597992 562498 598048
rect 562566 597992 562622 598048
rect 562194 597868 562250 597924
rect 562318 597868 562374 597924
rect 562442 597868 562498 597924
rect 562566 597868 562622 597924
rect 562194 597744 562250 597800
rect 562318 597744 562374 597800
rect 562442 597744 562498 597800
rect 562566 597744 562622 597800
rect 562194 586294 562250 586350
rect 562318 586294 562374 586350
rect 562442 586294 562498 586350
rect 562566 586294 562622 586350
rect 562194 586170 562250 586226
rect 562318 586170 562374 586226
rect 562442 586170 562498 586226
rect 562566 586170 562622 586226
rect 562194 586046 562250 586102
rect 562318 586046 562374 586102
rect 562442 586046 562498 586102
rect 562566 586046 562622 586102
rect 562194 585922 562250 585978
rect 562318 585922 562374 585978
rect 562442 585922 562498 585978
rect 562566 585922 562622 585978
rect 562194 568294 562250 568350
rect 562318 568294 562374 568350
rect 562442 568294 562498 568350
rect 562566 568294 562622 568350
rect 562194 568170 562250 568226
rect 562318 568170 562374 568226
rect 562442 568170 562498 568226
rect 562566 568170 562622 568226
rect 562194 568046 562250 568102
rect 562318 568046 562374 568102
rect 562442 568046 562498 568102
rect 562566 568046 562622 568102
rect 562194 567922 562250 567978
rect 562318 567922 562374 567978
rect 562442 567922 562498 567978
rect 562566 567922 562622 567978
rect 562194 550294 562250 550350
rect 562318 550294 562374 550350
rect 562442 550294 562498 550350
rect 562566 550294 562622 550350
rect 562194 550170 562250 550226
rect 562318 550170 562374 550226
rect 562442 550170 562498 550226
rect 562566 550170 562622 550226
rect 562194 550046 562250 550102
rect 562318 550046 562374 550102
rect 562442 550046 562498 550102
rect 562566 550046 562622 550102
rect 562194 549922 562250 549978
rect 562318 549922 562374 549978
rect 562442 549922 562498 549978
rect 562566 549922 562622 549978
rect 562194 532294 562250 532350
rect 562318 532294 562374 532350
rect 562442 532294 562498 532350
rect 562566 532294 562622 532350
rect 562194 532170 562250 532226
rect 562318 532170 562374 532226
rect 562442 532170 562498 532226
rect 562566 532170 562622 532226
rect 562194 532046 562250 532102
rect 562318 532046 562374 532102
rect 562442 532046 562498 532102
rect 562566 532046 562622 532102
rect 562194 531922 562250 531978
rect 562318 531922 562374 531978
rect 562442 531922 562498 531978
rect 562566 531922 562622 531978
rect 562194 514294 562250 514350
rect 562318 514294 562374 514350
rect 562442 514294 562498 514350
rect 562566 514294 562622 514350
rect 562194 514170 562250 514226
rect 562318 514170 562374 514226
rect 562442 514170 562498 514226
rect 562566 514170 562622 514226
rect 562194 514046 562250 514102
rect 562318 514046 562374 514102
rect 562442 514046 562498 514102
rect 562566 514046 562622 514102
rect 562194 513922 562250 513978
rect 562318 513922 562374 513978
rect 562442 513922 562498 513978
rect 562566 513922 562622 513978
rect 562194 496294 562250 496350
rect 562318 496294 562374 496350
rect 562442 496294 562498 496350
rect 562566 496294 562622 496350
rect 562194 496170 562250 496226
rect 562318 496170 562374 496226
rect 562442 496170 562498 496226
rect 562566 496170 562622 496226
rect 562194 496046 562250 496102
rect 562318 496046 562374 496102
rect 562442 496046 562498 496102
rect 562566 496046 562622 496102
rect 562194 495922 562250 495978
rect 562318 495922 562374 495978
rect 562442 495922 562498 495978
rect 562566 495922 562622 495978
rect 562194 478294 562250 478350
rect 562318 478294 562374 478350
rect 562442 478294 562498 478350
rect 562566 478294 562622 478350
rect 562194 478170 562250 478226
rect 562318 478170 562374 478226
rect 562442 478170 562498 478226
rect 562566 478170 562622 478226
rect 562194 478046 562250 478102
rect 562318 478046 562374 478102
rect 562442 478046 562498 478102
rect 562566 478046 562622 478102
rect 562194 477922 562250 477978
rect 562318 477922 562374 477978
rect 562442 477922 562498 477978
rect 562566 477922 562622 477978
rect 562194 460294 562250 460350
rect 562318 460294 562374 460350
rect 562442 460294 562498 460350
rect 562566 460294 562622 460350
rect 562194 460170 562250 460226
rect 562318 460170 562374 460226
rect 562442 460170 562498 460226
rect 562566 460170 562622 460226
rect 562194 460046 562250 460102
rect 562318 460046 562374 460102
rect 562442 460046 562498 460102
rect 562566 460046 562622 460102
rect 562194 459922 562250 459978
rect 562318 459922 562374 459978
rect 562442 459922 562498 459978
rect 562566 459922 562622 459978
rect 562194 442294 562250 442350
rect 562318 442294 562374 442350
rect 562442 442294 562498 442350
rect 562566 442294 562622 442350
rect 562194 442170 562250 442226
rect 562318 442170 562374 442226
rect 562442 442170 562498 442226
rect 562566 442170 562622 442226
rect 562194 442046 562250 442102
rect 562318 442046 562374 442102
rect 562442 442046 562498 442102
rect 562566 442046 562622 442102
rect 562194 441922 562250 441978
rect 562318 441922 562374 441978
rect 562442 441922 562498 441978
rect 562566 441922 562622 441978
rect 562194 424294 562250 424350
rect 562318 424294 562374 424350
rect 562442 424294 562498 424350
rect 562566 424294 562622 424350
rect 562194 424170 562250 424226
rect 562318 424170 562374 424226
rect 562442 424170 562498 424226
rect 562566 424170 562622 424226
rect 562194 424046 562250 424102
rect 562318 424046 562374 424102
rect 562442 424046 562498 424102
rect 562566 424046 562622 424102
rect 562194 423922 562250 423978
rect 562318 423922 562374 423978
rect 562442 423922 562498 423978
rect 562566 423922 562622 423978
rect 562194 406294 562250 406350
rect 562318 406294 562374 406350
rect 562442 406294 562498 406350
rect 562566 406294 562622 406350
rect 562194 406170 562250 406226
rect 562318 406170 562374 406226
rect 562442 406170 562498 406226
rect 562566 406170 562622 406226
rect 562194 406046 562250 406102
rect 562318 406046 562374 406102
rect 562442 406046 562498 406102
rect 562566 406046 562622 406102
rect 562194 405922 562250 405978
rect 562318 405922 562374 405978
rect 562442 405922 562498 405978
rect 562566 405922 562622 405978
rect 589194 597156 589250 597212
rect 589318 597156 589374 597212
rect 589442 597156 589498 597212
rect 589566 597156 589622 597212
rect 589194 597032 589250 597088
rect 589318 597032 589374 597088
rect 589442 597032 589498 597088
rect 589566 597032 589622 597088
rect 589194 596908 589250 596964
rect 589318 596908 589374 596964
rect 589442 596908 589498 596964
rect 589566 596908 589622 596964
rect 589194 596784 589250 596840
rect 589318 596784 589374 596840
rect 589442 596784 589498 596840
rect 589566 596784 589622 596840
rect 592914 598116 592970 598172
rect 593038 598116 593094 598172
rect 593162 598116 593218 598172
rect 593286 598116 593342 598172
rect 592914 597992 592970 598048
rect 593038 597992 593094 598048
rect 593162 597992 593218 598048
rect 593286 597992 593342 598048
rect 592914 597868 592970 597924
rect 593038 597868 593094 597924
rect 593162 597868 593218 597924
rect 593286 597868 593342 597924
rect 592914 597744 592970 597800
rect 593038 597744 593094 597800
rect 593162 597744 593218 597800
rect 593286 597744 593342 597800
rect 589194 580294 589250 580350
rect 589318 580294 589374 580350
rect 589442 580294 589498 580350
rect 589566 580294 589622 580350
rect 589194 580170 589250 580226
rect 589318 580170 589374 580226
rect 589442 580170 589498 580226
rect 589566 580170 589622 580226
rect 589194 580046 589250 580102
rect 589318 580046 589374 580102
rect 589442 580046 589498 580102
rect 589566 580046 589622 580102
rect 589194 579922 589250 579978
rect 589318 579922 589374 579978
rect 589442 579922 589498 579978
rect 589566 579922 589622 579978
rect 589194 562294 589250 562350
rect 589318 562294 589374 562350
rect 589442 562294 589498 562350
rect 589566 562294 589622 562350
rect 589194 562170 589250 562226
rect 589318 562170 589374 562226
rect 589442 562170 589498 562226
rect 589566 562170 589622 562226
rect 589194 562046 589250 562102
rect 589318 562046 589374 562102
rect 589442 562046 589498 562102
rect 589566 562046 589622 562102
rect 589194 561922 589250 561978
rect 589318 561922 589374 561978
rect 589442 561922 589498 561978
rect 589566 561922 589622 561978
rect 589194 544294 589250 544350
rect 589318 544294 589374 544350
rect 589442 544294 589498 544350
rect 589566 544294 589622 544350
rect 589194 544170 589250 544226
rect 589318 544170 589374 544226
rect 589442 544170 589498 544226
rect 589566 544170 589622 544226
rect 589194 544046 589250 544102
rect 589318 544046 589374 544102
rect 589442 544046 589498 544102
rect 589566 544046 589622 544102
rect 589194 543922 589250 543978
rect 589318 543922 589374 543978
rect 589442 543922 589498 543978
rect 589566 543922 589622 543978
rect 589194 526294 589250 526350
rect 589318 526294 589374 526350
rect 589442 526294 589498 526350
rect 589566 526294 589622 526350
rect 589194 526170 589250 526226
rect 589318 526170 589374 526226
rect 589442 526170 589498 526226
rect 589566 526170 589622 526226
rect 589194 526046 589250 526102
rect 589318 526046 589374 526102
rect 589442 526046 589498 526102
rect 589566 526046 589622 526102
rect 589194 525922 589250 525978
rect 589318 525922 589374 525978
rect 589442 525922 589498 525978
rect 589566 525922 589622 525978
rect 589194 508294 589250 508350
rect 589318 508294 589374 508350
rect 589442 508294 589498 508350
rect 589566 508294 589622 508350
rect 589194 508170 589250 508226
rect 589318 508170 589374 508226
rect 589442 508170 589498 508226
rect 589566 508170 589622 508226
rect 589194 508046 589250 508102
rect 589318 508046 589374 508102
rect 589442 508046 589498 508102
rect 589566 508046 589622 508102
rect 589194 507922 589250 507978
rect 589318 507922 589374 507978
rect 589442 507922 589498 507978
rect 589566 507922 589622 507978
rect 589194 490294 589250 490350
rect 589318 490294 589374 490350
rect 589442 490294 589498 490350
rect 589566 490294 589622 490350
rect 589194 490170 589250 490226
rect 589318 490170 589374 490226
rect 589442 490170 589498 490226
rect 589566 490170 589622 490226
rect 589194 490046 589250 490102
rect 589318 490046 589374 490102
rect 589442 490046 589498 490102
rect 589566 490046 589622 490102
rect 589194 489922 589250 489978
rect 589318 489922 589374 489978
rect 589442 489922 589498 489978
rect 589566 489922 589622 489978
rect 589194 472294 589250 472350
rect 589318 472294 589374 472350
rect 589442 472294 589498 472350
rect 589566 472294 589622 472350
rect 589194 472170 589250 472226
rect 589318 472170 589374 472226
rect 589442 472170 589498 472226
rect 589566 472170 589622 472226
rect 589194 472046 589250 472102
rect 589318 472046 589374 472102
rect 589442 472046 589498 472102
rect 589566 472046 589622 472102
rect 589194 471922 589250 471978
rect 589318 471922 589374 471978
rect 589442 471922 589498 471978
rect 589566 471922 589622 471978
rect 589194 454294 589250 454350
rect 589318 454294 589374 454350
rect 589442 454294 589498 454350
rect 589566 454294 589622 454350
rect 589194 454170 589250 454226
rect 589318 454170 589374 454226
rect 589442 454170 589498 454226
rect 589566 454170 589622 454226
rect 589194 454046 589250 454102
rect 589318 454046 589374 454102
rect 589442 454046 589498 454102
rect 589566 454046 589622 454102
rect 589194 453922 589250 453978
rect 589318 453922 589374 453978
rect 589442 453922 589498 453978
rect 589566 453922 589622 453978
rect 589194 436294 589250 436350
rect 589318 436294 589374 436350
rect 589442 436294 589498 436350
rect 589566 436294 589622 436350
rect 589194 436170 589250 436226
rect 589318 436170 589374 436226
rect 589442 436170 589498 436226
rect 589566 436170 589622 436226
rect 589194 436046 589250 436102
rect 589318 436046 589374 436102
rect 589442 436046 589498 436102
rect 589566 436046 589622 436102
rect 589194 435922 589250 435978
rect 589318 435922 589374 435978
rect 589442 435922 589498 435978
rect 589566 435922 589622 435978
rect 589194 418294 589250 418350
rect 589318 418294 589374 418350
rect 589442 418294 589498 418350
rect 589566 418294 589622 418350
rect 589194 418170 589250 418226
rect 589318 418170 589374 418226
rect 589442 418170 589498 418226
rect 589566 418170 589622 418226
rect 589194 418046 589250 418102
rect 589318 418046 589374 418102
rect 589442 418046 589498 418102
rect 589566 418046 589622 418102
rect 589194 417922 589250 417978
rect 589318 417922 589374 417978
rect 589442 417922 589498 417978
rect 589566 417922 589622 417978
rect 589194 400294 589250 400350
rect 589318 400294 589374 400350
rect 589442 400294 589498 400350
rect 589566 400294 589622 400350
rect 589194 400170 589250 400226
rect 589318 400170 589374 400226
rect 589442 400170 589498 400226
rect 589566 400170 589622 400226
rect 589194 400046 589250 400102
rect 589318 400046 589374 400102
rect 589442 400046 589498 400102
rect 589566 400046 589622 400102
rect 589194 399922 589250 399978
rect 589318 399922 589374 399978
rect 589442 399922 589498 399978
rect 589566 399922 589622 399978
rect 562194 388294 562250 388350
rect 562318 388294 562374 388350
rect 562442 388294 562498 388350
rect 562566 388294 562622 388350
rect 562194 388170 562250 388226
rect 562318 388170 562374 388226
rect 562442 388170 562498 388226
rect 562566 388170 562622 388226
rect 562194 388046 562250 388102
rect 562318 388046 562374 388102
rect 562442 388046 562498 388102
rect 562566 388046 562622 388102
rect 562194 387922 562250 387978
rect 562318 387922 562374 387978
rect 562442 387922 562498 387978
rect 562566 387922 562622 387978
rect 558474 364294 558530 364350
rect 558598 364294 558654 364350
rect 558722 364294 558778 364350
rect 558846 364294 558902 364350
rect 558474 364170 558530 364226
rect 558598 364170 558654 364226
rect 558722 364170 558778 364226
rect 558846 364170 558902 364226
rect 558474 364046 558530 364102
rect 558598 364046 558654 364102
rect 558722 364046 558778 364102
rect 558846 364046 558902 364102
rect 558474 363922 558530 363978
rect 558598 363922 558654 363978
rect 558722 363922 558778 363978
rect 558846 363922 558902 363978
rect 558474 346294 558530 346350
rect 558598 346294 558654 346350
rect 558722 346294 558778 346350
rect 558846 346294 558902 346350
rect 558474 346170 558530 346226
rect 558598 346170 558654 346226
rect 558722 346170 558778 346226
rect 558846 346170 558902 346226
rect 558474 346046 558530 346102
rect 558598 346046 558654 346102
rect 558722 346046 558778 346102
rect 558846 346046 558902 346102
rect 558474 345922 558530 345978
rect 558598 345922 558654 345978
rect 558722 345922 558778 345978
rect 558846 345922 558902 345978
rect 531474 334294 531530 334350
rect 531598 334294 531654 334350
rect 531722 334294 531778 334350
rect 531846 334294 531902 334350
rect 531474 334170 531530 334226
rect 531598 334170 531654 334226
rect 531722 334170 531778 334226
rect 531846 334170 531902 334226
rect 531474 334046 531530 334102
rect 531598 334046 531654 334102
rect 531722 334046 531778 334102
rect 531846 334046 531902 334102
rect 531474 333922 531530 333978
rect 531598 333922 531654 333978
rect 531722 333922 531778 333978
rect 531846 333922 531902 333978
rect 531474 316294 531530 316350
rect 531598 316294 531654 316350
rect 531722 316294 531778 316350
rect 531846 316294 531902 316350
rect 531474 316170 531530 316226
rect 531598 316170 531654 316226
rect 531722 316170 531778 316226
rect 531846 316170 531902 316226
rect 531474 316046 531530 316102
rect 531598 316046 531654 316102
rect 531722 316046 531778 316102
rect 531846 316046 531902 316102
rect 531474 315922 531530 315978
rect 531598 315922 531654 315978
rect 531722 315922 531778 315978
rect 531846 315922 531902 315978
rect 531474 298294 531530 298350
rect 531598 298294 531654 298350
rect 531722 298294 531778 298350
rect 531846 298294 531902 298350
rect 531474 298170 531530 298226
rect 531598 298170 531654 298226
rect 531722 298170 531778 298226
rect 531846 298170 531902 298226
rect 531474 298046 531530 298102
rect 531598 298046 531654 298102
rect 531722 298046 531778 298102
rect 531846 298046 531902 298102
rect 531474 297922 531530 297978
rect 531598 297922 531654 297978
rect 531722 297922 531778 297978
rect 531846 297922 531902 297978
rect 531474 280294 531530 280350
rect 531598 280294 531654 280350
rect 531722 280294 531778 280350
rect 531846 280294 531902 280350
rect 531474 280170 531530 280226
rect 531598 280170 531654 280226
rect 531722 280170 531778 280226
rect 531846 280170 531902 280226
rect 531474 280046 531530 280102
rect 531598 280046 531654 280102
rect 531722 280046 531778 280102
rect 531846 280046 531902 280102
rect 531474 279922 531530 279978
rect 531598 279922 531654 279978
rect 531722 279922 531778 279978
rect 531846 279922 531902 279978
rect 531474 262294 531530 262350
rect 531598 262294 531654 262350
rect 531722 262294 531778 262350
rect 531846 262294 531902 262350
rect 531474 262170 531530 262226
rect 531598 262170 531654 262226
rect 531722 262170 531778 262226
rect 531846 262170 531902 262226
rect 531474 262046 531530 262102
rect 531598 262046 531654 262102
rect 531722 262046 531778 262102
rect 531846 262046 531902 262102
rect 531474 261922 531530 261978
rect 531598 261922 531654 261978
rect 531722 261922 531778 261978
rect 531846 261922 531902 261978
rect 531474 244294 531530 244350
rect 531598 244294 531654 244350
rect 531722 244294 531778 244350
rect 531846 244294 531902 244350
rect 531474 244170 531530 244226
rect 531598 244170 531654 244226
rect 531722 244170 531778 244226
rect 531846 244170 531902 244226
rect 531474 244046 531530 244102
rect 531598 244046 531654 244102
rect 531722 244046 531778 244102
rect 531846 244046 531902 244102
rect 531474 243922 531530 243978
rect 531598 243922 531654 243978
rect 531722 243922 531778 243978
rect 531846 243922 531902 243978
rect 531474 226294 531530 226350
rect 531598 226294 531654 226350
rect 531722 226294 531778 226350
rect 531846 226294 531902 226350
rect 531474 226170 531530 226226
rect 531598 226170 531654 226226
rect 531722 226170 531778 226226
rect 531846 226170 531902 226226
rect 531474 226046 531530 226102
rect 531598 226046 531654 226102
rect 531722 226046 531778 226102
rect 531846 226046 531902 226102
rect 531474 225922 531530 225978
rect 531598 225922 531654 225978
rect 531722 225922 531778 225978
rect 531846 225922 531902 225978
rect 531474 208294 531530 208350
rect 531598 208294 531654 208350
rect 531722 208294 531778 208350
rect 531846 208294 531902 208350
rect 531474 208170 531530 208226
rect 531598 208170 531654 208226
rect 531722 208170 531778 208226
rect 531846 208170 531902 208226
rect 531474 208046 531530 208102
rect 531598 208046 531654 208102
rect 531722 208046 531778 208102
rect 531846 208046 531902 208102
rect 531474 207922 531530 207978
rect 531598 207922 531654 207978
rect 531722 207922 531778 207978
rect 531846 207922 531902 207978
rect 531474 190294 531530 190350
rect 531598 190294 531654 190350
rect 531722 190294 531778 190350
rect 531846 190294 531902 190350
rect 531474 190170 531530 190226
rect 531598 190170 531654 190226
rect 531722 190170 531778 190226
rect 531846 190170 531902 190226
rect 531474 190046 531530 190102
rect 531598 190046 531654 190102
rect 531722 190046 531778 190102
rect 531846 190046 531902 190102
rect 531474 189922 531530 189978
rect 531598 189922 531654 189978
rect 531722 189922 531778 189978
rect 531846 189922 531902 189978
rect 531474 172294 531530 172350
rect 531598 172294 531654 172350
rect 531722 172294 531778 172350
rect 531846 172294 531902 172350
rect 531474 172170 531530 172226
rect 531598 172170 531654 172226
rect 531722 172170 531778 172226
rect 531846 172170 531902 172226
rect 531474 172046 531530 172102
rect 531598 172046 531654 172102
rect 531722 172046 531778 172102
rect 531846 172046 531902 172102
rect 531474 171922 531530 171978
rect 531598 171922 531654 171978
rect 531722 171922 531778 171978
rect 531846 171922 531902 171978
rect 531474 154294 531530 154350
rect 531598 154294 531654 154350
rect 531722 154294 531778 154350
rect 531846 154294 531902 154350
rect 531474 154170 531530 154226
rect 531598 154170 531654 154226
rect 531722 154170 531778 154226
rect 531846 154170 531902 154226
rect 531474 154046 531530 154102
rect 531598 154046 531654 154102
rect 531722 154046 531778 154102
rect 531846 154046 531902 154102
rect 531474 153922 531530 153978
rect 531598 153922 531654 153978
rect 531722 153922 531778 153978
rect 531846 153922 531902 153978
rect 558474 328294 558530 328350
rect 558598 328294 558654 328350
rect 558722 328294 558778 328350
rect 558846 328294 558902 328350
rect 558474 328170 558530 328226
rect 558598 328170 558654 328226
rect 558722 328170 558778 328226
rect 558846 328170 558902 328226
rect 558474 328046 558530 328102
rect 558598 328046 558654 328102
rect 558722 328046 558778 328102
rect 558846 328046 558902 328102
rect 558474 327922 558530 327978
rect 558598 327922 558654 327978
rect 558722 327922 558778 327978
rect 558846 327922 558902 327978
rect 558474 310294 558530 310350
rect 558598 310294 558654 310350
rect 558722 310294 558778 310350
rect 558846 310294 558902 310350
rect 558474 310170 558530 310226
rect 558598 310170 558654 310226
rect 558722 310170 558778 310226
rect 558846 310170 558902 310226
rect 558474 310046 558530 310102
rect 558598 310046 558654 310102
rect 558722 310046 558778 310102
rect 558846 310046 558902 310102
rect 558474 309922 558530 309978
rect 558598 309922 558654 309978
rect 558722 309922 558778 309978
rect 558846 309922 558902 309978
rect 558474 292294 558530 292350
rect 558598 292294 558654 292350
rect 558722 292294 558778 292350
rect 558846 292294 558902 292350
rect 558474 292170 558530 292226
rect 558598 292170 558654 292226
rect 558722 292170 558778 292226
rect 558846 292170 558902 292226
rect 558474 292046 558530 292102
rect 558598 292046 558654 292102
rect 558722 292046 558778 292102
rect 558846 292046 558902 292102
rect 558474 291922 558530 291978
rect 558598 291922 558654 291978
rect 558722 291922 558778 291978
rect 558846 291922 558902 291978
rect 558474 274294 558530 274350
rect 558598 274294 558654 274350
rect 558722 274294 558778 274350
rect 558846 274294 558902 274350
rect 558474 274170 558530 274226
rect 558598 274170 558654 274226
rect 558722 274170 558778 274226
rect 558846 274170 558902 274226
rect 558474 274046 558530 274102
rect 558598 274046 558654 274102
rect 558722 274046 558778 274102
rect 558846 274046 558902 274102
rect 558474 273922 558530 273978
rect 558598 273922 558654 273978
rect 558722 273922 558778 273978
rect 558846 273922 558902 273978
rect 558474 256294 558530 256350
rect 558598 256294 558654 256350
rect 558722 256294 558778 256350
rect 558846 256294 558902 256350
rect 558474 256170 558530 256226
rect 558598 256170 558654 256226
rect 558722 256170 558778 256226
rect 558846 256170 558902 256226
rect 558474 256046 558530 256102
rect 558598 256046 558654 256102
rect 558722 256046 558778 256102
rect 558846 256046 558902 256102
rect 558474 255922 558530 255978
rect 558598 255922 558654 255978
rect 558722 255922 558778 255978
rect 558846 255922 558902 255978
rect 558474 238294 558530 238350
rect 558598 238294 558654 238350
rect 558722 238294 558778 238350
rect 558846 238294 558902 238350
rect 558474 238170 558530 238226
rect 558598 238170 558654 238226
rect 558722 238170 558778 238226
rect 558846 238170 558902 238226
rect 558474 238046 558530 238102
rect 558598 238046 558654 238102
rect 558722 238046 558778 238102
rect 558846 238046 558902 238102
rect 558474 237922 558530 237978
rect 558598 237922 558654 237978
rect 558722 237922 558778 237978
rect 558846 237922 558902 237978
rect 558474 220294 558530 220350
rect 558598 220294 558654 220350
rect 558722 220294 558778 220350
rect 558846 220294 558902 220350
rect 558474 220170 558530 220226
rect 558598 220170 558654 220226
rect 558722 220170 558778 220226
rect 558846 220170 558902 220226
rect 558474 220046 558530 220102
rect 558598 220046 558654 220102
rect 558722 220046 558778 220102
rect 558846 220046 558902 220102
rect 558474 219922 558530 219978
rect 558598 219922 558654 219978
rect 558722 219922 558778 219978
rect 558846 219922 558902 219978
rect 558474 202294 558530 202350
rect 558598 202294 558654 202350
rect 558722 202294 558778 202350
rect 558846 202294 558902 202350
rect 558474 202170 558530 202226
rect 558598 202170 558654 202226
rect 558722 202170 558778 202226
rect 558846 202170 558902 202226
rect 558474 202046 558530 202102
rect 558598 202046 558654 202102
rect 558722 202046 558778 202102
rect 558846 202046 558902 202102
rect 558474 201922 558530 201978
rect 558598 201922 558654 201978
rect 558722 201922 558778 201978
rect 558846 201922 558902 201978
rect 558474 184294 558530 184350
rect 558598 184294 558654 184350
rect 558722 184294 558778 184350
rect 558846 184294 558902 184350
rect 558474 184170 558530 184226
rect 558598 184170 558654 184226
rect 558722 184170 558778 184226
rect 558846 184170 558902 184226
rect 558474 184046 558530 184102
rect 558598 184046 558654 184102
rect 558722 184046 558778 184102
rect 558846 184046 558902 184102
rect 558474 183922 558530 183978
rect 558598 183922 558654 183978
rect 558722 183922 558778 183978
rect 558846 183922 558902 183978
rect 558474 166294 558530 166350
rect 558598 166294 558654 166350
rect 558722 166294 558778 166350
rect 558846 166294 558902 166350
rect 558474 166170 558530 166226
rect 558598 166170 558654 166226
rect 558722 166170 558778 166226
rect 558846 166170 558902 166226
rect 558474 166046 558530 166102
rect 558598 166046 558654 166102
rect 558722 166046 558778 166102
rect 558846 166046 558902 166102
rect 558474 165922 558530 165978
rect 558598 165922 558654 165978
rect 558722 165922 558778 165978
rect 558846 165922 558902 165978
rect 479878 136294 479934 136350
rect 480002 136294 480058 136350
rect 479878 136170 479934 136226
rect 480002 136170 480058 136226
rect 479878 136046 479934 136102
rect 480002 136046 480058 136102
rect 479878 135922 479934 135978
rect 480002 135922 480058 135978
rect 510598 136294 510654 136350
rect 510722 136294 510778 136350
rect 510598 136170 510654 136226
rect 510722 136170 510778 136226
rect 510598 136046 510654 136102
rect 510722 136046 510778 136102
rect 510598 135922 510654 135978
rect 510722 135922 510778 135978
rect 541318 136294 541374 136350
rect 541442 136294 541498 136350
rect 541318 136170 541374 136226
rect 541442 136170 541498 136226
rect 541318 136046 541374 136102
rect 541442 136046 541498 136102
rect 541318 135922 541374 135978
rect 541442 135922 541498 135978
rect 464518 130294 464574 130350
rect 464642 130294 464698 130350
rect 464518 130170 464574 130226
rect 464642 130170 464698 130226
rect 464518 130046 464574 130102
rect 464642 130046 464698 130102
rect 464518 129922 464574 129978
rect 464642 129922 464698 129978
rect 495238 130294 495294 130350
rect 495362 130294 495418 130350
rect 495238 130170 495294 130226
rect 495362 130170 495418 130226
rect 495238 130046 495294 130102
rect 495362 130046 495418 130102
rect 495238 129922 495294 129978
rect 495362 129922 495418 129978
rect 525958 130294 526014 130350
rect 526082 130294 526138 130350
rect 525958 130170 526014 130226
rect 526082 130170 526138 130226
rect 525958 130046 526014 130102
rect 526082 130046 526138 130102
rect 525958 129922 526014 129978
rect 526082 129922 526138 129978
rect 556678 130294 556734 130350
rect 556802 130294 556858 130350
rect 556678 130170 556734 130226
rect 556802 130170 556858 130226
rect 556678 130046 556734 130102
rect 556802 130046 556858 130102
rect 556678 129922 556734 129978
rect 556802 129922 556858 129978
rect 479878 118294 479934 118350
rect 480002 118294 480058 118350
rect 479878 118170 479934 118226
rect 480002 118170 480058 118226
rect 479878 118046 479934 118102
rect 480002 118046 480058 118102
rect 479878 117922 479934 117978
rect 480002 117922 480058 117978
rect 510598 118294 510654 118350
rect 510722 118294 510778 118350
rect 510598 118170 510654 118226
rect 510722 118170 510778 118226
rect 510598 118046 510654 118102
rect 510722 118046 510778 118102
rect 510598 117922 510654 117978
rect 510722 117922 510778 117978
rect 541318 118294 541374 118350
rect 541442 118294 541498 118350
rect 541318 118170 541374 118226
rect 541442 118170 541498 118226
rect 541318 118046 541374 118102
rect 541442 118046 541498 118102
rect 541318 117922 541374 117978
rect 541442 117922 541498 117978
rect 464518 112294 464574 112350
rect 464642 112294 464698 112350
rect 464518 112170 464574 112226
rect 464642 112170 464698 112226
rect 464518 112046 464574 112102
rect 464642 112046 464698 112102
rect 464518 111922 464574 111978
rect 464642 111922 464698 111978
rect 495238 112294 495294 112350
rect 495362 112294 495418 112350
rect 495238 112170 495294 112226
rect 495362 112170 495418 112226
rect 495238 112046 495294 112102
rect 495362 112046 495418 112102
rect 495238 111922 495294 111978
rect 495362 111922 495418 111978
rect 525958 112294 526014 112350
rect 526082 112294 526138 112350
rect 525958 112170 526014 112226
rect 526082 112170 526138 112226
rect 525958 112046 526014 112102
rect 526082 112046 526138 112102
rect 525958 111922 526014 111978
rect 526082 111922 526138 111978
rect 556678 112294 556734 112350
rect 556802 112294 556858 112350
rect 556678 112170 556734 112226
rect 556802 112170 556858 112226
rect 556678 112046 556734 112102
rect 556802 112046 556858 112102
rect 556678 111922 556734 111978
rect 556802 111922 556858 111978
rect 479878 100294 479934 100350
rect 480002 100294 480058 100350
rect 479878 100170 479934 100226
rect 480002 100170 480058 100226
rect 479878 100046 479934 100102
rect 480002 100046 480058 100102
rect 479878 99922 479934 99978
rect 480002 99922 480058 99978
rect 510598 100294 510654 100350
rect 510722 100294 510778 100350
rect 510598 100170 510654 100226
rect 510722 100170 510778 100226
rect 510598 100046 510654 100102
rect 510722 100046 510778 100102
rect 510598 99922 510654 99978
rect 510722 99922 510778 99978
rect 541318 100294 541374 100350
rect 541442 100294 541498 100350
rect 541318 100170 541374 100226
rect 541442 100170 541498 100226
rect 541318 100046 541374 100102
rect 541442 100046 541498 100102
rect 541318 99922 541374 99978
rect 541442 99922 541498 99978
rect 464518 94294 464574 94350
rect 464642 94294 464698 94350
rect 464518 94170 464574 94226
rect 464642 94170 464698 94226
rect 464518 94046 464574 94102
rect 464642 94046 464698 94102
rect 464518 93922 464574 93978
rect 464642 93922 464698 93978
rect 495238 94294 495294 94350
rect 495362 94294 495418 94350
rect 495238 94170 495294 94226
rect 495362 94170 495418 94226
rect 495238 94046 495294 94102
rect 495362 94046 495418 94102
rect 495238 93922 495294 93978
rect 495362 93922 495418 93978
rect 525958 94294 526014 94350
rect 526082 94294 526138 94350
rect 525958 94170 526014 94226
rect 526082 94170 526138 94226
rect 525958 94046 526014 94102
rect 526082 94046 526138 94102
rect 525958 93922 526014 93978
rect 526082 93922 526138 93978
rect 556678 94294 556734 94350
rect 556802 94294 556858 94350
rect 556678 94170 556734 94226
rect 556802 94170 556858 94226
rect 556678 94046 556734 94102
rect 556802 94046 556858 94102
rect 556678 93922 556734 93978
rect 556802 93922 556858 93978
rect 479878 82294 479934 82350
rect 480002 82294 480058 82350
rect 479878 82170 479934 82226
rect 480002 82170 480058 82226
rect 479878 82046 479934 82102
rect 480002 82046 480058 82102
rect 479878 81922 479934 81978
rect 480002 81922 480058 81978
rect 510598 82294 510654 82350
rect 510722 82294 510778 82350
rect 510598 82170 510654 82226
rect 510722 82170 510778 82226
rect 510598 82046 510654 82102
rect 510722 82046 510778 82102
rect 510598 81922 510654 81978
rect 510722 81922 510778 81978
rect 541318 82294 541374 82350
rect 541442 82294 541498 82350
rect 541318 82170 541374 82226
rect 541442 82170 541498 82226
rect 541318 82046 541374 82102
rect 541442 82046 541498 82102
rect 541318 81922 541374 81978
rect 541442 81922 541498 81978
rect 464518 76294 464574 76350
rect 464642 76294 464698 76350
rect 464518 76170 464574 76226
rect 464642 76170 464698 76226
rect 464518 76046 464574 76102
rect 464642 76046 464698 76102
rect 464518 75922 464574 75978
rect 464642 75922 464698 75978
rect 495238 76294 495294 76350
rect 495362 76294 495418 76350
rect 495238 76170 495294 76226
rect 495362 76170 495418 76226
rect 495238 76046 495294 76102
rect 495362 76046 495418 76102
rect 495238 75922 495294 75978
rect 495362 75922 495418 75978
rect 525958 76294 526014 76350
rect 526082 76294 526138 76350
rect 525958 76170 526014 76226
rect 526082 76170 526138 76226
rect 525958 76046 526014 76102
rect 526082 76046 526138 76102
rect 525958 75922 526014 75978
rect 526082 75922 526138 75978
rect 556678 76294 556734 76350
rect 556802 76294 556858 76350
rect 556678 76170 556734 76226
rect 556802 76170 556858 76226
rect 556678 76046 556734 76102
rect 556802 76046 556858 76102
rect 556678 75922 556734 75978
rect 556802 75922 556858 75978
rect 562194 370294 562250 370350
rect 562318 370294 562374 370350
rect 562442 370294 562498 370350
rect 562566 370294 562622 370350
rect 562194 370170 562250 370226
rect 562318 370170 562374 370226
rect 562442 370170 562498 370226
rect 562566 370170 562622 370226
rect 562194 370046 562250 370102
rect 562318 370046 562374 370102
rect 562442 370046 562498 370102
rect 562566 370046 562622 370102
rect 562194 369922 562250 369978
rect 562318 369922 562374 369978
rect 562442 369922 562498 369978
rect 562566 369922 562622 369978
rect 577052 389762 577108 389818
rect 562194 352294 562250 352350
rect 562318 352294 562374 352350
rect 562442 352294 562498 352350
rect 562566 352294 562622 352350
rect 562194 352170 562250 352226
rect 562318 352170 562374 352226
rect 562442 352170 562498 352226
rect 562566 352170 562622 352226
rect 562194 352046 562250 352102
rect 562318 352046 562374 352102
rect 562442 352046 562498 352102
rect 562566 352046 562622 352102
rect 562194 351922 562250 351978
rect 562318 351922 562374 351978
rect 562442 351922 562498 351978
rect 562566 351922 562622 351978
rect 562194 334294 562250 334350
rect 562318 334294 562374 334350
rect 562442 334294 562498 334350
rect 562566 334294 562622 334350
rect 562194 334170 562250 334226
rect 562318 334170 562374 334226
rect 562442 334170 562498 334226
rect 562566 334170 562622 334226
rect 562194 334046 562250 334102
rect 562318 334046 562374 334102
rect 562442 334046 562498 334102
rect 562566 334046 562622 334102
rect 562194 333922 562250 333978
rect 562318 333922 562374 333978
rect 562442 333922 562498 333978
rect 562566 333922 562622 333978
rect 562194 316294 562250 316350
rect 562318 316294 562374 316350
rect 562442 316294 562498 316350
rect 562566 316294 562622 316350
rect 562194 316170 562250 316226
rect 562318 316170 562374 316226
rect 562442 316170 562498 316226
rect 562566 316170 562622 316226
rect 562194 316046 562250 316102
rect 562318 316046 562374 316102
rect 562442 316046 562498 316102
rect 562566 316046 562622 316102
rect 562194 315922 562250 315978
rect 562318 315922 562374 315978
rect 562442 315922 562498 315978
rect 562566 315922 562622 315978
rect 562194 298294 562250 298350
rect 562318 298294 562374 298350
rect 562442 298294 562498 298350
rect 562566 298294 562622 298350
rect 562194 298170 562250 298226
rect 562318 298170 562374 298226
rect 562442 298170 562498 298226
rect 562566 298170 562622 298226
rect 562194 298046 562250 298102
rect 562318 298046 562374 298102
rect 562442 298046 562498 298102
rect 562566 298046 562622 298102
rect 562194 297922 562250 297978
rect 562318 297922 562374 297978
rect 562442 297922 562498 297978
rect 562566 297922 562622 297978
rect 562194 280294 562250 280350
rect 562318 280294 562374 280350
rect 562442 280294 562498 280350
rect 562566 280294 562622 280350
rect 562194 280170 562250 280226
rect 562318 280170 562374 280226
rect 562442 280170 562498 280226
rect 562566 280170 562622 280226
rect 562194 280046 562250 280102
rect 562318 280046 562374 280102
rect 562442 280046 562498 280102
rect 562566 280046 562622 280102
rect 562194 279922 562250 279978
rect 562318 279922 562374 279978
rect 562442 279922 562498 279978
rect 562566 279922 562622 279978
rect 562194 262294 562250 262350
rect 562318 262294 562374 262350
rect 562442 262294 562498 262350
rect 562566 262294 562622 262350
rect 562194 262170 562250 262226
rect 562318 262170 562374 262226
rect 562442 262170 562498 262226
rect 562566 262170 562622 262226
rect 562194 262046 562250 262102
rect 562318 262046 562374 262102
rect 562442 262046 562498 262102
rect 562566 262046 562622 262102
rect 562194 261922 562250 261978
rect 562318 261922 562374 261978
rect 562442 261922 562498 261978
rect 562566 261922 562622 261978
rect 562194 244294 562250 244350
rect 562318 244294 562374 244350
rect 562442 244294 562498 244350
rect 562566 244294 562622 244350
rect 562194 244170 562250 244226
rect 562318 244170 562374 244226
rect 562442 244170 562498 244226
rect 562566 244170 562622 244226
rect 562194 244046 562250 244102
rect 562318 244046 562374 244102
rect 562442 244046 562498 244102
rect 562566 244046 562622 244102
rect 562194 243922 562250 243978
rect 562318 243922 562374 243978
rect 562442 243922 562498 243978
rect 562566 243922 562622 243978
rect 562194 226294 562250 226350
rect 562318 226294 562374 226350
rect 562442 226294 562498 226350
rect 562566 226294 562622 226350
rect 562194 226170 562250 226226
rect 562318 226170 562374 226226
rect 562442 226170 562498 226226
rect 562566 226170 562622 226226
rect 562194 226046 562250 226102
rect 562318 226046 562374 226102
rect 562442 226046 562498 226102
rect 562566 226046 562622 226102
rect 562194 225922 562250 225978
rect 562318 225922 562374 225978
rect 562442 225922 562498 225978
rect 562566 225922 562622 225978
rect 562194 208294 562250 208350
rect 562318 208294 562374 208350
rect 562442 208294 562498 208350
rect 562566 208294 562622 208350
rect 562194 208170 562250 208226
rect 562318 208170 562374 208226
rect 562442 208170 562498 208226
rect 562566 208170 562622 208226
rect 562194 208046 562250 208102
rect 562318 208046 562374 208102
rect 562442 208046 562498 208102
rect 562566 208046 562622 208102
rect 562194 207922 562250 207978
rect 562318 207922 562374 207978
rect 562442 207922 562498 207978
rect 562566 207922 562622 207978
rect 562194 190294 562250 190350
rect 562318 190294 562374 190350
rect 562442 190294 562498 190350
rect 562566 190294 562622 190350
rect 562194 190170 562250 190226
rect 562318 190170 562374 190226
rect 562442 190170 562498 190226
rect 562566 190170 562622 190226
rect 562194 190046 562250 190102
rect 562318 190046 562374 190102
rect 562442 190046 562498 190102
rect 562566 190046 562622 190102
rect 562194 189922 562250 189978
rect 562318 189922 562374 189978
rect 562442 189922 562498 189978
rect 562566 189922 562622 189978
rect 562194 172294 562250 172350
rect 562318 172294 562374 172350
rect 562442 172294 562498 172350
rect 562566 172294 562622 172350
rect 562194 172170 562250 172226
rect 562318 172170 562374 172226
rect 562442 172170 562498 172226
rect 562566 172170 562622 172226
rect 562194 172046 562250 172102
rect 562318 172046 562374 172102
rect 562442 172046 562498 172102
rect 562566 172046 562622 172102
rect 562194 171922 562250 171978
rect 562318 171922 562374 171978
rect 562442 171922 562498 171978
rect 562566 171922 562622 171978
rect 562194 154294 562250 154350
rect 562318 154294 562374 154350
rect 562442 154294 562498 154350
rect 562566 154294 562622 154350
rect 562194 154170 562250 154226
rect 562318 154170 562374 154226
rect 562442 154170 562498 154226
rect 562566 154170 562622 154226
rect 562194 154046 562250 154102
rect 562318 154046 562374 154102
rect 562442 154046 562498 154102
rect 562566 154046 562622 154102
rect 562194 153922 562250 153978
rect 562318 153922 562374 153978
rect 562442 153922 562498 153978
rect 562566 153922 562622 153978
rect 562194 136294 562250 136350
rect 562318 136294 562374 136350
rect 562442 136294 562498 136350
rect 562566 136294 562622 136350
rect 562194 136170 562250 136226
rect 562318 136170 562374 136226
rect 562442 136170 562498 136226
rect 562566 136170 562622 136226
rect 562194 136046 562250 136102
rect 562318 136046 562374 136102
rect 562442 136046 562498 136102
rect 562566 136046 562622 136102
rect 562194 135922 562250 135978
rect 562318 135922 562374 135978
rect 562442 135922 562498 135978
rect 562566 135922 562622 135978
rect 562194 118294 562250 118350
rect 562318 118294 562374 118350
rect 562442 118294 562498 118350
rect 562566 118294 562622 118350
rect 562194 118170 562250 118226
rect 562318 118170 562374 118226
rect 562442 118170 562498 118226
rect 562566 118170 562622 118226
rect 562194 118046 562250 118102
rect 562318 118046 562374 118102
rect 562442 118046 562498 118102
rect 562566 118046 562622 118102
rect 562194 117922 562250 117978
rect 562318 117922 562374 117978
rect 562442 117922 562498 117978
rect 562566 117922 562622 117978
rect 562194 100294 562250 100350
rect 562318 100294 562374 100350
rect 562442 100294 562498 100350
rect 562566 100294 562622 100350
rect 562194 100170 562250 100226
rect 562318 100170 562374 100226
rect 562442 100170 562498 100226
rect 562566 100170 562622 100226
rect 562194 100046 562250 100102
rect 562318 100046 562374 100102
rect 562442 100046 562498 100102
rect 562566 100046 562622 100102
rect 562194 99922 562250 99978
rect 562318 99922 562374 99978
rect 562442 99922 562498 99978
rect 562566 99922 562622 99978
rect 562194 82294 562250 82350
rect 562318 82294 562374 82350
rect 562442 82294 562498 82350
rect 562566 82294 562622 82350
rect 562194 82170 562250 82226
rect 562318 82170 562374 82226
rect 562442 82170 562498 82226
rect 562566 82170 562622 82226
rect 562194 82046 562250 82102
rect 562318 82046 562374 82102
rect 562442 82046 562498 82102
rect 562566 82046 562622 82102
rect 562194 81922 562250 81978
rect 562318 81922 562374 81978
rect 562442 81922 562498 81978
rect 562566 81922 562622 81978
rect 479878 64294 479934 64350
rect 480002 64294 480058 64350
rect 479878 64170 479934 64226
rect 480002 64170 480058 64226
rect 479878 64046 479934 64102
rect 480002 64046 480058 64102
rect 479878 63922 479934 63978
rect 480002 63922 480058 63978
rect 510598 64294 510654 64350
rect 510722 64294 510778 64350
rect 510598 64170 510654 64226
rect 510722 64170 510778 64226
rect 510598 64046 510654 64102
rect 510722 64046 510778 64102
rect 510598 63922 510654 63978
rect 510722 63922 510778 63978
rect 541318 64294 541374 64350
rect 541442 64294 541498 64350
rect 541318 64170 541374 64226
rect 541442 64170 541498 64226
rect 541318 64046 541374 64102
rect 541442 64046 541498 64102
rect 541318 63922 541374 63978
rect 541442 63922 541498 63978
rect 562194 64294 562250 64350
rect 562318 64294 562374 64350
rect 562442 64294 562498 64350
rect 562566 64294 562622 64350
rect 562194 64170 562250 64226
rect 562318 64170 562374 64226
rect 562442 64170 562498 64226
rect 562566 64170 562622 64226
rect 562194 64046 562250 64102
rect 562318 64046 562374 64102
rect 562442 64046 562498 64102
rect 562566 64046 562622 64102
rect 562194 63922 562250 63978
rect 562318 63922 562374 63978
rect 562442 63922 562498 63978
rect 562566 63922 562622 63978
rect 464518 58294 464574 58350
rect 464642 58294 464698 58350
rect 464518 58170 464574 58226
rect 464642 58170 464698 58226
rect 464518 58046 464574 58102
rect 464642 58046 464698 58102
rect 464518 57922 464574 57978
rect 464642 57922 464698 57978
rect 495238 58294 495294 58350
rect 495362 58294 495418 58350
rect 495238 58170 495294 58226
rect 495362 58170 495418 58226
rect 495238 58046 495294 58102
rect 495362 58046 495418 58102
rect 495238 57922 495294 57978
rect 495362 57922 495418 57978
rect 525958 58294 526014 58350
rect 526082 58294 526138 58350
rect 525958 58170 526014 58226
rect 526082 58170 526138 58226
rect 525958 58046 526014 58102
rect 526082 58046 526138 58102
rect 525958 57922 526014 57978
rect 526082 57922 526138 57978
rect 556678 58294 556734 58350
rect 556802 58294 556858 58350
rect 556678 58170 556734 58226
rect 556802 58170 556858 58226
rect 556678 58046 556734 58102
rect 556802 58046 556858 58102
rect 556678 57922 556734 57978
rect 556802 57922 556858 57978
rect 439314 46294 439370 46350
rect 439438 46294 439494 46350
rect 439562 46294 439618 46350
rect 439686 46294 439742 46350
rect 439314 46170 439370 46226
rect 439438 46170 439494 46226
rect 439562 46170 439618 46226
rect 439686 46170 439742 46226
rect 439314 46046 439370 46102
rect 439438 46046 439494 46102
rect 439562 46046 439618 46102
rect 439686 46046 439742 46102
rect 439314 45922 439370 45978
rect 439438 45922 439494 45978
rect 439562 45922 439618 45978
rect 439686 45922 439742 45978
rect 439314 28294 439370 28350
rect 439438 28294 439494 28350
rect 439562 28294 439618 28350
rect 439686 28294 439742 28350
rect 439314 28170 439370 28226
rect 439438 28170 439494 28226
rect 439562 28170 439618 28226
rect 439686 28170 439742 28226
rect 439314 28046 439370 28102
rect 439438 28046 439494 28102
rect 439562 28046 439618 28102
rect 439686 28046 439742 28102
rect 439314 27922 439370 27978
rect 439438 27922 439494 27978
rect 439562 27922 439618 27978
rect 439686 27922 439742 27978
rect 439314 10294 439370 10350
rect 439438 10294 439494 10350
rect 439562 10294 439618 10350
rect 439686 10294 439742 10350
rect 439314 10170 439370 10226
rect 439438 10170 439494 10226
rect 439562 10170 439618 10226
rect 439686 10170 439742 10226
rect 439314 10046 439370 10102
rect 439438 10046 439494 10102
rect 439562 10046 439618 10102
rect 439686 10046 439742 10102
rect 439314 9922 439370 9978
rect 439438 9922 439494 9978
rect 439562 9922 439618 9978
rect 439686 9922 439742 9978
rect 439314 -1176 439370 -1120
rect 439438 -1176 439494 -1120
rect 439562 -1176 439618 -1120
rect 439686 -1176 439742 -1120
rect 439314 -1300 439370 -1244
rect 439438 -1300 439494 -1244
rect 439562 -1300 439618 -1244
rect 439686 -1300 439742 -1244
rect 439314 -1424 439370 -1368
rect 439438 -1424 439494 -1368
rect 439562 -1424 439618 -1368
rect 439686 -1424 439742 -1368
rect 439314 -1548 439370 -1492
rect 439438 -1548 439494 -1492
rect 439562 -1548 439618 -1492
rect 439686 -1548 439742 -1492
rect 466314 40294 466370 40350
rect 466438 40294 466494 40350
rect 466562 40294 466618 40350
rect 466686 40294 466742 40350
rect 466314 40170 466370 40226
rect 466438 40170 466494 40226
rect 466562 40170 466618 40226
rect 466686 40170 466742 40226
rect 466314 40046 466370 40102
rect 466438 40046 466494 40102
rect 466562 40046 466618 40102
rect 466686 40046 466742 40102
rect 466314 39922 466370 39978
rect 466438 39922 466494 39978
rect 466562 39922 466618 39978
rect 466686 39922 466742 39978
rect 466314 22294 466370 22350
rect 466438 22294 466494 22350
rect 466562 22294 466618 22350
rect 466686 22294 466742 22350
rect 466314 22170 466370 22226
rect 466438 22170 466494 22226
rect 466562 22170 466618 22226
rect 466686 22170 466742 22226
rect 466314 22046 466370 22102
rect 466438 22046 466494 22102
rect 466562 22046 466618 22102
rect 466686 22046 466742 22102
rect 466314 21922 466370 21978
rect 466438 21922 466494 21978
rect 466562 21922 466618 21978
rect 466686 21922 466742 21978
rect 466314 4294 466370 4350
rect 466438 4294 466494 4350
rect 466562 4294 466618 4350
rect 466686 4294 466742 4350
rect 466314 4170 466370 4226
rect 466438 4170 466494 4226
rect 466562 4170 466618 4226
rect 466686 4170 466742 4226
rect 466314 4046 466370 4102
rect 466438 4046 466494 4102
rect 466562 4046 466618 4102
rect 466686 4046 466742 4102
rect 466314 3922 466370 3978
rect 466438 3922 466494 3978
rect 466562 3922 466618 3978
rect 466686 3922 466742 3978
rect 466314 -216 466370 -160
rect 466438 -216 466494 -160
rect 466562 -216 466618 -160
rect 466686 -216 466742 -160
rect 466314 -340 466370 -284
rect 466438 -340 466494 -284
rect 466562 -340 466618 -284
rect 466686 -340 466742 -284
rect 466314 -464 466370 -408
rect 466438 -464 466494 -408
rect 466562 -464 466618 -408
rect 466686 -464 466742 -408
rect 466314 -588 466370 -532
rect 466438 -588 466494 -532
rect 466562 -588 466618 -532
rect 466686 -588 466742 -532
rect 470034 46294 470090 46350
rect 470158 46294 470214 46350
rect 470282 46294 470338 46350
rect 470406 46294 470462 46350
rect 470034 46170 470090 46226
rect 470158 46170 470214 46226
rect 470282 46170 470338 46226
rect 470406 46170 470462 46226
rect 470034 46046 470090 46102
rect 470158 46046 470214 46102
rect 470282 46046 470338 46102
rect 470406 46046 470462 46102
rect 470034 45922 470090 45978
rect 470158 45922 470214 45978
rect 470282 45922 470338 45978
rect 470406 45922 470462 45978
rect 470034 28294 470090 28350
rect 470158 28294 470214 28350
rect 470282 28294 470338 28350
rect 470406 28294 470462 28350
rect 470034 28170 470090 28226
rect 470158 28170 470214 28226
rect 470282 28170 470338 28226
rect 470406 28170 470462 28226
rect 470034 28046 470090 28102
rect 470158 28046 470214 28102
rect 470282 28046 470338 28102
rect 470406 28046 470462 28102
rect 470034 27922 470090 27978
rect 470158 27922 470214 27978
rect 470282 27922 470338 27978
rect 470406 27922 470462 27978
rect 470034 10294 470090 10350
rect 470158 10294 470214 10350
rect 470282 10294 470338 10350
rect 470406 10294 470462 10350
rect 470034 10170 470090 10226
rect 470158 10170 470214 10226
rect 470282 10170 470338 10226
rect 470406 10170 470462 10226
rect 470034 10046 470090 10102
rect 470158 10046 470214 10102
rect 470282 10046 470338 10102
rect 470406 10046 470462 10102
rect 470034 9922 470090 9978
rect 470158 9922 470214 9978
rect 470282 9922 470338 9978
rect 470406 9922 470462 9978
rect 470034 -1176 470090 -1120
rect 470158 -1176 470214 -1120
rect 470282 -1176 470338 -1120
rect 470406 -1176 470462 -1120
rect 470034 -1300 470090 -1244
rect 470158 -1300 470214 -1244
rect 470282 -1300 470338 -1244
rect 470406 -1300 470462 -1244
rect 470034 -1424 470090 -1368
rect 470158 -1424 470214 -1368
rect 470282 -1424 470338 -1368
rect 470406 -1424 470462 -1368
rect 470034 -1548 470090 -1492
rect 470158 -1548 470214 -1492
rect 470282 -1548 470338 -1492
rect 470406 -1548 470462 -1492
rect 497034 40294 497090 40350
rect 497158 40294 497214 40350
rect 497282 40294 497338 40350
rect 497406 40294 497462 40350
rect 497034 40170 497090 40226
rect 497158 40170 497214 40226
rect 497282 40170 497338 40226
rect 497406 40170 497462 40226
rect 497034 40046 497090 40102
rect 497158 40046 497214 40102
rect 497282 40046 497338 40102
rect 497406 40046 497462 40102
rect 497034 39922 497090 39978
rect 497158 39922 497214 39978
rect 497282 39922 497338 39978
rect 497406 39922 497462 39978
rect 497034 22294 497090 22350
rect 497158 22294 497214 22350
rect 497282 22294 497338 22350
rect 497406 22294 497462 22350
rect 497034 22170 497090 22226
rect 497158 22170 497214 22226
rect 497282 22170 497338 22226
rect 497406 22170 497462 22226
rect 497034 22046 497090 22102
rect 497158 22046 497214 22102
rect 497282 22046 497338 22102
rect 497406 22046 497462 22102
rect 497034 21922 497090 21978
rect 497158 21922 497214 21978
rect 497282 21922 497338 21978
rect 497406 21922 497462 21978
rect 497034 4294 497090 4350
rect 497158 4294 497214 4350
rect 497282 4294 497338 4350
rect 497406 4294 497462 4350
rect 497034 4170 497090 4226
rect 497158 4170 497214 4226
rect 497282 4170 497338 4226
rect 497406 4170 497462 4226
rect 497034 4046 497090 4102
rect 497158 4046 497214 4102
rect 497282 4046 497338 4102
rect 497406 4046 497462 4102
rect 497034 3922 497090 3978
rect 497158 3922 497214 3978
rect 497282 3922 497338 3978
rect 497406 3922 497462 3978
rect 497034 -216 497090 -160
rect 497158 -216 497214 -160
rect 497282 -216 497338 -160
rect 497406 -216 497462 -160
rect 497034 -340 497090 -284
rect 497158 -340 497214 -284
rect 497282 -340 497338 -284
rect 497406 -340 497462 -284
rect 497034 -464 497090 -408
rect 497158 -464 497214 -408
rect 497282 -464 497338 -408
rect 497406 -464 497462 -408
rect 497034 -588 497090 -532
rect 497158 -588 497214 -532
rect 497282 -588 497338 -532
rect 497406 -588 497462 -532
rect 500754 46294 500810 46350
rect 500878 46294 500934 46350
rect 501002 46294 501058 46350
rect 501126 46294 501182 46350
rect 500754 46170 500810 46226
rect 500878 46170 500934 46226
rect 501002 46170 501058 46226
rect 501126 46170 501182 46226
rect 500754 46046 500810 46102
rect 500878 46046 500934 46102
rect 501002 46046 501058 46102
rect 501126 46046 501182 46102
rect 500754 45922 500810 45978
rect 500878 45922 500934 45978
rect 501002 45922 501058 45978
rect 501126 45922 501182 45978
rect 500754 28294 500810 28350
rect 500878 28294 500934 28350
rect 501002 28294 501058 28350
rect 501126 28294 501182 28350
rect 500754 28170 500810 28226
rect 500878 28170 500934 28226
rect 501002 28170 501058 28226
rect 501126 28170 501182 28226
rect 500754 28046 500810 28102
rect 500878 28046 500934 28102
rect 501002 28046 501058 28102
rect 501126 28046 501182 28102
rect 500754 27922 500810 27978
rect 500878 27922 500934 27978
rect 501002 27922 501058 27978
rect 501126 27922 501182 27978
rect 500754 10294 500810 10350
rect 500878 10294 500934 10350
rect 501002 10294 501058 10350
rect 501126 10294 501182 10350
rect 500754 10170 500810 10226
rect 500878 10170 500934 10226
rect 501002 10170 501058 10226
rect 501126 10170 501182 10226
rect 500754 10046 500810 10102
rect 500878 10046 500934 10102
rect 501002 10046 501058 10102
rect 501126 10046 501182 10102
rect 500754 9922 500810 9978
rect 500878 9922 500934 9978
rect 501002 9922 501058 9978
rect 501126 9922 501182 9978
rect 500754 -1176 500810 -1120
rect 500878 -1176 500934 -1120
rect 501002 -1176 501058 -1120
rect 501126 -1176 501182 -1120
rect 500754 -1300 500810 -1244
rect 500878 -1300 500934 -1244
rect 501002 -1300 501058 -1244
rect 501126 -1300 501182 -1244
rect 500754 -1424 500810 -1368
rect 500878 -1424 500934 -1368
rect 501002 -1424 501058 -1368
rect 501126 -1424 501182 -1368
rect 500754 -1548 500810 -1492
rect 500878 -1548 500934 -1492
rect 501002 -1548 501058 -1492
rect 501126 -1548 501182 -1492
rect 527754 40294 527810 40350
rect 527878 40294 527934 40350
rect 528002 40294 528058 40350
rect 528126 40294 528182 40350
rect 527754 40170 527810 40226
rect 527878 40170 527934 40226
rect 528002 40170 528058 40226
rect 528126 40170 528182 40226
rect 527754 40046 527810 40102
rect 527878 40046 527934 40102
rect 528002 40046 528058 40102
rect 528126 40046 528182 40102
rect 527754 39922 527810 39978
rect 527878 39922 527934 39978
rect 528002 39922 528058 39978
rect 528126 39922 528182 39978
rect 527754 22294 527810 22350
rect 527878 22294 527934 22350
rect 528002 22294 528058 22350
rect 528126 22294 528182 22350
rect 527754 22170 527810 22226
rect 527878 22170 527934 22226
rect 528002 22170 528058 22226
rect 528126 22170 528182 22226
rect 527754 22046 527810 22102
rect 527878 22046 527934 22102
rect 528002 22046 528058 22102
rect 528126 22046 528182 22102
rect 527754 21922 527810 21978
rect 527878 21922 527934 21978
rect 528002 21922 528058 21978
rect 528126 21922 528182 21978
rect 527754 4294 527810 4350
rect 527878 4294 527934 4350
rect 528002 4294 528058 4350
rect 528126 4294 528182 4350
rect 527754 4170 527810 4226
rect 527878 4170 527934 4226
rect 528002 4170 528058 4226
rect 528126 4170 528182 4226
rect 527754 4046 527810 4102
rect 527878 4046 527934 4102
rect 528002 4046 528058 4102
rect 528126 4046 528182 4102
rect 527754 3922 527810 3978
rect 527878 3922 527934 3978
rect 528002 3922 528058 3978
rect 528126 3922 528182 3978
rect 527754 -216 527810 -160
rect 527878 -216 527934 -160
rect 528002 -216 528058 -160
rect 528126 -216 528182 -160
rect 527754 -340 527810 -284
rect 527878 -340 527934 -284
rect 528002 -340 528058 -284
rect 528126 -340 528182 -284
rect 527754 -464 527810 -408
rect 527878 -464 527934 -408
rect 528002 -464 528058 -408
rect 528126 -464 528182 -408
rect 527754 -588 527810 -532
rect 527878 -588 527934 -532
rect 528002 -588 528058 -532
rect 528126 -588 528182 -532
rect 531474 46294 531530 46350
rect 531598 46294 531654 46350
rect 531722 46294 531778 46350
rect 531846 46294 531902 46350
rect 531474 46170 531530 46226
rect 531598 46170 531654 46226
rect 531722 46170 531778 46226
rect 531846 46170 531902 46226
rect 531474 46046 531530 46102
rect 531598 46046 531654 46102
rect 531722 46046 531778 46102
rect 531846 46046 531902 46102
rect 531474 45922 531530 45978
rect 531598 45922 531654 45978
rect 531722 45922 531778 45978
rect 531846 45922 531902 45978
rect 531474 28294 531530 28350
rect 531598 28294 531654 28350
rect 531722 28294 531778 28350
rect 531846 28294 531902 28350
rect 531474 28170 531530 28226
rect 531598 28170 531654 28226
rect 531722 28170 531778 28226
rect 531846 28170 531902 28226
rect 531474 28046 531530 28102
rect 531598 28046 531654 28102
rect 531722 28046 531778 28102
rect 531846 28046 531902 28102
rect 531474 27922 531530 27978
rect 531598 27922 531654 27978
rect 531722 27922 531778 27978
rect 531846 27922 531902 27978
rect 531474 10294 531530 10350
rect 531598 10294 531654 10350
rect 531722 10294 531778 10350
rect 531846 10294 531902 10350
rect 531474 10170 531530 10226
rect 531598 10170 531654 10226
rect 531722 10170 531778 10226
rect 531846 10170 531902 10226
rect 531474 10046 531530 10102
rect 531598 10046 531654 10102
rect 531722 10046 531778 10102
rect 531846 10046 531902 10102
rect 531474 9922 531530 9978
rect 531598 9922 531654 9978
rect 531722 9922 531778 9978
rect 531846 9922 531902 9978
rect 531474 -1176 531530 -1120
rect 531598 -1176 531654 -1120
rect 531722 -1176 531778 -1120
rect 531846 -1176 531902 -1120
rect 531474 -1300 531530 -1244
rect 531598 -1300 531654 -1244
rect 531722 -1300 531778 -1244
rect 531846 -1300 531902 -1244
rect 531474 -1424 531530 -1368
rect 531598 -1424 531654 -1368
rect 531722 -1424 531778 -1368
rect 531846 -1424 531902 -1368
rect 531474 -1548 531530 -1492
rect 531598 -1548 531654 -1492
rect 531722 -1548 531778 -1492
rect 531846 -1548 531902 -1492
rect 558474 40294 558530 40350
rect 558598 40294 558654 40350
rect 558722 40294 558778 40350
rect 558846 40294 558902 40350
rect 558474 40170 558530 40226
rect 558598 40170 558654 40226
rect 558722 40170 558778 40226
rect 558846 40170 558902 40226
rect 558474 40046 558530 40102
rect 558598 40046 558654 40102
rect 558722 40046 558778 40102
rect 558846 40046 558902 40102
rect 558474 39922 558530 39978
rect 558598 39922 558654 39978
rect 558722 39922 558778 39978
rect 558846 39922 558902 39978
rect 558474 22294 558530 22350
rect 558598 22294 558654 22350
rect 558722 22294 558778 22350
rect 558846 22294 558902 22350
rect 558474 22170 558530 22226
rect 558598 22170 558654 22226
rect 558722 22170 558778 22226
rect 558846 22170 558902 22226
rect 558474 22046 558530 22102
rect 558598 22046 558654 22102
rect 558722 22046 558778 22102
rect 558846 22046 558902 22102
rect 558474 21922 558530 21978
rect 558598 21922 558654 21978
rect 558722 21922 558778 21978
rect 558846 21922 558902 21978
rect 558474 4294 558530 4350
rect 558598 4294 558654 4350
rect 558722 4294 558778 4350
rect 558846 4294 558902 4350
rect 558474 4170 558530 4226
rect 558598 4170 558654 4226
rect 558722 4170 558778 4226
rect 558846 4170 558902 4226
rect 558474 4046 558530 4102
rect 558598 4046 558654 4102
rect 558722 4046 558778 4102
rect 558846 4046 558902 4102
rect 558474 3922 558530 3978
rect 558598 3922 558654 3978
rect 558722 3922 558778 3978
rect 558846 3922 558902 3978
rect 558474 -216 558530 -160
rect 558598 -216 558654 -160
rect 558722 -216 558778 -160
rect 558846 -216 558902 -160
rect 558474 -340 558530 -284
rect 558598 -340 558654 -284
rect 558722 -340 558778 -284
rect 558846 -340 558902 -284
rect 558474 -464 558530 -408
rect 558598 -464 558654 -408
rect 558722 -464 558778 -408
rect 558846 -464 558902 -408
rect 558474 -588 558530 -532
rect 558598 -588 558654 -532
rect 558722 -588 558778 -532
rect 558846 -588 558902 -532
rect 582988 385442 583044 385498
rect 579628 385262 579684 385318
rect 562194 46294 562250 46350
rect 562318 46294 562374 46350
rect 562442 46294 562498 46350
rect 562566 46294 562622 46350
rect 562194 46170 562250 46226
rect 562318 46170 562374 46226
rect 562442 46170 562498 46226
rect 562566 46170 562622 46226
rect 562194 46046 562250 46102
rect 562318 46046 562374 46102
rect 562442 46046 562498 46102
rect 562566 46046 562622 46102
rect 562194 45922 562250 45978
rect 562318 45922 562374 45978
rect 562442 45922 562498 45978
rect 562566 45922 562622 45978
rect 562194 28294 562250 28350
rect 562318 28294 562374 28350
rect 562442 28294 562498 28350
rect 562566 28294 562622 28350
rect 562194 28170 562250 28226
rect 562318 28170 562374 28226
rect 562442 28170 562498 28226
rect 562566 28170 562622 28226
rect 562194 28046 562250 28102
rect 562318 28046 562374 28102
rect 562442 28046 562498 28102
rect 562566 28046 562622 28102
rect 562194 27922 562250 27978
rect 562318 27922 562374 27978
rect 562442 27922 562498 27978
rect 562566 27922 562622 27978
rect 562194 10294 562250 10350
rect 562318 10294 562374 10350
rect 562442 10294 562498 10350
rect 562566 10294 562622 10350
rect 562194 10170 562250 10226
rect 562318 10170 562374 10226
rect 562442 10170 562498 10226
rect 562566 10170 562622 10226
rect 562194 10046 562250 10102
rect 562318 10046 562374 10102
rect 562442 10046 562498 10102
rect 562566 10046 562622 10102
rect 562194 9922 562250 9978
rect 562318 9922 562374 9978
rect 562442 9922 562498 9978
rect 562566 9922 562622 9978
rect 597456 598116 597512 598172
rect 597580 598116 597636 598172
rect 597704 598116 597760 598172
rect 597828 598116 597884 598172
rect 597456 597992 597512 598048
rect 597580 597992 597636 598048
rect 597704 597992 597760 598048
rect 597828 597992 597884 598048
rect 597456 597868 597512 597924
rect 597580 597868 597636 597924
rect 597704 597868 597760 597924
rect 597828 597868 597884 597924
rect 597456 597744 597512 597800
rect 597580 597744 597636 597800
rect 597704 597744 597760 597800
rect 597828 597744 597884 597800
rect 592914 586294 592970 586350
rect 593038 586294 593094 586350
rect 593162 586294 593218 586350
rect 593286 586294 593342 586350
rect 592914 586170 592970 586226
rect 593038 586170 593094 586226
rect 593162 586170 593218 586226
rect 593286 586170 593342 586226
rect 592914 586046 592970 586102
rect 593038 586046 593094 586102
rect 593162 586046 593218 586102
rect 593286 586046 593342 586102
rect 592914 585922 592970 585978
rect 593038 585922 593094 585978
rect 593162 585922 593218 585978
rect 593286 585922 593342 585978
rect 592914 568294 592970 568350
rect 593038 568294 593094 568350
rect 593162 568294 593218 568350
rect 593286 568294 593342 568350
rect 592914 568170 592970 568226
rect 593038 568170 593094 568226
rect 593162 568170 593218 568226
rect 593286 568170 593342 568226
rect 592914 568046 592970 568102
rect 593038 568046 593094 568102
rect 593162 568046 593218 568102
rect 593286 568046 593342 568102
rect 592914 567922 592970 567978
rect 593038 567922 593094 567978
rect 593162 567922 593218 567978
rect 593286 567922 593342 567978
rect 592914 550294 592970 550350
rect 593038 550294 593094 550350
rect 593162 550294 593218 550350
rect 593286 550294 593342 550350
rect 592914 550170 592970 550226
rect 593038 550170 593094 550226
rect 593162 550170 593218 550226
rect 593286 550170 593342 550226
rect 592914 550046 592970 550102
rect 593038 550046 593094 550102
rect 593162 550046 593218 550102
rect 593286 550046 593342 550102
rect 592914 549922 592970 549978
rect 593038 549922 593094 549978
rect 593162 549922 593218 549978
rect 593286 549922 593342 549978
rect 592914 532294 592970 532350
rect 593038 532294 593094 532350
rect 593162 532294 593218 532350
rect 593286 532294 593342 532350
rect 592914 532170 592970 532226
rect 593038 532170 593094 532226
rect 593162 532170 593218 532226
rect 593286 532170 593342 532226
rect 592914 532046 592970 532102
rect 593038 532046 593094 532102
rect 593162 532046 593218 532102
rect 593286 532046 593342 532102
rect 592914 531922 592970 531978
rect 593038 531922 593094 531978
rect 593162 531922 593218 531978
rect 593286 531922 593342 531978
rect 592914 514294 592970 514350
rect 593038 514294 593094 514350
rect 593162 514294 593218 514350
rect 593286 514294 593342 514350
rect 592914 514170 592970 514226
rect 593038 514170 593094 514226
rect 593162 514170 593218 514226
rect 593286 514170 593342 514226
rect 592914 514046 592970 514102
rect 593038 514046 593094 514102
rect 593162 514046 593218 514102
rect 593286 514046 593342 514102
rect 592914 513922 592970 513978
rect 593038 513922 593094 513978
rect 593162 513922 593218 513978
rect 593286 513922 593342 513978
rect 592914 496294 592970 496350
rect 593038 496294 593094 496350
rect 593162 496294 593218 496350
rect 593286 496294 593342 496350
rect 592914 496170 592970 496226
rect 593038 496170 593094 496226
rect 593162 496170 593218 496226
rect 593286 496170 593342 496226
rect 592914 496046 592970 496102
rect 593038 496046 593094 496102
rect 593162 496046 593218 496102
rect 593286 496046 593342 496102
rect 592914 495922 592970 495978
rect 593038 495922 593094 495978
rect 593162 495922 593218 495978
rect 593286 495922 593342 495978
rect 592914 478294 592970 478350
rect 593038 478294 593094 478350
rect 593162 478294 593218 478350
rect 593286 478294 593342 478350
rect 592914 478170 592970 478226
rect 593038 478170 593094 478226
rect 593162 478170 593218 478226
rect 593286 478170 593342 478226
rect 592914 478046 592970 478102
rect 593038 478046 593094 478102
rect 593162 478046 593218 478102
rect 593286 478046 593342 478102
rect 592914 477922 592970 477978
rect 593038 477922 593094 477978
rect 593162 477922 593218 477978
rect 593286 477922 593342 477978
rect 592914 460294 592970 460350
rect 593038 460294 593094 460350
rect 593162 460294 593218 460350
rect 593286 460294 593342 460350
rect 592914 460170 592970 460226
rect 593038 460170 593094 460226
rect 593162 460170 593218 460226
rect 593286 460170 593342 460226
rect 592914 460046 592970 460102
rect 593038 460046 593094 460102
rect 593162 460046 593218 460102
rect 593286 460046 593342 460102
rect 592914 459922 592970 459978
rect 593038 459922 593094 459978
rect 593162 459922 593218 459978
rect 593286 459922 593342 459978
rect 592914 442294 592970 442350
rect 593038 442294 593094 442350
rect 593162 442294 593218 442350
rect 593286 442294 593342 442350
rect 592914 442170 592970 442226
rect 593038 442170 593094 442226
rect 593162 442170 593218 442226
rect 593286 442170 593342 442226
rect 592914 442046 592970 442102
rect 593038 442046 593094 442102
rect 593162 442046 593218 442102
rect 593286 442046 593342 442102
rect 592914 441922 592970 441978
rect 593038 441922 593094 441978
rect 593162 441922 593218 441978
rect 593286 441922 593342 441978
rect 590828 403982 590884 404038
rect 592914 424294 592970 424350
rect 593038 424294 593094 424350
rect 593162 424294 593218 424350
rect 593286 424294 593342 424350
rect 592914 424170 592970 424226
rect 593038 424170 593094 424226
rect 593162 424170 593218 424226
rect 593286 424170 593342 424226
rect 592914 424046 592970 424102
rect 593038 424046 593094 424102
rect 593162 424046 593218 424102
rect 593286 424046 593342 424102
rect 592914 423922 592970 423978
rect 593038 423922 593094 423978
rect 593162 423922 593218 423978
rect 593286 423922 593342 423978
rect 592914 406294 592970 406350
rect 593038 406294 593094 406350
rect 593162 406294 593218 406350
rect 593286 406294 593342 406350
rect 592914 406170 592970 406226
rect 593038 406170 593094 406226
rect 593162 406170 593218 406226
rect 593286 406170 593342 406226
rect 592914 406046 592970 406102
rect 593038 406046 593094 406102
rect 593162 406046 593218 406102
rect 593286 406046 593342 406102
rect 592914 405922 592970 405978
rect 593038 405922 593094 405978
rect 593162 405922 593218 405978
rect 593286 405922 593342 405978
rect 592914 388294 592970 388350
rect 593038 388294 593094 388350
rect 593162 388294 593218 388350
rect 593286 388294 593342 388350
rect 592914 388170 592970 388226
rect 593038 388170 593094 388226
rect 593162 388170 593218 388226
rect 593286 388170 593342 388226
rect 592914 388046 592970 388102
rect 593038 388046 593094 388102
rect 593162 388046 593218 388102
rect 593286 388046 593342 388102
rect 592914 387922 592970 387978
rect 593038 387922 593094 387978
rect 593162 387922 593218 387978
rect 593286 387922 593342 387978
rect 589194 382294 589250 382350
rect 589318 382294 589374 382350
rect 589442 382294 589498 382350
rect 589566 382294 589622 382350
rect 589194 382170 589250 382226
rect 589318 382170 589374 382226
rect 589442 382170 589498 382226
rect 589566 382170 589622 382226
rect 589194 382046 589250 382102
rect 589318 382046 589374 382102
rect 589442 382046 589498 382102
rect 589566 382046 589622 382102
rect 589194 381922 589250 381978
rect 589318 381922 589374 381978
rect 589442 381922 589498 381978
rect 589566 381922 589622 381978
rect 589194 364294 589250 364350
rect 589318 364294 589374 364350
rect 589442 364294 589498 364350
rect 589566 364294 589622 364350
rect 589194 364170 589250 364226
rect 589318 364170 589374 364226
rect 589442 364170 589498 364226
rect 589566 364170 589622 364226
rect 589194 364046 589250 364102
rect 589318 364046 589374 364102
rect 589442 364046 589498 364102
rect 589566 364046 589622 364102
rect 589194 363922 589250 363978
rect 589318 363922 589374 363978
rect 589442 363922 589498 363978
rect 589566 363922 589622 363978
rect 592914 370294 592970 370350
rect 593038 370294 593094 370350
rect 593162 370294 593218 370350
rect 593286 370294 593342 370350
rect 592914 370170 592970 370226
rect 593038 370170 593094 370226
rect 593162 370170 593218 370226
rect 593286 370170 593342 370226
rect 592914 370046 592970 370102
rect 593038 370046 593094 370102
rect 593162 370046 593218 370102
rect 593286 370046 593342 370102
rect 592914 369922 592970 369978
rect 593038 369922 593094 369978
rect 593162 369922 593218 369978
rect 593286 369922 593342 369978
rect 592914 352294 592970 352350
rect 593038 352294 593094 352350
rect 593162 352294 593218 352350
rect 593286 352294 593342 352350
rect 592914 352170 592970 352226
rect 593038 352170 593094 352226
rect 593162 352170 593218 352226
rect 593286 352170 593342 352226
rect 592914 352046 592970 352102
rect 593038 352046 593094 352102
rect 593162 352046 593218 352102
rect 593286 352046 593342 352102
rect 592914 351922 592970 351978
rect 593038 351922 593094 351978
rect 593162 351922 593218 351978
rect 593286 351922 593342 351978
rect 589194 346294 589250 346350
rect 589318 346294 589374 346350
rect 589442 346294 589498 346350
rect 589566 346294 589622 346350
rect 589194 346170 589250 346226
rect 589318 346170 589374 346226
rect 589442 346170 589498 346226
rect 589566 346170 589622 346226
rect 589194 346046 589250 346102
rect 589318 346046 589374 346102
rect 589442 346046 589498 346102
rect 589566 346046 589622 346102
rect 589194 345922 589250 345978
rect 589318 345922 589374 345978
rect 589442 345922 589498 345978
rect 589566 345922 589622 345978
rect 589194 328294 589250 328350
rect 589318 328294 589374 328350
rect 589442 328294 589498 328350
rect 589566 328294 589622 328350
rect 589194 328170 589250 328226
rect 589318 328170 589374 328226
rect 589442 328170 589498 328226
rect 589566 328170 589622 328226
rect 589194 328046 589250 328102
rect 589318 328046 589374 328102
rect 589442 328046 589498 328102
rect 589566 328046 589622 328102
rect 589194 327922 589250 327978
rect 589318 327922 589374 327978
rect 589442 327922 589498 327978
rect 589566 327922 589622 327978
rect 589194 310294 589250 310350
rect 589318 310294 589374 310350
rect 589442 310294 589498 310350
rect 589566 310294 589622 310350
rect 589194 310170 589250 310226
rect 589318 310170 589374 310226
rect 589442 310170 589498 310226
rect 589566 310170 589622 310226
rect 589194 310046 589250 310102
rect 589318 310046 589374 310102
rect 589442 310046 589498 310102
rect 589566 310046 589622 310102
rect 589194 309922 589250 309978
rect 589318 309922 589374 309978
rect 589442 309922 589498 309978
rect 589566 309922 589622 309978
rect 589194 292294 589250 292350
rect 589318 292294 589374 292350
rect 589442 292294 589498 292350
rect 589566 292294 589622 292350
rect 589194 292170 589250 292226
rect 589318 292170 589374 292226
rect 589442 292170 589498 292226
rect 589566 292170 589622 292226
rect 589194 292046 589250 292102
rect 589318 292046 589374 292102
rect 589442 292046 589498 292102
rect 589566 292046 589622 292102
rect 589194 291922 589250 291978
rect 589318 291922 589374 291978
rect 589442 291922 589498 291978
rect 589566 291922 589622 291978
rect 589194 274294 589250 274350
rect 589318 274294 589374 274350
rect 589442 274294 589498 274350
rect 589566 274294 589622 274350
rect 589194 274170 589250 274226
rect 589318 274170 589374 274226
rect 589442 274170 589498 274226
rect 589566 274170 589622 274226
rect 589194 274046 589250 274102
rect 589318 274046 589374 274102
rect 589442 274046 589498 274102
rect 589566 274046 589622 274102
rect 589194 273922 589250 273978
rect 589318 273922 589374 273978
rect 589442 273922 589498 273978
rect 589566 273922 589622 273978
rect 592914 334294 592970 334350
rect 593038 334294 593094 334350
rect 593162 334294 593218 334350
rect 593286 334294 593342 334350
rect 592914 334170 592970 334226
rect 593038 334170 593094 334226
rect 593162 334170 593218 334226
rect 593286 334170 593342 334226
rect 592914 334046 592970 334102
rect 593038 334046 593094 334102
rect 593162 334046 593218 334102
rect 593286 334046 593342 334102
rect 592914 333922 592970 333978
rect 593038 333922 593094 333978
rect 593162 333922 593218 333978
rect 593286 333922 593342 333978
rect 592914 316294 592970 316350
rect 593038 316294 593094 316350
rect 593162 316294 593218 316350
rect 593286 316294 593342 316350
rect 592914 316170 592970 316226
rect 593038 316170 593094 316226
rect 593162 316170 593218 316226
rect 593286 316170 593342 316226
rect 592914 316046 592970 316102
rect 593038 316046 593094 316102
rect 593162 316046 593218 316102
rect 593286 316046 593342 316102
rect 592914 315922 592970 315978
rect 593038 315922 593094 315978
rect 593162 315922 593218 315978
rect 593286 315922 593342 315978
rect 589194 256294 589250 256350
rect 589318 256294 589374 256350
rect 589442 256294 589498 256350
rect 589566 256294 589622 256350
rect 589194 256170 589250 256226
rect 589318 256170 589374 256226
rect 589442 256170 589498 256226
rect 589566 256170 589622 256226
rect 589194 256046 589250 256102
rect 589318 256046 589374 256102
rect 589442 256046 589498 256102
rect 589566 256046 589622 256102
rect 589194 255922 589250 255978
rect 589318 255922 589374 255978
rect 589442 255922 589498 255978
rect 589566 255922 589622 255978
rect 592914 298294 592970 298350
rect 593038 298294 593094 298350
rect 593162 298294 593218 298350
rect 593286 298294 593342 298350
rect 592914 298170 592970 298226
rect 593038 298170 593094 298226
rect 593162 298170 593218 298226
rect 593286 298170 593342 298226
rect 592914 298046 592970 298102
rect 593038 298046 593094 298102
rect 593162 298046 593218 298102
rect 593286 298046 593342 298102
rect 592914 297922 592970 297978
rect 593038 297922 593094 297978
rect 593162 297922 593218 297978
rect 593286 297922 593342 297978
rect 592914 280294 592970 280350
rect 593038 280294 593094 280350
rect 593162 280294 593218 280350
rect 593286 280294 593342 280350
rect 592914 280170 592970 280226
rect 593038 280170 593094 280226
rect 593162 280170 593218 280226
rect 593286 280170 593342 280226
rect 592914 280046 592970 280102
rect 593038 280046 593094 280102
rect 593162 280046 593218 280102
rect 593286 280046 593342 280102
rect 592914 279922 592970 279978
rect 593038 279922 593094 279978
rect 593162 279922 593218 279978
rect 593286 279922 593342 279978
rect 592914 262294 592970 262350
rect 593038 262294 593094 262350
rect 593162 262294 593218 262350
rect 593286 262294 593342 262350
rect 592914 262170 592970 262226
rect 593038 262170 593094 262226
rect 593162 262170 593218 262226
rect 593286 262170 593342 262226
rect 592914 262046 592970 262102
rect 593038 262046 593094 262102
rect 593162 262046 593218 262102
rect 593286 262046 593342 262102
rect 592914 261922 592970 261978
rect 593038 261922 593094 261978
rect 593162 261922 593218 261978
rect 593286 261922 593342 261978
rect 592914 244294 592970 244350
rect 593038 244294 593094 244350
rect 593162 244294 593218 244350
rect 593286 244294 593342 244350
rect 592914 244170 592970 244226
rect 593038 244170 593094 244226
rect 593162 244170 593218 244226
rect 593286 244170 593342 244226
rect 592914 244046 592970 244102
rect 593038 244046 593094 244102
rect 593162 244046 593218 244102
rect 593286 244046 593342 244102
rect 592914 243922 592970 243978
rect 593038 243922 593094 243978
rect 593162 243922 593218 243978
rect 593286 243922 593342 243978
rect 589194 238294 589250 238350
rect 589318 238294 589374 238350
rect 589442 238294 589498 238350
rect 589566 238294 589622 238350
rect 589194 238170 589250 238226
rect 589318 238170 589374 238226
rect 589442 238170 589498 238226
rect 589566 238170 589622 238226
rect 589194 238046 589250 238102
rect 589318 238046 589374 238102
rect 589442 238046 589498 238102
rect 589566 238046 589622 238102
rect 589194 237922 589250 237978
rect 589318 237922 589374 237978
rect 589442 237922 589498 237978
rect 589566 237922 589622 237978
rect 589194 220294 589250 220350
rect 589318 220294 589374 220350
rect 589442 220294 589498 220350
rect 589566 220294 589622 220350
rect 589194 220170 589250 220226
rect 589318 220170 589374 220226
rect 589442 220170 589498 220226
rect 589566 220170 589622 220226
rect 589194 220046 589250 220102
rect 589318 220046 589374 220102
rect 589442 220046 589498 220102
rect 589566 220046 589622 220102
rect 589194 219922 589250 219978
rect 589318 219922 589374 219978
rect 589442 219922 589498 219978
rect 589566 219922 589622 219978
rect 589194 202294 589250 202350
rect 589318 202294 589374 202350
rect 589442 202294 589498 202350
rect 589566 202294 589622 202350
rect 589194 202170 589250 202226
rect 589318 202170 589374 202226
rect 589442 202170 589498 202226
rect 589566 202170 589622 202226
rect 589194 202046 589250 202102
rect 589318 202046 589374 202102
rect 589442 202046 589498 202102
rect 589566 202046 589622 202102
rect 589194 201922 589250 201978
rect 589318 201922 589374 201978
rect 589442 201922 589498 201978
rect 589566 201922 589622 201978
rect 589194 184294 589250 184350
rect 589318 184294 589374 184350
rect 589442 184294 589498 184350
rect 589566 184294 589622 184350
rect 589194 184170 589250 184226
rect 589318 184170 589374 184226
rect 589442 184170 589498 184226
rect 589566 184170 589622 184226
rect 589194 184046 589250 184102
rect 589318 184046 589374 184102
rect 589442 184046 589498 184102
rect 589566 184046 589622 184102
rect 589194 183922 589250 183978
rect 589318 183922 589374 183978
rect 589442 183922 589498 183978
rect 589566 183922 589622 183978
rect 589194 166294 589250 166350
rect 589318 166294 589374 166350
rect 589442 166294 589498 166350
rect 589566 166294 589622 166350
rect 589194 166170 589250 166226
rect 589318 166170 589374 166226
rect 589442 166170 589498 166226
rect 589566 166170 589622 166226
rect 589194 166046 589250 166102
rect 589318 166046 589374 166102
rect 589442 166046 589498 166102
rect 589566 166046 589622 166102
rect 589194 165922 589250 165978
rect 589318 165922 589374 165978
rect 589442 165922 589498 165978
rect 589566 165922 589622 165978
rect 589194 148294 589250 148350
rect 589318 148294 589374 148350
rect 589442 148294 589498 148350
rect 589566 148294 589622 148350
rect 589194 148170 589250 148226
rect 589318 148170 589374 148226
rect 589442 148170 589498 148226
rect 589566 148170 589622 148226
rect 589194 148046 589250 148102
rect 589318 148046 589374 148102
rect 589442 148046 589498 148102
rect 589566 148046 589622 148102
rect 589194 147922 589250 147978
rect 589318 147922 589374 147978
rect 589442 147922 589498 147978
rect 589566 147922 589622 147978
rect 589194 130294 589250 130350
rect 589318 130294 589374 130350
rect 589442 130294 589498 130350
rect 589566 130294 589622 130350
rect 589194 130170 589250 130226
rect 589318 130170 589374 130226
rect 589442 130170 589498 130226
rect 589566 130170 589622 130226
rect 589194 130046 589250 130102
rect 589318 130046 589374 130102
rect 589442 130046 589498 130102
rect 589566 130046 589622 130102
rect 589194 129922 589250 129978
rect 589318 129922 589374 129978
rect 589442 129922 589498 129978
rect 589566 129922 589622 129978
rect 589194 112294 589250 112350
rect 589318 112294 589374 112350
rect 589442 112294 589498 112350
rect 589566 112294 589622 112350
rect 589194 112170 589250 112226
rect 589318 112170 589374 112226
rect 589442 112170 589498 112226
rect 589566 112170 589622 112226
rect 589194 112046 589250 112102
rect 589318 112046 589374 112102
rect 589442 112046 589498 112102
rect 589566 112046 589622 112102
rect 589194 111922 589250 111978
rect 589318 111922 589374 111978
rect 589442 111922 589498 111978
rect 589566 111922 589622 111978
rect 589194 94294 589250 94350
rect 589318 94294 589374 94350
rect 589442 94294 589498 94350
rect 589566 94294 589622 94350
rect 589194 94170 589250 94226
rect 589318 94170 589374 94226
rect 589442 94170 589498 94226
rect 589566 94170 589622 94226
rect 589194 94046 589250 94102
rect 589318 94046 589374 94102
rect 589442 94046 589498 94102
rect 589566 94046 589622 94102
rect 589194 93922 589250 93978
rect 589318 93922 589374 93978
rect 589442 93922 589498 93978
rect 589566 93922 589622 93978
rect 589194 76294 589250 76350
rect 589318 76294 589374 76350
rect 589442 76294 589498 76350
rect 589566 76294 589622 76350
rect 589194 76170 589250 76226
rect 589318 76170 589374 76226
rect 589442 76170 589498 76226
rect 589566 76170 589622 76226
rect 589194 76046 589250 76102
rect 589318 76046 589374 76102
rect 589442 76046 589498 76102
rect 589566 76046 589622 76102
rect 589194 75922 589250 75978
rect 589318 75922 589374 75978
rect 589442 75922 589498 75978
rect 589566 75922 589622 75978
rect 592914 226294 592970 226350
rect 593038 226294 593094 226350
rect 593162 226294 593218 226350
rect 593286 226294 593342 226350
rect 592914 226170 592970 226226
rect 593038 226170 593094 226226
rect 593162 226170 593218 226226
rect 593286 226170 593342 226226
rect 592914 226046 592970 226102
rect 593038 226046 593094 226102
rect 593162 226046 593218 226102
rect 593286 226046 593342 226102
rect 592914 225922 592970 225978
rect 593038 225922 593094 225978
rect 593162 225922 593218 225978
rect 593286 225922 593342 225978
rect 592914 208294 592970 208350
rect 593038 208294 593094 208350
rect 593162 208294 593218 208350
rect 593286 208294 593342 208350
rect 592914 208170 592970 208226
rect 593038 208170 593094 208226
rect 593162 208170 593218 208226
rect 593286 208170 593342 208226
rect 592914 208046 592970 208102
rect 593038 208046 593094 208102
rect 593162 208046 593218 208102
rect 593286 208046 593342 208102
rect 592914 207922 592970 207978
rect 593038 207922 593094 207978
rect 593162 207922 593218 207978
rect 593286 207922 593342 207978
rect 592914 190294 592970 190350
rect 593038 190294 593094 190350
rect 593162 190294 593218 190350
rect 593286 190294 593342 190350
rect 592914 190170 592970 190226
rect 593038 190170 593094 190226
rect 593162 190170 593218 190226
rect 593286 190170 593342 190226
rect 592914 190046 592970 190102
rect 593038 190046 593094 190102
rect 593162 190046 593218 190102
rect 593286 190046 593342 190102
rect 592914 189922 592970 189978
rect 593038 189922 593094 189978
rect 593162 189922 593218 189978
rect 593286 189922 593342 189978
rect 592914 172294 592970 172350
rect 593038 172294 593094 172350
rect 593162 172294 593218 172350
rect 593286 172294 593342 172350
rect 592914 172170 592970 172226
rect 593038 172170 593094 172226
rect 593162 172170 593218 172226
rect 593286 172170 593342 172226
rect 592914 172046 592970 172102
rect 593038 172046 593094 172102
rect 593162 172046 593218 172102
rect 593286 172046 593342 172102
rect 592914 171922 592970 171978
rect 593038 171922 593094 171978
rect 593162 171922 593218 171978
rect 593286 171922 593342 171978
rect 592914 154294 592970 154350
rect 593038 154294 593094 154350
rect 593162 154294 593218 154350
rect 593286 154294 593342 154350
rect 592914 154170 592970 154226
rect 593038 154170 593094 154226
rect 593162 154170 593218 154226
rect 593286 154170 593342 154226
rect 592914 154046 592970 154102
rect 593038 154046 593094 154102
rect 593162 154046 593218 154102
rect 593286 154046 593342 154102
rect 592914 153922 592970 153978
rect 593038 153922 593094 153978
rect 593162 153922 593218 153978
rect 593286 153922 593342 153978
rect 592914 136294 592970 136350
rect 593038 136294 593094 136350
rect 593162 136294 593218 136350
rect 593286 136294 593342 136350
rect 592914 136170 592970 136226
rect 593038 136170 593094 136226
rect 593162 136170 593218 136226
rect 593286 136170 593342 136226
rect 592914 136046 592970 136102
rect 593038 136046 593094 136102
rect 593162 136046 593218 136102
rect 593286 136046 593342 136102
rect 592914 135922 592970 135978
rect 593038 135922 593094 135978
rect 593162 135922 593218 135978
rect 593286 135922 593342 135978
rect 592914 118294 592970 118350
rect 593038 118294 593094 118350
rect 593162 118294 593218 118350
rect 593286 118294 593342 118350
rect 592914 118170 592970 118226
rect 593038 118170 593094 118226
rect 593162 118170 593218 118226
rect 593286 118170 593342 118226
rect 592914 118046 592970 118102
rect 593038 118046 593094 118102
rect 593162 118046 593218 118102
rect 593286 118046 593342 118102
rect 592914 117922 592970 117978
rect 593038 117922 593094 117978
rect 593162 117922 593218 117978
rect 593286 117922 593342 117978
rect 592914 100294 592970 100350
rect 593038 100294 593094 100350
rect 593162 100294 593218 100350
rect 593286 100294 593342 100350
rect 592914 100170 592970 100226
rect 593038 100170 593094 100226
rect 593162 100170 593218 100226
rect 593286 100170 593342 100226
rect 592914 100046 592970 100102
rect 593038 100046 593094 100102
rect 593162 100046 593218 100102
rect 593286 100046 593342 100102
rect 592914 99922 592970 99978
rect 593038 99922 593094 99978
rect 593162 99922 593218 99978
rect 593286 99922 593342 99978
rect 592914 82294 592970 82350
rect 593038 82294 593094 82350
rect 593162 82294 593218 82350
rect 593286 82294 593342 82350
rect 592914 82170 592970 82226
rect 593038 82170 593094 82226
rect 593162 82170 593218 82226
rect 593286 82170 593342 82226
rect 592914 82046 592970 82102
rect 593038 82046 593094 82102
rect 593162 82046 593218 82102
rect 593286 82046 593342 82102
rect 592914 81922 592970 81978
rect 593038 81922 593094 81978
rect 593162 81922 593218 81978
rect 593286 81922 593342 81978
rect 589194 58294 589250 58350
rect 589318 58294 589374 58350
rect 589442 58294 589498 58350
rect 589566 58294 589622 58350
rect 589194 58170 589250 58226
rect 589318 58170 589374 58226
rect 589442 58170 589498 58226
rect 589566 58170 589622 58226
rect 589194 58046 589250 58102
rect 589318 58046 589374 58102
rect 589442 58046 589498 58102
rect 589566 58046 589622 58102
rect 589194 57922 589250 57978
rect 589318 57922 589374 57978
rect 589442 57922 589498 57978
rect 589566 57922 589622 57978
rect 589194 40294 589250 40350
rect 589318 40294 589374 40350
rect 589442 40294 589498 40350
rect 589566 40294 589622 40350
rect 589194 40170 589250 40226
rect 589318 40170 589374 40226
rect 589442 40170 589498 40226
rect 589566 40170 589622 40226
rect 589194 40046 589250 40102
rect 589318 40046 589374 40102
rect 589442 40046 589498 40102
rect 589566 40046 589622 40102
rect 589194 39922 589250 39978
rect 589318 39922 589374 39978
rect 589442 39922 589498 39978
rect 589566 39922 589622 39978
rect 589194 22294 589250 22350
rect 589318 22294 589374 22350
rect 589442 22294 589498 22350
rect 589566 22294 589622 22350
rect 589194 22170 589250 22226
rect 589318 22170 589374 22226
rect 589442 22170 589498 22226
rect 589566 22170 589622 22226
rect 589194 22046 589250 22102
rect 589318 22046 589374 22102
rect 589442 22046 589498 22102
rect 589566 22046 589622 22102
rect 589194 21922 589250 21978
rect 589318 21922 589374 21978
rect 589442 21922 589498 21978
rect 589566 21922 589622 21978
rect 589194 4294 589250 4350
rect 589318 4294 589374 4350
rect 589442 4294 589498 4350
rect 589566 4294 589622 4350
rect 589194 4170 589250 4226
rect 589318 4170 589374 4226
rect 589442 4170 589498 4226
rect 589566 4170 589622 4226
rect 562194 -1176 562250 -1120
rect 562318 -1176 562374 -1120
rect 562442 -1176 562498 -1120
rect 562566 -1176 562622 -1120
rect 562194 -1300 562250 -1244
rect 562318 -1300 562374 -1244
rect 562442 -1300 562498 -1244
rect 562566 -1300 562622 -1244
rect 562194 -1424 562250 -1368
rect 562318 -1424 562374 -1368
rect 562442 -1424 562498 -1368
rect 562566 -1424 562622 -1368
rect 562194 -1548 562250 -1492
rect 562318 -1548 562374 -1492
rect 562442 -1548 562498 -1492
rect 562566 -1548 562622 -1492
rect 589194 4046 589250 4102
rect 589318 4046 589374 4102
rect 589442 4046 589498 4102
rect 589566 4046 589622 4102
rect 589194 3922 589250 3978
rect 589318 3922 589374 3978
rect 589442 3922 589498 3978
rect 589566 3922 589622 3978
rect 589194 -216 589250 -160
rect 589318 -216 589374 -160
rect 589442 -216 589498 -160
rect 589566 -216 589622 -160
rect 589194 -340 589250 -284
rect 589318 -340 589374 -284
rect 589442 -340 589498 -284
rect 589566 -340 589622 -284
rect 589194 -464 589250 -408
rect 589318 -464 589374 -408
rect 589442 -464 589498 -408
rect 589566 -464 589622 -408
rect 589194 -588 589250 -532
rect 589318 -588 589374 -532
rect 589442 -588 589498 -532
rect 589566 -588 589622 -532
rect 592914 64294 592970 64350
rect 593038 64294 593094 64350
rect 593162 64294 593218 64350
rect 593286 64294 593342 64350
rect 592914 64170 592970 64226
rect 593038 64170 593094 64226
rect 593162 64170 593218 64226
rect 593286 64170 593342 64226
rect 592914 64046 592970 64102
rect 593038 64046 593094 64102
rect 593162 64046 593218 64102
rect 593286 64046 593342 64102
rect 592914 63922 592970 63978
rect 593038 63922 593094 63978
rect 593162 63922 593218 63978
rect 593286 63922 593342 63978
rect 592914 46294 592970 46350
rect 593038 46294 593094 46350
rect 593162 46294 593218 46350
rect 593286 46294 593342 46350
rect 592914 46170 592970 46226
rect 593038 46170 593094 46226
rect 593162 46170 593218 46226
rect 593286 46170 593342 46226
rect 592914 46046 592970 46102
rect 593038 46046 593094 46102
rect 593162 46046 593218 46102
rect 593286 46046 593342 46102
rect 592914 45922 592970 45978
rect 593038 45922 593094 45978
rect 593162 45922 593218 45978
rect 593286 45922 593342 45978
rect 592914 28294 592970 28350
rect 593038 28294 593094 28350
rect 593162 28294 593218 28350
rect 593286 28294 593342 28350
rect 592914 28170 592970 28226
rect 593038 28170 593094 28226
rect 593162 28170 593218 28226
rect 593286 28170 593342 28226
rect 592914 28046 592970 28102
rect 593038 28046 593094 28102
rect 593162 28046 593218 28102
rect 593286 28046 593342 28102
rect 592914 27922 592970 27978
rect 593038 27922 593094 27978
rect 593162 27922 593218 27978
rect 593286 27922 593342 27978
rect 592914 10294 592970 10350
rect 593038 10294 593094 10350
rect 593162 10294 593218 10350
rect 593286 10294 593342 10350
rect 592914 10170 592970 10226
rect 593038 10170 593094 10226
rect 593162 10170 593218 10226
rect 593286 10170 593342 10226
rect 592914 10046 592970 10102
rect 593038 10046 593094 10102
rect 593162 10046 593218 10102
rect 593286 10046 593342 10102
rect 592914 9922 592970 9978
rect 593038 9922 593094 9978
rect 593162 9922 593218 9978
rect 593286 9922 593342 9978
rect 596496 597156 596552 597212
rect 596620 597156 596676 597212
rect 596744 597156 596800 597212
rect 596868 597156 596924 597212
rect 596496 597032 596552 597088
rect 596620 597032 596676 597088
rect 596744 597032 596800 597088
rect 596868 597032 596924 597088
rect 596496 596908 596552 596964
rect 596620 596908 596676 596964
rect 596744 596908 596800 596964
rect 596868 596908 596924 596964
rect 596496 596784 596552 596840
rect 596620 596784 596676 596840
rect 596744 596784 596800 596840
rect 596868 596784 596924 596840
rect 596496 580294 596552 580350
rect 596620 580294 596676 580350
rect 596744 580294 596800 580350
rect 596868 580294 596924 580350
rect 596496 580170 596552 580226
rect 596620 580170 596676 580226
rect 596744 580170 596800 580226
rect 596868 580170 596924 580226
rect 596496 580046 596552 580102
rect 596620 580046 596676 580102
rect 596744 580046 596800 580102
rect 596868 580046 596924 580102
rect 596496 579922 596552 579978
rect 596620 579922 596676 579978
rect 596744 579922 596800 579978
rect 596868 579922 596924 579978
rect 596496 562294 596552 562350
rect 596620 562294 596676 562350
rect 596744 562294 596800 562350
rect 596868 562294 596924 562350
rect 596496 562170 596552 562226
rect 596620 562170 596676 562226
rect 596744 562170 596800 562226
rect 596868 562170 596924 562226
rect 596496 562046 596552 562102
rect 596620 562046 596676 562102
rect 596744 562046 596800 562102
rect 596868 562046 596924 562102
rect 596496 561922 596552 561978
rect 596620 561922 596676 561978
rect 596744 561922 596800 561978
rect 596868 561922 596924 561978
rect 596496 544294 596552 544350
rect 596620 544294 596676 544350
rect 596744 544294 596800 544350
rect 596868 544294 596924 544350
rect 596496 544170 596552 544226
rect 596620 544170 596676 544226
rect 596744 544170 596800 544226
rect 596868 544170 596924 544226
rect 596496 544046 596552 544102
rect 596620 544046 596676 544102
rect 596744 544046 596800 544102
rect 596868 544046 596924 544102
rect 596496 543922 596552 543978
rect 596620 543922 596676 543978
rect 596744 543922 596800 543978
rect 596868 543922 596924 543978
rect 596496 526294 596552 526350
rect 596620 526294 596676 526350
rect 596744 526294 596800 526350
rect 596868 526294 596924 526350
rect 596496 526170 596552 526226
rect 596620 526170 596676 526226
rect 596744 526170 596800 526226
rect 596868 526170 596924 526226
rect 596496 526046 596552 526102
rect 596620 526046 596676 526102
rect 596744 526046 596800 526102
rect 596868 526046 596924 526102
rect 596496 525922 596552 525978
rect 596620 525922 596676 525978
rect 596744 525922 596800 525978
rect 596868 525922 596924 525978
rect 596496 508294 596552 508350
rect 596620 508294 596676 508350
rect 596744 508294 596800 508350
rect 596868 508294 596924 508350
rect 596496 508170 596552 508226
rect 596620 508170 596676 508226
rect 596744 508170 596800 508226
rect 596868 508170 596924 508226
rect 596496 508046 596552 508102
rect 596620 508046 596676 508102
rect 596744 508046 596800 508102
rect 596868 508046 596924 508102
rect 596496 507922 596552 507978
rect 596620 507922 596676 507978
rect 596744 507922 596800 507978
rect 596868 507922 596924 507978
rect 596496 490294 596552 490350
rect 596620 490294 596676 490350
rect 596744 490294 596800 490350
rect 596868 490294 596924 490350
rect 596496 490170 596552 490226
rect 596620 490170 596676 490226
rect 596744 490170 596800 490226
rect 596868 490170 596924 490226
rect 596496 490046 596552 490102
rect 596620 490046 596676 490102
rect 596744 490046 596800 490102
rect 596868 490046 596924 490102
rect 596496 489922 596552 489978
rect 596620 489922 596676 489978
rect 596744 489922 596800 489978
rect 596868 489922 596924 489978
rect 596496 472294 596552 472350
rect 596620 472294 596676 472350
rect 596744 472294 596800 472350
rect 596868 472294 596924 472350
rect 596496 472170 596552 472226
rect 596620 472170 596676 472226
rect 596744 472170 596800 472226
rect 596868 472170 596924 472226
rect 596496 472046 596552 472102
rect 596620 472046 596676 472102
rect 596744 472046 596800 472102
rect 596868 472046 596924 472102
rect 596496 471922 596552 471978
rect 596620 471922 596676 471978
rect 596744 471922 596800 471978
rect 596868 471922 596924 471978
rect 596496 454294 596552 454350
rect 596620 454294 596676 454350
rect 596744 454294 596800 454350
rect 596868 454294 596924 454350
rect 596496 454170 596552 454226
rect 596620 454170 596676 454226
rect 596744 454170 596800 454226
rect 596868 454170 596924 454226
rect 596496 454046 596552 454102
rect 596620 454046 596676 454102
rect 596744 454046 596800 454102
rect 596868 454046 596924 454102
rect 596496 453922 596552 453978
rect 596620 453922 596676 453978
rect 596744 453922 596800 453978
rect 596868 453922 596924 453978
rect 596496 436294 596552 436350
rect 596620 436294 596676 436350
rect 596744 436294 596800 436350
rect 596868 436294 596924 436350
rect 596496 436170 596552 436226
rect 596620 436170 596676 436226
rect 596744 436170 596800 436226
rect 596868 436170 596924 436226
rect 596496 436046 596552 436102
rect 596620 436046 596676 436102
rect 596744 436046 596800 436102
rect 596868 436046 596924 436102
rect 596496 435922 596552 435978
rect 596620 435922 596676 435978
rect 596744 435922 596800 435978
rect 596868 435922 596924 435978
rect 596496 418294 596552 418350
rect 596620 418294 596676 418350
rect 596744 418294 596800 418350
rect 596868 418294 596924 418350
rect 596496 418170 596552 418226
rect 596620 418170 596676 418226
rect 596744 418170 596800 418226
rect 596868 418170 596924 418226
rect 596496 418046 596552 418102
rect 596620 418046 596676 418102
rect 596744 418046 596800 418102
rect 596868 418046 596924 418102
rect 596496 417922 596552 417978
rect 596620 417922 596676 417978
rect 596744 417922 596800 417978
rect 596868 417922 596924 417978
rect 596496 400294 596552 400350
rect 596620 400294 596676 400350
rect 596744 400294 596800 400350
rect 596868 400294 596924 400350
rect 596496 400170 596552 400226
rect 596620 400170 596676 400226
rect 596744 400170 596800 400226
rect 596868 400170 596924 400226
rect 596496 400046 596552 400102
rect 596620 400046 596676 400102
rect 596744 400046 596800 400102
rect 596868 400046 596924 400102
rect 596496 399922 596552 399978
rect 596620 399922 596676 399978
rect 596744 399922 596800 399978
rect 596868 399922 596924 399978
rect 596496 382294 596552 382350
rect 596620 382294 596676 382350
rect 596744 382294 596800 382350
rect 596868 382294 596924 382350
rect 596496 382170 596552 382226
rect 596620 382170 596676 382226
rect 596744 382170 596800 382226
rect 596868 382170 596924 382226
rect 596496 382046 596552 382102
rect 596620 382046 596676 382102
rect 596744 382046 596800 382102
rect 596868 382046 596924 382102
rect 596496 381922 596552 381978
rect 596620 381922 596676 381978
rect 596744 381922 596800 381978
rect 596868 381922 596924 381978
rect 596496 364294 596552 364350
rect 596620 364294 596676 364350
rect 596744 364294 596800 364350
rect 596868 364294 596924 364350
rect 596496 364170 596552 364226
rect 596620 364170 596676 364226
rect 596744 364170 596800 364226
rect 596868 364170 596924 364226
rect 596496 364046 596552 364102
rect 596620 364046 596676 364102
rect 596744 364046 596800 364102
rect 596868 364046 596924 364102
rect 596496 363922 596552 363978
rect 596620 363922 596676 363978
rect 596744 363922 596800 363978
rect 596868 363922 596924 363978
rect 596496 346294 596552 346350
rect 596620 346294 596676 346350
rect 596744 346294 596800 346350
rect 596868 346294 596924 346350
rect 596496 346170 596552 346226
rect 596620 346170 596676 346226
rect 596744 346170 596800 346226
rect 596868 346170 596924 346226
rect 596496 346046 596552 346102
rect 596620 346046 596676 346102
rect 596744 346046 596800 346102
rect 596868 346046 596924 346102
rect 596496 345922 596552 345978
rect 596620 345922 596676 345978
rect 596744 345922 596800 345978
rect 596868 345922 596924 345978
rect 596496 328294 596552 328350
rect 596620 328294 596676 328350
rect 596744 328294 596800 328350
rect 596868 328294 596924 328350
rect 596496 328170 596552 328226
rect 596620 328170 596676 328226
rect 596744 328170 596800 328226
rect 596868 328170 596924 328226
rect 596496 328046 596552 328102
rect 596620 328046 596676 328102
rect 596744 328046 596800 328102
rect 596868 328046 596924 328102
rect 596496 327922 596552 327978
rect 596620 327922 596676 327978
rect 596744 327922 596800 327978
rect 596868 327922 596924 327978
rect 596496 310294 596552 310350
rect 596620 310294 596676 310350
rect 596744 310294 596800 310350
rect 596868 310294 596924 310350
rect 596496 310170 596552 310226
rect 596620 310170 596676 310226
rect 596744 310170 596800 310226
rect 596868 310170 596924 310226
rect 596496 310046 596552 310102
rect 596620 310046 596676 310102
rect 596744 310046 596800 310102
rect 596868 310046 596924 310102
rect 596496 309922 596552 309978
rect 596620 309922 596676 309978
rect 596744 309922 596800 309978
rect 596868 309922 596924 309978
rect 596496 292294 596552 292350
rect 596620 292294 596676 292350
rect 596744 292294 596800 292350
rect 596868 292294 596924 292350
rect 596496 292170 596552 292226
rect 596620 292170 596676 292226
rect 596744 292170 596800 292226
rect 596868 292170 596924 292226
rect 596496 292046 596552 292102
rect 596620 292046 596676 292102
rect 596744 292046 596800 292102
rect 596868 292046 596924 292102
rect 596496 291922 596552 291978
rect 596620 291922 596676 291978
rect 596744 291922 596800 291978
rect 596868 291922 596924 291978
rect 596496 274294 596552 274350
rect 596620 274294 596676 274350
rect 596744 274294 596800 274350
rect 596868 274294 596924 274350
rect 596496 274170 596552 274226
rect 596620 274170 596676 274226
rect 596744 274170 596800 274226
rect 596868 274170 596924 274226
rect 596496 274046 596552 274102
rect 596620 274046 596676 274102
rect 596744 274046 596800 274102
rect 596868 274046 596924 274102
rect 596496 273922 596552 273978
rect 596620 273922 596676 273978
rect 596744 273922 596800 273978
rect 596868 273922 596924 273978
rect 596496 256294 596552 256350
rect 596620 256294 596676 256350
rect 596744 256294 596800 256350
rect 596868 256294 596924 256350
rect 596496 256170 596552 256226
rect 596620 256170 596676 256226
rect 596744 256170 596800 256226
rect 596868 256170 596924 256226
rect 596496 256046 596552 256102
rect 596620 256046 596676 256102
rect 596744 256046 596800 256102
rect 596868 256046 596924 256102
rect 596496 255922 596552 255978
rect 596620 255922 596676 255978
rect 596744 255922 596800 255978
rect 596868 255922 596924 255978
rect 596496 238294 596552 238350
rect 596620 238294 596676 238350
rect 596744 238294 596800 238350
rect 596868 238294 596924 238350
rect 596496 238170 596552 238226
rect 596620 238170 596676 238226
rect 596744 238170 596800 238226
rect 596868 238170 596924 238226
rect 596496 238046 596552 238102
rect 596620 238046 596676 238102
rect 596744 238046 596800 238102
rect 596868 238046 596924 238102
rect 596496 237922 596552 237978
rect 596620 237922 596676 237978
rect 596744 237922 596800 237978
rect 596868 237922 596924 237978
rect 596496 220294 596552 220350
rect 596620 220294 596676 220350
rect 596744 220294 596800 220350
rect 596868 220294 596924 220350
rect 596496 220170 596552 220226
rect 596620 220170 596676 220226
rect 596744 220170 596800 220226
rect 596868 220170 596924 220226
rect 596496 220046 596552 220102
rect 596620 220046 596676 220102
rect 596744 220046 596800 220102
rect 596868 220046 596924 220102
rect 596496 219922 596552 219978
rect 596620 219922 596676 219978
rect 596744 219922 596800 219978
rect 596868 219922 596924 219978
rect 596496 202294 596552 202350
rect 596620 202294 596676 202350
rect 596744 202294 596800 202350
rect 596868 202294 596924 202350
rect 596496 202170 596552 202226
rect 596620 202170 596676 202226
rect 596744 202170 596800 202226
rect 596868 202170 596924 202226
rect 596496 202046 596552 202102
rect 596620 202046 596676 202102
rect 596744 202046 596800 202102
rect 596868 202046 596924 202102
rect 596496 201922 596552 201978
rect 596620 201922 596676 201978
rect 596744 201922 596800 201978
rect 596868 201922 596924 201978
rect 596496 184294 596552 184350
rect 596620 184294 596676 184350
rect 596744 184294 596800 184350
rect 596868 184294 596924 184350
rect 596496 184170 596552 184226
rect 596620 184170 596676 184226
rect 596744 184170 596800 184226
rect 596868 184170 596924 184226
rect 596496 184046 596552 184102
rect 596620 184046 596676 184102
rect 596744 184046 596800 184102
rect 596868 184046 596924 184102
rect 596496 183922 596552 183978
rect 596620 183922 596676 183978
rect 596744 183922 596800 183978
rect 596868 183922 596924 183978
rect 596496 166294 596552 166350
rect 596620 166294 596676 166350
rect 596744 166294 596800 166350
rect 596868 166294 596924 166350
rect 596496 166170 596552 166226
rect 596620 166170 596676 166226
rect 596744 166170 596800 166226
rect 596868 166170 596924 166226
rect 596496 166046 596552 166102
rect 596620 166046 596676 166102
rect 596744 166046 596800 166102
rect 596868 166046 596924 166102
rect 596496 165922 596552 165978
rect 596620 165922 596676 165978
rect 596744 165922 596800 165978
rect 596868 165922 596924 165978
rect 596496 148294 596552 148350
rect 596620 148294 596676 148350
rect 596744 148294 596800 148350
rect 596868 148294 596924 148350
rect 596496 148170 596552 148226
rect 596620 148170 596676 148226
rect 596744 148170 596800 148226
rect 596868 148170 596924 148226
rect 596496 148046 596552 148102
rect 596620 148046 596676 148102
rect 596744 148046 596800 148102
rect 596868 148046 596924 148102
rect 596496 147922 596552 147978
rect 596620 147922 596676 147978
rect 596744 147922 596800 147978
rect 596868 147922 596924 147978
rect 596496 130294 596552 130350
rect 596620 130294 596676 130350
rect 596744 130294 596800 130350
rect 596868 130294 596924 130350
rect 596496 130170 596552 130226
rect 596620 130170 596676 130226
rect 596744 130170 596800 130226
rect 596868 130170 596924 130226
rect 596496 130046 596552 130102
rect 596620 130046 596676 130102
rect 596744 130046 596800 130102
rect 596868 130046 596924 130102
rect 596496 129922 596552 129978
rect 596620 129922 596676 129978
rect 596744 129922 596800 129978
rect 596868 129922 596924 129978
rect 596496 112294 596552 112350
rect 596620 112294 596676 112350
rect 596744 112294 596800 112350
rect 596868 112294 596924 112350
rect 596496 112170 596552 112226
rect 596620 112170 596676 112226
rect 596744 112170 596800 112226
rect 596868 112170 596924 112226
rect 596496 112046 596552 112102
rect 596620 112046 596676 112102
rect 596744 112046 596800 112102
rect 596868 112046 596924 112102
rect 596496 111922 596552 111978
rect 596620 111922 596676 111978
rect 596744 111922 596800 111978
rect 596868 111922 596924 111978
rect 596496 94294 596552 94350
rect 596620 94294 596676 94350
rect 596744 94294 596800 94350
rect 596868 94294 596924 94350
rect 596496 94170 596552 94226
rect 596620 94170 596676 94226
rect 596744 94170 596800 94226
rect 596868 94170 596924 94226
rect 596496 94046 596552 94102
rect 596620 94046 596676 94102
rect 596744 94046 596800 94102
rect 596868 94046 596924 94102
rect 596496 93922 596552 93978
rect 596620 93922 596676 93978
rect 596744 93922 596800 93978
rect 596868 93922 596924 93978
rect 596496 76294 596552 76350
rect 596620 76294 596676 76350
rect 596744 76294 596800 76350
rect 596868 76294 596924 76350
rect 596496 76170 596552 76226
rect 596620 76170 596676 76226
rect 596744 76170 596800 76226
rect 596868 76170 596924 76226
rect 596496 76046 596552 76102
rect 596620 76046 596676 76102
rect 596744 76046 596800 76102
rect 596868 76046 596924 76102
rect 596496 75922 596552 75978
rect 596620 75922 596676 75978
rect 596744 75922 596800 75978
rect 596868 75922 596924 75978
rect 596496 58294 596552 58350
rect 596620 58294 596676 58350
rect 596744 58294 596800 58350
rect 596868 58294 596924 58350
rect 596496 58170 596552 58226
rect 596620 58170 596676 58226
rect 596744 58170 596800 58226
rect 596868 58170 596924 58226
rect 596496 58046 596552 58102
rect 596620 58046 596676 58102
rect 596744 58046 596800 58102
rect 596868 58046 596924 58102
rect 596496 57922 596552 57978
rect 596620 57922 596676 57978
rect 596744 57922 596800 57978
rect 596868 57922 596924 57978
rect 596496 40294 596552 40350
rect 596620 40294 596676 40350
rect 596744 40294 596800 40350
rect 596868 40294 596924 40350
rect 596496 40170 596552 40226
rect 596620 40170 596676 40226
rect 596744 40170 596800 40226
rect 596868 40170 596924 40226
rect 596496 40046 596552 40102
rect 596620 40046 596676 40102
rect 596744 40046 596800 40102
rect 596868 40046 596924 40102
rect 596496 39922 596552 39978
rect 596620 39922 596676 39978
rect 596744 39922 596800 39978
rect 596868 39922 596924 39978
rect 596496 22294 596552 22350
rect 596620 22294 596676 22350
rect 596744 22294 596800 22350
rect 596868 22294 596924 22350
rect 596496 22170 596552 22226
rect 596620 22170 596676 22226
rect 596744 22170 596800 22226
rect 596868 22170 596924 22226
rect 596496 22046 596552 22102
rect 596620 22046 596676 22102
rect 596744 22046 596800 22102
rect 596868 22046 596924 22102
rect 596496 21922 596552 21978
rect 596620 21922 596676 21978
rect 596744 21922 596800 21978
rect 596868 21922 596924 21978
rect 596496 4294 596552 4350
rect 596620 4294 596676 4350
rect 596744 4294 596800 4350
rect 596868 4294 596924 4350
rect 596496 4170 596552 4226
rect 596620 4170 596676 4226
rect 596744 4170 596800 4226
rect 596868 4170 596924 4226
rect 596496 4046 596552 4102
rect 596620 4046 596676 4102
rect 596744 4046 596800 4102
rect 596868 4046 596924 4102
rect 596496 3922 596552 3978
rect 596620 3922 596676 3978
rect 596744 3922 596800 3978
rect 596868 3922 596924 3978
rect 596496 -216 596552 -160
rect 596620 -216 596676 -160
rect 596744 -216 596800 -160
rect 596868 -216 596924 -160
rect 596496 -340 596552 -284
rect 596620 -340 596676 -284
rect 596744 -340 596800 -284
rect 596868 -340 596924 -284
rect 596496 -464 596552 -408
rect 596620 -464 596676 -408
rect 596744 -464 596800 -408
rect 596868 -464 596924 -408
rect 596496 -588 596552 -532
rect 596620 -588 596676 -532
rect 596744 -588 596800 -532
rect 596868 -588 596924 -532
rect 597456 586294 597512 586350
rect 597580 586294 597636 586350
rect 597704 586294 597760 586350
rect 597828 586294 597884 586350
rect 597456 586170 597512 586226
rect 597580 586170 597636 586226
rect 597704 586170 597760 586226
rect 597828 586170 597884 586226
rect 597456 586046 597512 586102
rect 597580 586046 597636 586102
rect 597704 586046 597760 586102
rect 597828 586046 597884 586102
rect 597456 585922 597512 585978
rect 597580 585922 597636 585978
rect 597704 585922 597760 585978
rect 597828 585922 597884 585978
rect 597456 568294 597512 568350
rect 597580 568294 597636 568350
rect 597704 568294 597760 568350
rect 597828 568294 597884 568350
rect 597456 568170 597512 568226
rect 597580 568170 597636 568226
rect 597704 568170 597760 568226
rect 597828 568170 597884 568226
rect 597456 568046 597512 568102
rect 597580 568046 597636 568102
rect 597704 568046 597760 568102
rect 597828 568046 597884 568102
rect 597456 567922 597512 567978
rect 597580 567922 597636 567978
rect 597704 567922 597760 567978
rect 597828 567922 597884 567978
rect 597456 550294 597512 550350
rect 597580 550294 597636 550350
rect 597704 550294 597760 550350
rect 597828 550294 597884 550350
rect 597456 550170 597512 550226
rect 597580 550170 597636 550226
rect 597704 550170 597760 550226
rect 597828 550170 597884 550226
rect 597456 550046 597512 550102
rect 597580 550046 597636 550102
rect 597704 550046 597760 550102
rect 597828 550046 597884 550102
rect 597456 549922 597512 549978
rect 597580 549922 597636 549978
rect 597704 549922 597760 549978
rect 597828 549922 597884 549978
rect 597456 532294 597512 532350
rect 597580 532294 597636 532350
rect 597704 532294 597760 532350
rect 597828 532294 597884 532350
rect 597456 532170 597512 532226
rect 597580 532170 597636 532226
rect 597704 532170 597760 532226
rect 597828 532170 597884 532226
rect 597456 532046 597512 532102
rect 597580 532046 597636 532102
rect 597704 532046 597760 532102
rect 597828 532046 597884 532102
rect 597456 531922 597512 531978
rect 597580 531922 597636 531978
rect 597704 531922 597760 531978
rect 597828 531922 597884 531978
rect 597456 514294 597512 514350
rect 597580 514294 597636 514350
rect 597704 514294 597760 514350
rect 597828 514294 597884 514350
rect 597456 514170 597512 514226
rect 597580 514170 597636 514226
rect 597704 514170 597760 514226
rect 597828 514170 597884 514226
rect 597456 514046 597512 514102
rect 597580 514046 597636 514102
rect 597704 514046 597760 514102
rect 597828 514046 597884 514102
rect 597456 513922 597512 513978
rect 597580 513922 597636 513978
rect 597704 513922 597760 513978
rect 597828 513922 597884 513978
rect 597456 496294 597512 496350
rect 597580 496294 597636 496350
rect 597704 496294 597760 496350
rect 597828 496294 597884 496350
rect 597456 496170 597512 496226
rect 597580 496170 597636 496226
rect 597704 496170 597760 496226
rect 597828 496170 597884 496226
rect 597456 496046 597512 496102
rect 597580 496046 597636 496102
rect 597704 496046 597760 496102
rect 597828 496046 597884 496102
rect 597456 495922 597512 495978
rect 597580 495922 597636 495978
rect 597704 495922 597760 495978
rect 597828 495922 597884 495978
rect 597456 478294 597512 478350
rect 597580 478294 597636 478350
rect 597704 478294 597760 478350
rect 597828 478294 597884 478350
rect 597456 478170 597512 478226
rect 597580 478170 597636 478226
rect 597704 478170 597760 478226
rect 597828 478170 597884 478226
rect 597456 478046 597512 478102
rect 597580 478046 597636 478102
rect 597704 478046 597760 478102
rect 597828 478046 597884 478102
rect 597456 477922 597512 477978
rect 597580 477922 597636 477978
rect 597704 477922 597760 477978
rect 597828 477922 597884 477978
rect 597456 460294 597512 460350
rect 597580 460294 597636 460350
rect 597704 460294 597760 460350
rect 597828 460294 597884 460350
rect 597456 460170 597512 460226
rect 597580 460170 597636 460226
rect 597704 460170 597760 460226
rect 597828 460170 597884 460226
rect 597456 460046 597512 460102
rect 597580 460046 597636 460102
rect 597704 460046 597760 460102
rect 597828 460046 597884 460102
rect 597456 459922 597512 459978
rect 597580 459922 597636 459978
rect 597704 459922 597760 459978
rect 597828 459922 597884 459978
rect 597456 442294 597512 442350
rect 597580 442294 597636 442350
rect 597704 442294 597760 442350
rect 597828 442294 597884 442350
rect 597456 442170 597512 442226
rect 597580 442170 597636 442226
rect 597704 442170 597760 442226
rect 597828 442170 597884 442226
rect 597456 442046 597512 442102
rect 597580 442046 597636 442102
rect 597704 442046 597760 442102
rect 597828 442046 597884 442102
rect 597456 441922 597512 441978
rect 597580 441922 597636 441978
rect 597704 441922 597760 441978
rect 597828 441922 597884 441978
rect 597456 424294 597512 424350
rect 597580 424294 597636 424350
rect 597704 424294 597760 424350
rect 597828 424294 597884 424350
rect 597456 424170 597512 424226
rect 597580 424170 597636 424226
rect 597704 424170 597760 424226
rect 597828 424170 597884 424226
rect 597456 424046 597512 424102
rect 597580 424046 597636 424102
rect 597704 424046 597760 424102
rect 597828 424046 597884 424102
rect 597456 423922 597512 423978
rect 597580 423922 597636 423978
rect 597704 423922 597760 423978
rect 597828 423922 597884 423978
rect 597456 406294 597512 406350
rect 597580 406294 597636 406350
rect 597704 406294 597760 406350
rect 597828 406294 597884 406350
rect 597456 406170 597512 406226
rect 597580 406170 597636 406226
rect 597704 406170 597760 406226
rect 597828 406170 597884 406226
rect 597456 406046 597512 406102
rect 597580 406046 597636 406102
rect 597704 406046 597760 406102
rect 597828 406046 597884 406102
rect 597456 405922 597512 405978
rect 597580 405922 597636 405978
rect 597704 405922 597760 405978
rect 597828 405922 597884 405978
rect 597456 388294 597512 388350
rect 597580 388294 597636 388350
rect 597704 388294 597760 388350
rect 597828 388294 597884 388350
rect 597456 388170 597512 388226
rect 597580 388170 597636 388226
rect 597704 388170 597760 388226
rect 597828 388170 597884 388226
rect 597456 388046 597512 388102
rect 597580 388046 597636 388102
rect 597704 388046 597760 388102
rect 597828 388046 597884 388102
rect 597456 387922 597512 387978
rect 597580 387922 597636 387978
rect 597704 387922 597760 387978
rect 597828 387922 597884 387978
rect 597456 370294 597512 370350
rect 597580 370294 597636 370350
rect 597704 370294 597760 370350
rect 597828 370294 597884 370350
rect 597456 370170 597512 370226
rect 597580 370170 597636 370226
rect 597704 370170 597760 370226
rect 597828 370170 597884 370226
rect 597456 370046 597512 370102
rect 597580 370046 597636 370102
rect 597704 370046 597760 370102
rect 597828 370046 597884 370102
rect 597456 369922 597512 369978
rect 597580 369922 597636 369978
rect 597704 369922 597760 369978
rect 597828 369922 597884 369978
rect 597456 352294 597512 352350
rect 597580 352294 597636 352350
rect 597704 352294 597760 352350
rect 597828 352294 597884 352350
rect 597456 352170 597512 352226
rect 597580 352170 597636 352226
rect 597704 352170 597760 352226
rect 597828 352170 597884 352226
rect 597456 352046 597512 352102
rect 597580 352046 597636 352102
rect 597704 352046 597760 352102
rect 597828 352046 597884 352102
rect 597456 351922 597512 351978
rect 597580 351922 597636 351978
rect 597704 351922 597760 351978
rect 597828 351922 597884 351978
rect 597456 334294 597512 334350
rect 597580 334294 597636 334350
rect 597704 334294 597760 334350
rect 597828 334294 597884 334350
rect 597456 334170 597512 334226
rect 597580 334170 597636 334226
rect 597704 334170 597760 334226
rect 597828 334170 597884 334226
rect 597456 334046 597512 334102
rect 597580 334046 597636 334102
rect 597704 334046 597760 334102
rect 597828 334046 597884 334102
rect 597456 333922 597512 333978
rect 597580 333922 597636 333978
rect 597704 333922 597760 333978
rect 597828 333922 597884 333978
rect 597456 316294 597512 316350
rect 597580 316294 597636 316350
rect 597704 316294 597760 316350
rect 597828 316294 597884 316350
rect 597456 316170 597512 316226
rect 597580 316170 597636 316226
rect 597704 316170 597760 316226
rect 597828 316170 597884 316226
rect 597456 316046 597512 316102
rect 597580 316046 597636 316102
rect 597704 316046 597760 316102
rect 597828 316046 597884 316102
rect 597456 315922 597512 315978
rect 597580 315922 597636 315978
rect 597704 315922 597760 315978
rect 597828 315922 597884 315978
rect 597456 298294 597512 298350
rect 597580 298294 597636 298350
rect 597704 298294 597760 298350
rect 597828 298294 597884 298350
rect 597456 298170 597512 298226
rect 597580 298170 597636 298226
rect 597704 298170 597760 298226
rect 597828 298170 597884 298226
rect 597456 298046 597512 298102
rect 597580 298046 597636 298102
rect 597704 298046 597760 298102
rect 597828 298046 597884 298102
rect 597456 297922 597512 297978
rect 597580 297922 597636 297978
rect 597704 297922 597760 297978
rect 597828 297922 597884 297978
rect 597456 280294 597512 280350
rect 597580 280294 597636 280350
rect 597704 280294 597760 280350
rect 597828 280294 597884 280350
rect 597456 280170 597512 280226
rect 597580 280170 597636 280226
rect 597704 280170 597760 280226
rect 597828 280170 597884 280226
rect 597456 280046 597512 280102
rect 597580 280046 597636 280102
rect 597704 280046 597760 280102
rect 597828 280046 597884 280102
rect 597456 279922 597512 279978
rect 597580 279922 597636 279978
rect 597704 279922 597760 279978
rect 597828 279922 597884 279978
rect 597456 262294 597512 262350
rect 597580 262294 597636 262350
rect 597704 262294 597760 262350
rect 597828 262294 597884 262350
rect 597456 262170 597512 262226
rect 597580 262170 597636 262226
rect 597704 262170 597760 262226
rect 597828 262170 597884 262226
rect 597456 262046 597512 262102
rect 597580 262046 597636 262102
rect 597704 262046 597760 262102
rect 597828 262046 597884 262102
rect 597456 261922 597512 261978
rect 597580 261922 597636 261978
rect 597704 261922 597760 261978
rect 597828 261922 597884 261978
rect 597456 244294 597512 244350
rect 597580 244294 597636 244350
rect 597704 244294 597760 244350
rect 597828 244294 597884 244350
rect 597456 244170 597512 244226
rect 597580 244170 597636 244226
rect 597704 244170 597760 244226
rect 597828 244170 597884 244226
rect 597456 244046 597512 244102
rect 597580 244046 597636 244102
rect 597704 244046 597760 244102
rect 597828 244046 597884 244102
rect 597456 243922 597512 243978
rect 597580 243922 597636 243978
rect 597704 243922 597760 243978
rect 597828 243922 597884 243978
rect 597456 226294 597512 226350
rect 597580 226294 597636 226350
rect 597704 226294 597760 226350
rect 597828 226294 597884 226350
rect 597456 226170 597512 226226
rect 597580 226170 597636 226226
rect 597704 226170 597760 226226
rect 597828 226170 597884 226226
rect 597456 226046 597512 226102
rect 597580 226046 597636 226102
rect 597704 226046 597760 226102
rect 597828 226046 597884 226102
rect 597456 225922 597512 225978
rect 597580 225922 597636 225978
rect 597704 225922 597760 225978
rect 597828 225922 597884 225978
rect 597456 208294 597512 208350
rect 597580 208294 597636 208350
rect 597704 208294 597760 208350
rect 597828 208294 597884 208350
rect 597456 208170 597512 208226
rect 597580 208170 597636 208226
rect 597704 208170 597760 208226
rect 597828 208170 597884 208226
rect 597456 208046 597512 208102
rect 597580 208046 597636 208102
rect 597704 208046 597760 208102
rect 597828 208046 597884 208102
rect 597456 207922 597512 207978
rect 597580 207922 597636 207978
rect 597704 207922 597760 207978
rect 597828 207922 597884 207978
rect 597456 190294 597512 190350
rect 597580 190294 597636 190350
rect 597704 190294 597760 190350
rect 597828 190294 597884 190350
rect 597456 190170 597512 190226
rect 597580 190170 597636 190226
rect 597704 190170 597760 190226
rect 597828 190170 597884 190226
rect 597456 190046 597512 190102
rect 597580 190046 597636 190102
rect 597704 190046 597760 190102
rect 597828 190046 597884 190102
rect 597456 189922 597512 189978
rect 597580 189922 597636 189978
rect 597704 189922 597760 189978
rect 597828 189922 597884 189978
rect 597456 172294 597512 172350
rect 597580 172294 597636 172350
rect 597704 172294 597760 172350
rect 597828 172294 597884 172350
rect 597456 172170 597512 172226
rect 597580 172170 597636 172226
rect 597704 172170 597760 172226
rect 597828 172170 597884 172226
rect 597456 172046 597512 172102
rect 597580 172046 597636 172102
rect 597704 172046 597760 172102
rect 597828 172046 597884 172102
rect 597456 171922 597512 171978
rect 597580 171922 597636 171978
rect 597704 171922 597760 171978
rect 597828 171922 597884 171978
rect 597456 154294 597512 154350
rect 597580 154294 597636 154350
rect 597704 154294 597760 154350
rect 597828 154294 597884 154350
rect 597456 154170 597512 154226
rect 597580 154170 597636 154226
rect 597704 154170 597760 154226
rect 597828 154170 597884 154226
rect 597456 154046 597512 154102
rect 597580 154046 597636 154102
rect 597704 154046 597760 154102
rect 597828 154046 597884 154102
rect 597456 153922 597512 153978
rect 597580 153922 597636 153978
rect 597704 153922 597760 153978
rect 597828 153922 597884 153978
rect 597456 136294 597512 136350
rect 597580 136294 597636 136350
rect 597704 136294 597760 136350
rect 597828 136294 597884 136350
rect 597456 136170 597512 136226
rect 597580 136170 597636 136226
rect 597704 136170 597760 136226
rect 597828 136170 597884 136226
rect 597456 136046 597512 136102
rect 597580 136046 597636 136102
rect 597704 136046 597760 136102
rect 597828 136046 597884 136102
rect 597456 135922 597512 135978
rect 597580 135922 597636 135978
rect 597704 135922 597760 135978
rect 597828 135922 597884 135978
rect 597456 118294 597512 118350
rect 597580 118294 597636 118350
rect 597704 118294 597760 118350
rect 597828 118294 597884 118350
rect 597456 118170 597512 118226
rect 597580 118170 597636 118226
rect 597704 118170 597760 118226
rect 597828 118170 597884 118226
rect 597456 118046 597512 118102
rect 597580 118046 597636 118102
rect 597704 118046 597760 118102
rect 597828 118046 597884 118102
rect 597456 117922 597512 117978
rect 597580 117922 597636 117978
rect 597704 117922 597760 117978
rect 597828 117922 597884 117978
rect 597456 100294 597512 100350
rect 597580 100294 597636 100350
rect 597704 100294 597760 100350
rect 597828 100294 597884 100350
rect 597456 100170 597512 100226
rect 597580 100170 597636 100226
rect 597704 100170 597760 100226
rect 597828 100170 597884 100226
rect 597456 100046 597512 100102
rect 597580 100046 597636 100102
rect 597704 100046 597760 100102
rect 597828 100046 597884 100102
rect 597456 99922 597512 99978
rect 597580 99922 597636 99978
rect 597704 99922 597760 99978
rect 597828 99922 597884 99978
rect 597456 82294 597512 82350
rect 597580 82294 597636 82350
rect 597704 82294 597760 82350
rect 597828 82294 597884 82350
rect 597456 82170 597512 82226
rect 597580 82170 597636 82226
rect 597704 82170 597760 82226
rect 597828 82170 597884 82226
rect 597456 82046 597512 82102
rect 597580 82046 597636 82102
rect 597704 82046 597760 82102
rect 597828 82046 597884 82102
rect 597456 81922 597512 81978
rect 597580 81922 597636 81978
rect 597704 81922 597760 81978
rect 597828 81922 597884 81978
rect 597456 64294 597512 64350
rect 597580 64294 597636 64350
rect 597704 64294 597760 64350
rect 597828 64294 597884 64350
rect 597456 64170 597512 64226
rect 597580 64170 597636 64226
rect 597704 64170 597760 64226
rect 597828 64170 597884 64226
rect 597456 64046 597512 64102
rect 597580 64046 597636 64102
rect 597704 64046 597760 64102
rect 597828 64046 597884 64102
rect 597456 63922 597512 63978
rect 597580 63922 597636 63978
rect 597704 63922 597760 63978
rect 597828 63922 597884 63978
rect 597456 46294 597512 46350
rect 597580 46294 597636 46350
rect 597704 46294 597760 46350
rect 597828 46294 597884 46350
rect 597456 46170 597512 46226
rect 597580 46170 597636 46226
rect 597704 46170 597760 46226
rect 597828 46170 597884 46226
rect 597456 46046 597512 46102
rect 597580 46046 597636 46102
rect 597704 46046 597760 46102
rect 597828 46046 597884 46102
rect 597456 45922 597512 45978
rect 597580 45922 597636 45978
rect 597704 45922 597760 45978
rect 597828 45922 597884 45978
rect 597456 28294 597512 28350
rect 597580 28294 597636 28350
rect 597704 28294 597760 28350
rect 597828 28294 597884 28350
rect 597456 28170 597512 28226
rect 597580 28170 597636 28226
rect 597704 28170 597760 28226
rect 597828 28170 597884 28226
rect 597456 28046 597512 28102
rect 597580 28046 597636 28102
rect 597704 28046 597760 28102
rect 597828 28046 597884 28102
rect 597456 27922 597512 27978
rect 597580 27922 597636 27978
rect 597704 27922 597760 27978
rect 597828 27922 597884 27978
rect 597456 10294 597512 10350
rect 597580 10294 597636 10350
rect 597704 10294 597760 10350
rect 597828 10294 597884 10350
rect 597456 10170 597512 10226
rect 597580 10170 597636 10226
rect 597704 10170 597760 10226
rect 597828 10170 597884 10226
rect 597456 10046 597512 10102
rect 597580 10046 597636 10102
rect 597704 10046 597760 10102
rect 597828 10046 597884 10102
rect 597456 9922 597512 9978
rect 597580 9922 597636 9978
rect 597704 9922 597760 9978
rect 597828 9922 597884 9978
rect 592914 -1176 592970 -1120
rect 593038 -1176 593094 -1120
rect 593162 -1176 593218 -1120
rect 593286 -1176 593342 -1120
rect 592914 -1300 592970 -1244
rect 593038 -1300 593094 -1244
rect 593162 -1300 593218 -1244
rect 593286 -1300 593342 -1244
rect 592914 -1424 592970 -1368
rect 593038 -1424 593094 -1368
rect 593162 -1424 593218 -1368
rect 593286 -1424 593342 -1368
rect 592914 -1548 592970 -1492
rect 593038 -1548 593094 -1492
rect 593162 -1548 593218 -1492
rect 593286 -1548 593342 -1492
rect 597456 -1176 597512 -1120
rect 597580 -1176 597636 -1120
rect 597704 -1176 597760 -1120
rect 597828 -1176 597884 -1120
rect 597456 -1300 597512 -1244
rect 597580 -1300 597636 -1244
rect 597704 -1300 597760 -1244
rect 597828 -1300 597884 -1244
rect 597456 -1424 597512 -1368
rect 597580 -1424 597636 -1368
rect 597704 -1424 597760 -1368
rect 597828 -1424 597884 -1368
rect 597456 -1548 597512 -1492
rect 597580 -1548 597636 -1492
rect 597704 -1548 597760 -1492
rect 597828 -1548 597884 -1492
<< metal5 >>
rect -1916 598172 597980 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 39954 598172
rect 40010 598116 40078 598172
rect 40134 598116 40202 598172
rect 40258 598116 40326 598172
rect 40382 598116 70674 598172
rect 70730 598116 70798 598172
rect 70854 598116 70922 598172
rect 70978 598116 71046 598172
rect 71102 598116 101394 598172
rect 101450 598116 101518 598172
rect 101574 598116 101642 598172
rect 101698 598116 101766 598172
rect 101822 598116 132114 598172
rect 132170 598116 132238 598172
rect 132294 598116 132362 598172
rect 132418 598116 132486 598172
rect 132542 598116 162834 598172
rect 162890 598116 162958 598172
rect 163014 598116 163082 598172
rect 163138 598116 163206 598172
rect 163262 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect -1916 598048 597980 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 39954 598048
rect 40010 597992 40078 598048
rect 40134 597992 40202 598048
rect 40258 597992 40326 598048
rect 40382 597992 70674 598048
rect 70730 597992 70798 598048
rect 70854 597992 70922 598048
rect 70978 597992 71046 598048
rect 71102 597992 101394 598048
rect 101450 597992 101518 598048
rect 101574 597992 101642 598048
rect 101698 597992 101766 598048
rect 101822 597992 132114 598048
rect 132170 597992 132238 598048
rect 132294 597992 132362 598048
rect 132418 597992 132486 598048
rect 132542 597992 162834 598048
rect 162890 597992 162958 598048
rect 163014 597992 163082 598048
rect 163138 597992 163206 598048
rect 163262 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect -1916 597924 597980 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 39954 597924
rect 40010 597868 40078 597924
rect 40134 597868 40202 597924
rect 40258 597868 40326 597924
rect 40382 597868 70674 597924
rect 70730 597868 70798 597924
rect 70854 597868 70922 597924
rect 70978 597868 71046 597924
rect 71102 597868 101394 597924
rect 101450 597868 101518 597924
rect 101574 597868 101642 597924
rect 101698 597868 101766 597924
rect 101822 597868 132114 597924
rect 132170 597868 132238 597924
rect 132294 597868 132362 597924
rect 132418 597868 132486 597924
rect 132542 597868 162834 597924
rect 162890 597868 162958 597924
rect 163014 597868 163082 597924
rect 163138 597868 163206 597924
rect 163262 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect -1916 597800 597980 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 39954 597800
rect 40010 597744 40078 597800
rect 40134 597744 40202 597800
rect 40258 597744 40326 597800
rect 40382 597744 70674 597800
rect 70730 597744 70798 597800
rect 70854 597744 70922 597800
rect 70978 597744 71046 597800
rect 71102 597744 101394 597800
rect 101450 597744 101518 597800
rect 101574 597744 101642 597800
rect 101698 597744 101766 597800
rect 101822 597744 132114 597800
rect 132170 597744 132238 597800
rect 132294 597744 132362 597800
rect 132418 597744 132486 597800
rect 132542 597744 162834 597800
rect 162890 597744 162958 597800
rect 163014 597744 163082 597800
rect 163138 597744 163206 597800
rect 163262 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect -1916 597648 597980 597744
rect -956 597212 597020 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 36234 597212
rect 36290 597156 36358 597212
rect 36414 597156 36482 597212
rect 36538 597156 36606 597212
rect 36662 597156 66954 597212
rect 67010 597156 67078 597212
rect 67134 597156 67202 597212
rect 67258 597156 67326 597212
rect 67382 597156 97674 597212
rect 97730 597156 97798 597212
rect 97854 597156 97922 597212
rect 97978 597156 98046 597212
rect 98102 597156 128394 597212
rect 128450 597156 128518 597212
rect 128574 597156 128642 597212
rect 128698 597156 128766 597212
rect 128822 597156 159114 597212
rect 159170 597156 159238 597212
rect 159294 597156 159362 597212
rect 159418 597156 159486 597212
rect 159542 597156 189834 597212
rect 189890 597156 189958 597212
rect 190014 597156 190082 597212
rect 190138 597156 190206 597212
rect 190262 597156 220554 597212
rect 220610 597156 220678 597212
rect 220734 597156 220802 597212
rect 220858 597156 220926 597212
rect 220982 597156 251274 597212
rect 251330 597156 251398 597212
rect 251454 597156 251522 597212
rect 251578 597156 251646 597212
rect 251702 597156 281994 597212
rect 282050 597156 282118 597212
rect 282174 597156 282242 597212
rect 282298 597156 282366 597212
rect 282422 597156 312714 597212
rect 312770 597156 312838 597212
rect 312894 597156 312962 597212
rect 313018 597156 313086 597212
rect 313142 597156 343434 597212
rect 343490 597156 343558 597212
rect 343614 597156 343682 597212
rect 343738 597156 343806 597212
rect 343862 597156 374154 597212
rect 374210 597156 374278 597212
rect 374334 597156 374402 597212
rect 374458 597156 374526 597212
rect 374582 597156 404874 597212
rect 404930 597156 404998 597212
rect 405054 597156 405122 597212
rect 405178 597156 405246 597212
rect 405302 597156 435594 597212
rect 435650 597156 435718 597212
rect 435774 597156 435842 597212
rect 435898 597156 435966 597212
rect 436022 597156 466314 597212
rect 466370 597156 466438 597212
rect 466494 597156 466562 597212
rect 466618 597156 466686 597212
rect 466742 597156 497034 597212
rect 497090 597156 497158 597212
rect 497214 597156 497282 597212
rect 497338 597156 497406 597212
rect 497462 597156 527754 597212
rect 527810 597156 527878 597212
rect 527934 597156 528002 597212
rect 528058 597156 528126 597212
rect 528182 597156 558474 597212
rect 558530 597156 558598 597212
rect 558654 597156 558722 597212
rect 558778 597156 558846 597212
rect 558902 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect -956 597088 597020 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 36234 597088
rect 36290 597032 36358 597088
rect 36414 597032 36482 597088
rect 36538 597032 36606 597088
rect 36662 597032 66954 597088
rect 67010 597032 67078 597088
rect 67134 597032 67202 597088
rect 67258 597032 67326 597088
rect 67382 597032 97674 597088
rect 97730 597032 97798 597088
rect 97854 597032 97922 597088
rect 97978 597032 98046 597088
rect 98102 597032 128394 597088
rect 128450 597032 128518 597088
rect 128574 597032 128642 597088
rect 128698 597032 128766 597088
rect 128822 597032 159114 597088
rect 159170 597032 159238 597088
rect 159294 597032 159362 597088
rect 159418 597032 159486 597088
rect 159542 597032 189834 597088
rect 189890 597032 189958 597088
rect 190014 597032 190082 597088
rect 190138 597032 190206 597088
rect 190262 597032 220554 597088
rect 220610 597032 220678 597088
rect 220734 597032 220802 597088
rect 220858 597032 220926 597088
rect 220982 597032 251274 597088
rect 251330 597032 251398 597088
rect 251454 597032 251522 597088
rect 251578 597032 251646 597088
rect 251702 597032 281994 597088
rect 282050 597032 282118 597088
rect 282174 597032 282242 597088
rect 282298 597032 282366 597088
rect 282422 597032 312714 597088
rect 312770 597032 312838 597088
rect 312894 597032 312962 597088
rect 313018 597032 313086 597088
rect 313142 597032 343434 597088
rect 343490 597032 343558 597088
rect 343614 597032 343682 597088
rect 343738 597032 343806 597088
rect 343862 597032 374154 597088
rect 374210 597032 374278 597088
rect 374334 597032 374402 597088
rect 374458 597032 374526 597088
rect 374582 597032 404874 597088
rect 404930 597032 404998 597088
rect 405054 597032 405122 597088
rect 405178 597032 405246 597088
rect 405302 597032 435594 597088
rect 435650 597032 435718 597088
rect 435774 597032 435842 597088
rect 435898 597032 435966 597088
rect 436022 597032 466314 597088
rect 466370 597032 466438 597088
rect 466494 597032 466562 597088
rect 466618 597032 466686 597088
rect 466742 597032 497034 597088
rect 497090 597032 497158 597088
rect 497214 597032 497282 597088
rect 497338 597032 497406 597088
rect 497462 597032 527754 597088
rect 527810 597032 527878 597088
rect 527934 597032 528002 597088
rect 528058 597032 528126 597088
rect 528182 597032 558474 597088
rect 558530 597032 558598 597088
rect 558654 597032 558722 597088
rect 558778 597032 558846 597088
rect 558902 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect -956 596964 597020 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 36234 596964
rect 36290 596908 36358 596964
rect 36414 596908 36482 596964
rect 36538 596908 36606 596964
rect 36662 596908 66954 596964
rect 67010 596908 67078 596964
rect 67134 596908 67202 596964
rect 67258 596908 67326 596964
rect 67382 596908 97674 596964
rect 97730 596908 97798 596964
rect 97854 596908 97922 596964
rect 97978 596908 98046 596964
rect 98102 596908 128394 596964
rect 128450 596908 128518 596964
rect 128574 596908 128642 596964
rect 128698 596908 128766 596964
rect 128822 596908 159114 596964
rect 159170 596908 159238 596964
rect 159294 596908 159362 596964
rect 159418 596908 159486 596964
rect 159542 596908 189834 596964
rect 189890 596908 189958 596964
rect 190014 596908 190082 596964
rect 190138 596908 190206 596964
rect 190262 596908 220554 596964
rect 220610 596908 220678 596964
rect 220734 596908 220802 596964
rect 220858 596908 220926 596964
rect 220982 596908 251274 596964
rect 251330 596908 251398 596964
rect 251454 596908 251522 596964
rect 251578 596908 251646 596964
rect 251702 596908 281994 596964
rect 282050 596908 282118 596964
rect 282174 596908 282242 596964
rect 282298 596908 282366 596964
rect 282422 596908 312714 596964
rect 312770 596908 312838 596964
rect 312894 596908 312962 596964
rect 313018 596908 313086 596964
rect 313142 596908 343434 596964
rect 343490 596908 343558 596964
rect 343614 596908 343682 596964
rect 343738 596908 343806 596964
rect 343862 596908 374154 596964
rect 374210 596908 374278 596964
rect 374334 596908 374402 596964
rect 374458 596908 374526 596964
rect 374582 596908 404874 596964
rect 404930 596908 404998 596964
rect 405054 596908 405122 596964
rect 405178 596908 405246 596964
rect 405302 596908 435594 596964
rect 435650 596908 435718 596964
rect 435774 596908 435842 596964
rect 435898 596908 435966 596964
rect 436022 596908 466314 596964
rect 466370 596908 466438 596964
rect 466494 596908 466562 596964
rect 466618 596908 466686 596964
rect 466742 596908 497034 596964
rect 497090 596908 497158 596964
rect 497214 596908 497282 596964
rect 497338 596908 497406 596964
rect 497462 596908 527754 596964
rect 527810 596908 527878 596964
rect 527934 596908 528002 596964
rect 528058 596908 528126 596964
rect 528182 596908 558474 596964
rect 558530 596908 558598 596964
rect 558654 596908 558722 596964
rect 558778 596908 558846 596964
rect 558902 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect -956 596840 597020 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 36234 596840
rect 36290 596784 36358 596840
rect 36414 596784 36482 596840
rect 36538 596784 36606 596840
rect 36662 596784 66954 596840
rect 67010 596784 67078 596840
rect 67134 596784 67202 596840
rect 67258 596784 67326 596840
rect 67382 596784 97674 596840
rect 97730 596784 97798 596840
rect 97854 596784 97922 596840
rect 97978 596784 98046 596840
rect 98102 596784 128394 596840
rect 128450 596784 128518 596840
rect 128574 596784 128642 596840
rect 128698 596784 128766 596840
rect 128822 596784 159114 596840
rect 159170 596784 159238 596840
rect 159294 596784 159362 596840
rect 159418 596784 159486 596840
rect 159542 596784 189834 596840
rect 189890 596784 189958 596840
rect 190014 596784 190082 596840
rect 190138 596784 190206 596840
rect 190262 596784 220554 596840
rect 220610 596784 220678 596840
rect 220734 596784 220802 596840
rect 220858 596784 220926 596840
rect 220982 596784 251274 596840
rect 251330 596784 251398 596840
rect 251454 596784 251522 596840
rect 251578 596784 251646 596840
rect 251702 596784 281994 596840
rect 282050 596784 282118 596840
rect 282174 596784 282242 596840
rect 282298 596784 282366 596840
rect 282422 596784 312714 596840
rect 312770 596784 312838 596840
rect 312894 596784 312962 596840
rect 313018 596784 313086 596840
rect 313142 596784 343434 596840
rect 343490 596784 343558 596840
rect 343614 596784 343682 596840
rect 343738 596784 343806 596840
rect 343862 596784 374154 596840
rect 374210 596784 374278 596840
rect 374334 596784 374402 596840
rect 374458 596784 374526 596840
rect 374582 596784 404874 596840
rect 404930 596784 404998 596840
rect 405054 596784 405122 596840
rect 405178 596784 405246 596840
rect 405302 596784 435594 596840
rect 435650 596784 435718 596840
rect 435774 596784 435842 596840
rect 435898 596784 435966 596840
rect 436022 596784 466314 596840
rect 466370 596784 466438 596840
rect 466494 596784 466562 596840
rect 466618 596784 466686 596840
rect 466742 596784 497034 596840
rect 497090 596784 497158 596840
rect 497214 596784 497282 596840
rect 497338 596784 497406 596840
rect 497462 596784 527754 596840
rect 527810 596784 527878 596840
rect 527934 596784 528002 596840
rect 528058 596784 528126 596840
rect 528182 596784 558474 596840
rect 558530 596784 558598 596840
rect 558654 596784 558722 596840
rect 558778 596784 558846 596840
rect 558902 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect -956 596688 597020 596784
rect 190636 589978 408340 589994
rect 190636 589922 190652 589978
rect 190708 589922 408268 589978
rect 408324 589922 408340 589978
rect 190636 589906 408340 589922
rect 193100 589798 474420 589814
rect 193100 589742 193116 589798
rect 193172 589742 474348 589798
rect 474404 589742 474420 589798
rect 193100 589726 474420 589742
rect -1916 586350 597980 586446
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 39954 586350
rect 40010 586294 40078 586350
rect 40134 586294 40202 586350
rect 40258 586294 40326 586350
rect 40382 586294 70674 586350
rect 70730 586294 70798 586350
rect 70854 586294 70922 586350
rect 70978 586294 71046 586350
rect 71102 586294 101394 586350
rect 101450 586294 101518 586350
rect 101574 586294 101642 586350
rect 101698 586294 101766 586350
rect 101822 586294 132114 586350
rect 132170 586294 132238 586350
rect 132294 586294 132362 586350
rect 132418 586294 132486 586350
rect 132542 586294 162834 586350
rect 162890 586294 162958 586350
rect 163014 586294 163082 586350
rect 163138 586294 163206 586350
rect 163262 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect -1916 586226 597980 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 39954 586226
rect 40010 586170 40078 586226
rect 40134 586170 40202 586226
rect 40258 586170 40326 586226
rect 40382 586170 70674 586226
rect 70730 586170 70798 586226
rect 70854 586170 70922 586226
rect 70978 586170 71046 586226
rect 71102 586170 101394 586226
rect 101450 586170 101518 586226
rect 101574 586170 101642 586226
rect 101698 586170 101766 586226
rect 101822 586170 132114 586226
rect 132170 586170 132238 586226
rect 132294 586170 132362 586226
rect 132418 586170 132486 586226
rect 132542 586170 162834 586226
rect 162890 586170 162958 586226
rect 163014 586170 163082 586226
rect 163138 586170 163206 586226
rect 163262 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect -1916 586102 597980 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 39954 586102
rect 40010 586046 40078 586102
rect 40134 586046 40202 586102
rect 40258 586046 40326 586102
rect 40382 586046 70674 586102
rect 70730 586046 70798 586102
rect 70854 586046 70922 586102
rect 70978 586046 71046 586102
rect 71102 586046 101394 586102
rect 101450 586046 101518 586102
rect 101574 586046 101642 586102
rect 101698 586046 101766 586102
rect 101822 586046 132114 586102
rect 132170 586046 132238 586102
rect 132294 586046 132362 586102
rect 132418 586046 132486 586102
rect 132542 586046 162834 586102
rect 162890 586046 162958 586102
rect 163014 586046 163082 586102
rect 163138 586046 163206 586102
rect 163262 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect -1916 585978 597980 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 39954 585978
rect 40010 585922 40078 585978
rect 40134 585922 40202 585978
rect 40258 585922 40326 585978
rect 40382 585922 70674 585978
rect 70730 585922 70798 585978
rect 70854 585922 70922 585978
rect 70978 585922 71046 585978
rect 71102 585922 101394 585978
rect 101450 585922 101518 585978
rect 101574 585922 101642 585978
rect 101698 585922 101766 585978
rect 101822 585922 132114 585978
rect 132170 585922 132238 585978
rect 132294 585922 132362 585978
rect 132418 585922 132486 585978
rect 132542 585922 162834 585978
rect 162890 585922 162958 585978
rect 163014 585922 163082 585978
rect 163138 585922 163206 585978
rect 163262 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect -1916 585826 597980 585922
rect -1916 580350 597980 580446
rect -1916 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 36234 580350
rect 36290 580294 36358 580350
rect 36414 580294 36482 580350
rect 36538 580294 36606 580350
rect 36662 580294 66954 580350
rect 67010 580294 67078 580350
rect 67134 580294 67202 580350
rect 67258 580294 67326 580350
rect 67382 580294 97674 580350
rect 97730 580294 97798 580350
rect 97854 580294 97922 580350
rect 97978 580294 98046 580350
rect 98102 580294 128394 580350
rect 128450 580294 128518 580350
rect 128574 580294 128642 580350
rect 128698 580294 128766 580350
rect 128822 580294 159114 580350
rect 159170 580294 159238 580350
rect 159294 580294 159362 580350
rect 159418 580294 159486 580350
rect 159542 580294 189834 580350
rect 189890 580294 189958 580350
rect 190014 580294 190082 580350
rect 190138 580294 190206 580350
rect 190262 580294 220554 580350
rect 220610 580294 220678 580350
rect 220734 580294 220802 580350
rect 220858 580294 220926 580350
rect 220982 580294 251274 580350
rect 251330 580294 251398 580350
rect 251454 580294 251522 580350
rect 251578 580294 251646 580350
rect 251702 580294 281994 580350
rect 282050 580294 282118 580350
rect 282174 580294 282242 580350
rect 282298 580294 282366 580350
rect 282422 580294 312714 580350
rect 312770 580294 312838 580350
rect 312894 580294 312962 580350
rect 313018 580294 313086 580350
rect 313142 580294 343434 580350
rect 343490 580294 343558 580350
rect 343614 580294 343682 580350
rect 343738 580294 343806 580350
rect 343862 580294 374154 580350
rect 374210 580294 374278 580350
rect 374334 580294 374402 580350
rect 374458 580294 374526 580350
rect 374582 580294 404874 580350
rect 404930 580294 404998 580350
rect 405054 580294 405122 580350
rect 405178 580294 405246 580350
rect 405302 580294 435594 580350
rect 435650 580294 435718 580350
rect 435774 580294 435842 580350
rect 435898 580294 435966 580350
rect 436022 580294 466314 580350
rect 466370 580294 466438 580350
rect 466494 580294 466562 580350
rect 466618 580294 466686 580350
rect 466742 580294 497034 580350
rect 497090 580294 497158 580350
rect 497214 580294 497282 580350
rect 497338 580294 497406 580350
rect 497462 580294 527754 580350
rect 527810 580294 527878 580350
rect 527934 580294 528002 580350
rect 528058 580294 528126 580350
rect 528182 580294 558474 580350
rect 558530 580294 558598 580350
rect 558654 580294 558722 580350
rect 558778 580294 558846 580350
rect 558902 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597980 580350
rect -1916 580226 597980 580294
rect -1916 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 36234 580226
rect 36290 580170 36358 580226
rect 36414 580170 36482 580226
rect 36538 580170 36606 580226
rect 36662 580170 66954 580226
rect 67010 580170 67078 580226
rect 67134 580170 67202 580226
rect 67258 580170 67326 580226
rect 67382 580170 97674 580226
rect 97730 580170 97798 580226
rect 97854 580170 97922 580226
rect 97978 580170 98046 580226
rect 98102 580170 128394 580226
rect 128450 580170 128518 580226
rect 128574 580170 128642 580226
rect 128698 580170 128766 580226
rect 128822 580170 159114 580226
rect 159170 580170 159238 580226
rect 159294 580170 159362 580226
rect 159418 580170 159486 580226
rect 159542 580170 189834 580226
rect 189890 580170 189958 580226
rect 190014 580170 190082 580226
rect 190138 580170 190206 580226
rect 190262 580170 220554 580226
rect 220610 580170 220678 580226
rect 220734 580170 220802 580226
rect 220858 580170 220926 580226
rect 220982 580170 251274 580226
rect 251330 580170 251398 580226
rect 251454 580170 251522 580226
rect 251578 580170 251646 580226
rect 251702 580170 281994 580226
rect 282050 580170 282118 580226
rect 282174 580170 282242 580226
rect 282298 580170 282366 580226
rect 282422 580170 312714 580226
rect 312770 580170 312838 580226
rect 312894 580170 312962 580226
rect 313018 580170 313086 580226
rect 313142 580170 343434 580226
rect 343490 580170 343558 580226
rect 343614 580170 343682 580226
rect 343738 580170 343806 580226
rect 343862 580170 374154 580226
rect 374210 580170 374278 580226
rect 374334 580170 374402 580226
rect 374458 580170 374526 580226
rect 374582 580170 404874 580226
rect 404930 580170 404998 580226
rect 405054 580170 405122 580226
rect 405178 580170 405246 580226
rect 405302 580170 435594 580226
rect 435650 580170 435718 580226
rect 435774 580170 435842 580226
rect 435898 580170 435966 580226
rect 436022 580170 466314 580226
rect 466370 580170 466438 580226
rect 466494 580170 466562 580226
rect 466618 580170 466686 580226
rect 466742 580170 497034 580226
rect 497090 580170 497158 580226
rect 497214 580170 497282 580226
rect 497338 580170 497406 580226
rect 497462 580170 527754 580226
rect 527810 580170 527878 580226
rect 527934 580170 528002 580226
rect 528058 580170 528126 580226
rect 528182 580170 558474 580226
rect 558530 580170 558598 580226
rect 558654 580170 558722 580226
rect 558778 580170 558846 580226
rect 558902 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597980 580226
rect -1916 580102 597980 580170
rect -1916 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 36234 580102
rect 36290 580046 36358 580102
rect 36414 580046 36482 580102
rect 36538 580046 36606 580102
rect 36662 580046 66954 580102
rect 67010 580046 67078 580102
rect 67134 580046 67202 580102
rect 67258 580046 67326 580102
rect 67382 580046 97674 580102
rect 97730 580046 97798 580102
rect 97854 580046 97922 580102
rect 97978 580046 98046 580102
rect 98102 580046 128394 580102
rect 128450 580046 128518 580102
rect 128574 580046 128642 580102
rect 128698 580046 128766 580102
rect 128822 580046 159114 580102
rect 159170 580046 159238 580102
rect 159294 580046 159362 580102
rect 159418 580046 159486 580102
rect 159542 580046 189834 580102
rect 189890 580046 189958 580102
rect 190014 580046 190082 580102
rect 190138 580046 190206 580102
rect 190262 580046 220554 580102
rect 220610 580046 220678 580102
rect 220734 580046 220802 580102
rect 220858 580046 220926 580102
rect 220982 580046 251274 580102
rect 251330 580046 251398 580102
rect 251454 580046 251522 580102
rect 251578 580046 251646 580102
rect 251702 580046 281994 580102
rect 282050 580046 282118 580102
rect 282174 580046 282242 580102
rect 282298 580046 282366 580102
rect 282422 580046 312714 580102
rect 312770 580046 312838 580102
rect 312894 580046 312962 580102
rect 313018 580046 313086 580102
rect 313142 580046 343434 580102
rect 343490 580046 343558 580102
rect 343614 580046 343682 580102
rect 343738 580046 343806 580102
rect 343862 580046 374154 580102
rect 374210 580046 374278 580102
rect 374334 580046 374402 580102
rect 374458 580046 374526 580102
rect 374582 580046 404874 580102
rect 404930 580046 404998 580102
rect 405054 580046 405122 580102
rect 405178 580046 405246 580102
rect 405302 580046 435594 580102
rect 435650 580046 435718 580102
rect 435774 580046 435842 580102
rect 435898 580046 435966 580102
rect 436022 580046 466314 580102
rect 466370 580046 466438 580102
rect 466494 580046 466562 580102
rect 466618 580046 466686 580102
rect 466742 580046 497034 580102
rect 497090 580046 497158 580102
rect 497214 580046 497282 580102
rect 497338 580046 497406 580102
rect 497462 580046 527754 580102
rect 527810 580046 527878 580102
rect 527934 580046 528002 580102
rect 528058 580046 528126 580102
rect 528182 580046 558474 580102
rect 558530 580046 558598 580102
rect 558654 580046 558722 580102
rect 558778 580046 558846 580102
rect 558902 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597980 580102
rect -1916 579978 597980 580046
rect -1916 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 36234 579978
rect 36290 579922 36358 579978
rect 36414 579922 36482 579978
rect 36538 579922 36606 579978
rect 36662 579922 66954 579978
rect 67010 579922 67078 579978
rect 67134 579922 67202 579978
rect 67258 579922 67326 579978
rect 67382 579922 97674 579978
rect 97730 579922 97798 579978
rect 97854 579922 97922 579978
rect 97978 579922 98046 579978
rect 98102 579922 128394 579978
rect 128450 579922 128518 579978
rect 128574 579922 128642 579978
rect 128698 579922 128766 579978
rect 128822 579922 159114 579978
rect 159170 579922 159238 579978
rect 159294 579922 159362 579978
rect 159418 579922 159486 579978
rect 159542 579922 189834 579978
rect 189890 579922 189958 579978
rect 190014 579922 190082 579978
rect 190138 579922 190206 579978
rect 190262 579922 220554 579978
rect 220610 579922 220678 579978
rect 220734 579922 220802 579978
rect 220858 579922 220926 579978
rect 220982 579922 251274 579978
rect 251330 579922 251398 579978
rect 251454 579922 251522 579978
rect 251578 579922 251646 579978
rect 251702 579922 281994 579978
rect 282050 579922 282118 579978
rect 282174 579922 282242 579978
rect 282298 579922 282366 579978
rect 282422 579922 312714 579978
rect 312770 579922 312838 579978
rect 312894 579922 312962 579978
rect 313018 579922 313086 579978
rect 313142 579922 343434 579978
rect 343490 579922 343558 579978
rect 343614 579922 343682 579978
rect 343738 579922 343806 579978
rect 343862 579922 374154 579978
rect 374210 579922 374278 579978
rect 374334 579922 374402 579978
rect 374458 579922 374526 579978
rect 374582 579922 404874 579978
rect 404930 579922 404998 579978
rect 405054 579922 405122 579978
rect 405178 579922 405246 579978
rect 405302 579922 435594 579978
rect 435650 579922 435718 579978
rect 435774 579922 435842 579978
rect 435898 579922 435966 579978
rect 436022 579922 466314 579978
rect 466370 579922 466438 579978
rect 466494 579922 466562 579978
rect 466618 579922 466686 579978
rect 466742 579922 497034 579978
rect 497090 579922 497158 579978
rect 497214 579922 497282 579978
rect 497338 579922 497406 579978
rect 497462 579922 527754 579978
rect 527810 579922 527878 579978
rect 527934 579922 528002 579978
rect 528058 579922 528126 579978
rect 528182 579922 558474 579978
rect 558530 579922 558598 579978
rect 558654 579922 558722 579978
rect 558778 579922 558846 579978
rect 558902 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597980 579978
rect -1916 579826 597980 579922
rect -1916 568350 597980 568446
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 9234 568350
rect 9290 568294 9358 568350
rect 9414 568294 9482 568350
rect 9538 568294 9606 568350
rect 9662 568294 39954 568350
rect 40010 568294 40078 568350
rect 40134 568294 40202 568350
rect 40258 568294 40326 568350
rect 40382 568294 70674 568350
rect 70730 568294 70798 568350
rect 70854 568294 70922 568350
rect 70978 568294 71046 568350
rect 71102 568294 101394 568350
rect 101450 568294 101518 568350
rect 101574 568294 101642 568350
rect 101698 568294 101766 568350
rect 101822 568294 132114 568350
rect 132170 568294 132238 568350
rect 132294 568294 132362 568350
rect 132418 568294 132486 568350
rect 132542 568294 162834 568350
rect 162890 568294 162958 568350
rect 163014 568294 163082 568350
rect 163138 568294 163206 568350
rect 163262 568294 562194 568350
rect 562250 568294 562318 568350
rect 562374 568294 562442 568350
rect 562498 568294 562566 568350
rect 562622 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect -1916 568226 597980 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 9234 568226
rect 9290 568170 9358 568226
rect 9414 568170 9482 568226
rect 9538 568170 9606 568226
rect 9662 568170 39954 568226
rect 40010 568170 40078 568226
rect 40134 568170 40202 568226
rect 40258 568170 40326 568226
rect 40382 568170 70674 568226
rect 70730 568170 70798 568226
rect 70854 568170 70922 568226
rect 70978 568170 71046 568226
rect 71102 568170 101394 568226
rect 101450 568170 101518 568226
rect 101574 568170 101642 568226
rect 101698 568170 101766 568226
rect 101822 568170 132114 568226
rect 132170 568170 132238 568226
rect 132294 568170 132362 568226
rect 132418 568170 132486 568226
rect 132542 568170 162834 568226
rect 162890 568170 162958 568226
rect 163014 568170 163082 568226
rect 163138 568170 163206 568226
rect 163262 568170 562194 568226
rect 562250 568170 562318 568226
rect 562374 568170 562442 568226
rect 562498 568170 562566 568226
rect 562622 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect -1916 568102 597980 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 9234 568102
rect 9290 568046 9358 568102
rect 9414 568046 9482 568102
rect 9538 568046 9606 568102
rect 9662 568046 39954 568102
rect 40010 568046 40078 568102
rect 40134 568046 40202 568102
rect 40258 568046 40326 568102
rect 40382 568046 70674 568102
rect 70730 568046 70798 568102
rect 70854 568046 70922 568102
rect 70978 568046 71046 568102
rect 71102 568046 101394 568102
rect 101450 568046 101518 568102
rect 101574 568046 101642 568102
rect 101698 568046 101766 568102
rect 101822 568046 132114 568102
rect 132170 568046 132238 568102
rect 132294 568046 132362 568102
rect 132418 568046 132486 568102
rect 132542 568046 162834 568102
rect 162890 568046 162958 568102
rect 163014 568046 163082 568102
rect 163138 568046 163206 568102
rect 163262 568046 562194 568102
rect 562250 568046 562318 568102
rect 562374 568046 562442 568102
rect 562498 568046 562566 568102
rect 562622 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect -1916 567978 597980 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 9234 567978
rect 9290 567922 9358 567978
rect 9414 567922 9482 567978
rect 9538 567922 9606 567978
rect 9662 567922 39954 567978
rect 40010 567922 40078 567978
rect 40134 567922 40202 567978
rect 40258 567922 40326 567978
rect 40382 567922 70674 567978
rect 70730 567922 70798 567978
rect 70854 567922 70922 567978
rect 70978 567922 71046 567978
rect 71102 567922 101394 567978
rect 101450 567922 101518 567978
rect 101574 567922 101642 567978
rect 101698 567922 101766 567978
rect 101822 567922 132114 567978
rect 132170 567922 132238 567978
rect 132294 567922 132362 567978
rect 132418 567922 132486 567978
rect 132542 567922 162834 567978
rect 162890 567922 162958 567978
rect 163014 567922 163082 567978
rect 163138 567922 163206 567978
rect 163262 567922 562194 567978
rect 562250 567922 562318 567978
rect 562374 567922 562442 567978
rect 562498 567922 562566 567978
rect 562622 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect -1916 567826 597980 567922
rect -1916 562350 597980 562446
rect -1916 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 36234 562350
rect 36290 562294 36358 562350
rect 36414 562294 36482 562350
rect 36538 562294 36606 562350
rect 36662 562294 66954 562350
rect 67010 562294 67078 562350
rect 67134 562294 67202 562350
rect 67258 562294 67326 562350
rect 67382 562294 97674 562350
rect 97730 562294 97798 562350
rect 97854 562294 97922 562350
rect 97978 562294 98046 562350
rect 98102 562294 128394 562350
rect 128450 562294 128518 562350
rect 128574 562294 128642 562350
rect 128698 562294 128766 562350
rect 128822 562294 159114 562350
rect 159170 562294 159238 562350
rect 159294 562294 159362 562350
rect 159418 562294 159486 562350
rect 159542 562294 189834 562350
rect 189890 562294 189958 562350
rect 190014 562294 190082 562350
rect 190138 562294 190206 562350
rect 190262 562294 194518 562350
rect 194574 562294 194642 562350
rect 194698 562294 225238 562350
rect 225294 562294 225362 562350
rect 225418 562294 255958 562350
rect 256014 562294 256082 562350
rect 256138 562294 286678 562350
rect 286734 562294 286802 562350
rect 286858 562294 317398 562350
rect 317454 562294 317522 562350
rect 317578 562294 348118 562350
rect 348174 562294 348242 562350
rect 348298 562294 378838 562350
rect 378894 562294 378962 562350
rect 379018 562294 409558 562350
rect 409614 562294 409682 562350
rect 409738 562294 440278 562350
rect 440334 562294 440402 562350
rect 440458 562294 470998 562350
rect 471054 562294 471122 562350
rect 471178 562294 501718 562350
rect 501774 562294 501842 562350
rect 501898 562294 532438 562350
rect 532494 562294 532562 562350
rect 532618 562294 558474 562350
rect 558530 562294 558598 562350
rect 558654 562294 558722 562350
rect 558778 562294 558846 562350
rect 558902 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597980 562350
rect -1916 562226 597980 562294
rect -1916 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 36234 562226
rect 36290 562170 36358 562226
rect 36414 562170 36482 562226
rect 36538 562170 36606 562226
rect 36662 562170 66954 562226
rect 67010 562170 67078 562226
rect 67134 562170 67202 562226
rect 67258 562170 67326 562226
rect 67382 562170 97674 562226
rect 97730 562170 97798 562226
rect 97854 562170 97922 562226
rect 97978 562170 98046 562226
rect 98102 562170 128394 562226
rect 128450 562170 128518 562226
rect 128574 562170 128642 562226
rect 128698 562170 128766 562226
rect 128822 562170 159114 562226
rect 159170 562170 159238 562226
rect 159294 562170 159362 562226
rect 159418 562170 159486 562226
rect 159542 562170 189834 562226
rect 189890 562170 189958 562226
rect 190014 562170 190082 562226
rect 190138 562170 190206 562226
rect 190262 562170 194518 562226
rect 194574 562170 194642 562226
rect 194698 562170 225238 562226
rect 225294 562170 225362 562226
rect 225418 562170 255958 562226
rect 256014 562170 256082 562226
rect 256138 562170 286678 562226
rect 286734 562170 286802 562226
rect 286858 562170 317398 562226
rect 317454 562170 317522 562226
rect 317578 562170 348118 562226
rect 348174 562170 348242 562226
rect 348298 562170 378838 562226
rect 378894 562170 378962 562226
rect 379018 562170 409558 562226
rect 409614 562170 409682 562226
rect 409738 562170 440278 562226
rect 440334 562170 440402 562226
rect 440458 562170 470998 562226
rect 471054 562170 471122 562226
rect 471178 562170 501718 562226
rect 501774 562170 501842 562226
rect 501898 562170 532438 562226
rect 532494 562170 532562 562226
rect 532618 562170 558474 562226
rect 558530 562170 558598 562226
rect 558654 562170 558722 562226
rect 558778 562170 558846 562226
rect 558902 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597980 562226
rect -1916 562102 597980 562170
rect -1916 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 36234 562102
rect 36290 562046 36358 562102
rect 36414 562046 36482 562102
rect 36538 562046 36606 562102
rect 36662 562046 66954 562102
rect 67010 562046 67078 562102
rect 67134 562046 67202 562102
rect 67258 562046 67326 562102
rect 67382 562046 97674 562102
rect 97730 562046 97798 562102
rect 97854 562046 97922 562102
rect 97978 562046 98046 562102
rect 98102 562046 128394 562102
rect 128450 562046 128518 562102
rect 128574 562046 128642 562102
rect 128698 562046 128766 562102
rect 128822 562046 159114 562102
rect 159170 562046 159238 562102
rect 159294 562046 159362 562102
rect 159418 562046 159486 562102
rect 159542 562046 189834 562102
rect 189890 562046 189958 562102
rect 190014 562046 190082 562102
rect 190138 562046 190206 562102
rect 190262 562046 194518 562102
rect 194574 562046 194642 562102
rect 194698 562046 225238 562102
rect 225294 562046 225362 562102
rect 225418 562046 255958 562102
rect 256014 562046 256082 562102
rect 256138 562046 286678 562102
rect 286734 562046 286802 562102
rect 286858 562046 317398 562102
rect 317454 562046 317522 562102
rect 317578 562046 348118 562102
rect 348174 562046 348242 562102
rect 348298 562046 378838 562102
rect 378894 562046 378962 562102
rect 379018 562046 409558 562102
rect 409614 562046 409682 562102
rect 409738 562046 440278 562102
rect 440334 562046 440402 562102
rect 440458 562046 470998 562102
rect 471054 562046 471122 562102
rect 471178 562046 501718 562102
rect 501774 562046 501842 562102
rect 501898 562046 532438 562102
rect 532494 562046 532562 562102
rect 532618 562046 558474 562102
rect 558530 562046 558598 562102
rect 558654 562046 558722 562102
rect 558778 562046 558846 562102
rect 558902 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597980 562102
rect -1916 562003 597980 562046
rect -1916 561978 114035 562003
rect -1916 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 36234 561978
rect 36290 561922 36358 561978
rect 36414 561922 36482 561978
rect 36538 561922 36606 561978
rect 36662 561922 66954 561978
rect 67010 561922 67078 561978
rect 67134 561922 67202 561978
rect 67258 561922 67326 561978
rect 67382 561922 97674 561978
rect 97730 561922 97798 561978
rect 97854 561922 97922 561978
rect 97978 561922 98046 561978
rect 98102 561947 114035 561978
rect 114091 561947 114159 562003
rect 114215 561947 114283 562003
rect 114339 561947 114407 562003
rect 114463 561947 114531 562003
rect 114587 561947 114655 562003
rect 114711 561947 114779 562003
rect 114835 561947 114903 562003
rect 114959 561947 115027 562003
rect 115083 561947 115151 562003
rect 115207 561947 115275 562003
rect 115331 561947 115399 562003
rect 115455 561947 115523 562003
rect 115579 561947 115647 562003
rect 115703 561947 115771 562003
rect 115827 561947 115895 562003
rect 115951 561947 116019 562003
rect 116075 561947 116143 562003
rect 116199 561947 116267 562003
rect 116323 561947 116391 562003
rect 116447 561947 116515 562003
rect 116571 561947 116639 562003
rect 116695 561947 116763 562003
rect 116819 561947 116887 562003
rect 116943 561947 117011 562003
rect 117067 561947 117135 562003
rect 117191 561947 117259 562003
rect 117315 561947 117383 562003
rect 117439 561947 117507 562003
rect 117563 561947 117631 562003
rect 117687 561947 117755 562003
rect 117811 561947 117879 562003
rect 117935 561947 118003 562003
rect 118059 561947 118127 562003
rect 118183 561947 118251 562003
rect 118307 561947 118375 562003
rect 118431 561947 118499 562003
rect 118555 561947 118623 562003
rect 118679 561947 118747 562003
rect 118803 561947 118871 562003
rect 118927 561947 118995 562003
rect 119051 561947 119119 562003
rect 119175 561947 119243 562003
rect 119299 561947 119367 562003
rect 119423 561947 119491 562003
rect 119547 561947 119615 562003
rect 119671 561947 119739 562003
rect 119795 561947 119863 562003
rect 119919 561947 119987 562003
rect 120043 561947 120111 562003
rect 120167 561947 120235 562003
rect 120291 561947 120359 562003
rect 120415 561978 597980 562003
rect 120415 561947 128394 561978
rect 98102 561922 128394 561947
rect 128450 561922 128518 561978
rect 128574 561922 128642 561978
rect 128698 561922 128766 561978
rect 128822 561922 159114 561978
rect 159170 561922 159238 561978
rect 159294 561922 159362 561978
rect 159418 561922 159486 561978
rect 159542 561922 189834 561978
rect 189890 561922 189958 561978
rect 190014 561922 190082 561978
rect 190138 561922 190206 561978
rect 190262 561922 194518 561978
rect 194574 561922 194642 561978
rect 194698 561922 225238 561978
rect 225294 561922 225362 561978
rect 225418 561922 255958 561978
rect 256014 561922 256082 561978
rect 256138 561922 286678 561978
rect 286734 561922 286802 561978
rect 286858 561922 317398 561978
rect 317454 561922 317522 561978
rect 317578 561922 348118 561978
rect 348174 561922 348242 561978
rect 348298 561922 378838 561978
rect 378894 561922 378962 561978
rect 379018 561922 409558 561978
rect 409614 561922 409682 561978
rect 409738 561922 440278 561978
rect 440334 561922 440402 561978
rect 440458 561922 470998 561978
rect 471054 561922 471122 561978
rect 471178 561922 501718 561978
rect 501774 561922 501842 561978
rect 501898 561922 532438 561978
rect 532494 561922 532562 561978
rect 532618 561922 558474 561978
rect 558530 561922 558598 561978
rect 558654 561922 558722 561978
rect 558778 561922 558846 561978
rect 558902 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597980 561978
rect -1916 561826 597980 561922
rect -1916 550350 597980 550446
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 9234 550350
rect 9290 550294 9358 550350
rect 9414 550294 9482 550350
rect 9538 550294 9606 550350
rect 9662 550294 39954 550350
rect 40010 550294 40078 550350
rect 40134 550294 40202 550350
rect 40258 550294 40326 550350
rect 40382 550294 70674 550350
rect 70730 550294 70798 550350
rect 70854 550294 70922 550350
rect 70978 550294 71046 550350
rect 71102 550294 101394 550350
rect 101450 550294 101518 550350
rect 101574 550294 101642 550350
rect 101698 550294 101766 550350
rect 101822 550294 132114 550350
rect 132170 550294 132238 550350
rect 132294 550294 132362 550350
rect 132418 550294 132486 550350
rect 132542 550294 162834 550350
rect 162890 550294 162958 550350
rect 163014 550294 163082 550350
rect 163138 550294 163206 550350
rect 163262 550294 209878 550350
rect 209934 550294 210002 550350
rect 210058 550294 240598 550350
rect 240654 550294 240722 550350
rect 240778 550294 271318 550350
rect 271374 550294 271442 550350
rect 271498 550294 302038 550350
rect 302094 550294 302162 550350
rect 302218 550294 332758 550350
rect 332814 550294 332882 550350
rect 332938 550294 363478 550350
rect 363534 550294 363602 550350
rect 363658 550294 394198 550350
rect 394254 550294 394322 550350
rect 394378 550294 424918 550350
rect 424974 550294 425042 550350
rect 425098 550294 455638 550350
rect 455694 550294 455762 550350
rect 455818 550294 486358 550350
rect 486414 550294 486482 550350
rect 486538 550294 517078 550350
rect 517134 550294 517202 550350
rect 517258 550294 547798 550350
rect 547854 550294 547922 550350
rect 547978 550294 562194 550350
rect 562250 550294 562318 550350
rect 562374 550294 562442 550350
rect 562498 550294 562566 550350
rect 562622 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect -1916 550226 597980 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 9234 550226
rect 9290 550170 9358 550226
rect 9414 550170 9482 550226
rect 9538 550170 9606 550226
rect 9662 550170 39954 550226
rect 40010 550170 40078 550226
rect 40134 550170 40202 550226
rect 40258 550170 40326 550226
rect 40382 550170 70674 550226
rect 70730 550170 70798 550226
rect 70854 550170 70922 550226
rect 70978 550170 71046 550226
rect 71102 550170 101394 550226
rect 101450 550170 101518 550226
rect 101574 550170 101642 550226
rect 101698 550170 101766 550226
rect 101822 550170 132114 550226
rect 132170 550170 132238 550226
rect 132294 550170 132362 550226
rect 132418 550170 132486 550226
rect 132542 550170 162834 550226
rect 162890 550170 162958 550226
rect 163014 550170 163082 550226
rect 163138 550170 163206 550226
rect 163262 550170 209878 550226
rect 209934 550170 210002 550226
rect 210058 550170 240598 550226
rect 240654 550170 240722 550226
rect 240778 550170 271318 550226
rect 271374 550170 271442 550226
rect 271498 550170 302038 550226
rect 302094 550170 302162 550226
rect 302218 550170 332758 550226
rect 332814 550170 332882 550226
rect 332938 550170 363478 550226
rect 363534 550170 363602 550226
rect 363658 550170 394198 550226
rect 394254 550170 394322 550226
rect 394378 550170 424918 550226
rect 424974 550170 425042 550226
rect 425098 550170 455638 550226
rect 455694 550170 455762 550226
rect 455818 550170 486358 550226
rect 486414 550170 486482 550226
rect 486538 550170 517078 550226
rect 517134 550170 517202 550226
rect 517258 550170 547798 550226
rect 547854 550170 547922 550226
rect 547978 550170 562194 550226
rect 562250 550170 562318 550226
rect 562374 550170 562442 550226
rect 562498 550170 562566 550226
rect 562622 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect -1916 550102 597980 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 9234 550102
rect 9290 550046 9358 550102
rect 9414 550046 9482 550102
rect 9538 550046 9606 550102
rect 9662 550046 39954 550102
rect 40010 550046 40078 550102
rect 40134 550046 40202 550102
rect 40258 550046 40326 550102
rect 40382 550046 70674 550102
rect 70730 550046 70798 550102
rect 70854 550046 70922 550102
rect 70978 550046 71046 550102
rect 71102 550046 101394 550102
rect 101450 550046 101518 550102
rect 101574 550046 101642 550102
rect 101698 550046 101766 550102
rect 101822 550046 132114 550102
rect 132170 550046 132238 550102
rect 132294 550046 132362 550102
rect 132418 550046 132486 550102
rect 132542 550046 162834 550102
rect 162890 550046 162958 550102
rect 163014 550046 163082 550102
rect 163138 550046 163206 550102
rect 163262 550046 209878 550102
rect 209934 550046 210002 550102
rect 210058 550046 240598 550102
rect 240654 550046 240722 550102
rect 240778 550046 271318 550102
rect 271374 550046 271442 550102
rect 271498 550046 302038 550102
rect 302094 550046 302162 550102
rect 302218 550046 332758 550102
rect 332814 550046 332882 550102
rect 332938 550046 363478 550102
rect 363534 550046 363602 550102
rect 363658 550046 394198 550102
rect 394254 550046 394322 550102
rect 394378 550046 424918 550102
rect 424974 550046 425042 550102
rect 425098 550046 455638 550102
rect 455694 550046 455762 550102
rect 455818 550046 486358 550102
rect 486414 550046 486482 550102
rect 486538 550046 517078 550102
rect 517134 550046 517202 550102
rect 517258 550046 547798 550102
rect 547854 550046 547922 550102
rect 547978 550046 562194 550102
rect 562250 550046 562318 550102
rect 562374 550046 562442 550102
rect 562498 550046 562566 550102
rect 562622 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect -1916 549978 597980 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 9234 549978
rect 9290 549922 9358 549978
rect 9414 549922 9482 549978
rect 9538 549922 9606 549978
rect 9662 549922 39954 549978
rect 40010 549922 40078 549978
rect 40134 549922 40202 549978
rect 40258 549922 40326 549978
rect 40382 549922 70674 549978
rect 70730 549922 70798 549978
rect 70854 549922 70922 549978
rect 70978 549922 71046 549978
rect 71102 549922 101394 549978
rect 101450 549922 101518 549978
rect 101574 549922 101642 549978
rect 101698 549922 101766 549978
rect 101822 549922 132114 549978
rect 132170 549922 132238 549978
rect 132294 549922 132362 549978
rect 132418 549922 132486 549978
rect 132542 549922 162834 549978
rect 162890 549922 162958 549978
rect 163014 549922 163082 549978
rect 163138 549922 163206 549978
rect 163262 549922 209878 549978
rect 209934 549922 210002 549978
rect 210058 549922 240598 549978
rect 240654 549922 240722 549978
rect 240778 549922 271318 549978
rect 271374 549922 271442 549978
rect 271498 549922 302038 549978
rect 302094 549922 302162 549978
rect 302218 549922 332758 549978
rect 332814 549922 332882 549978
rect 332938 549922 363478 549978
rect 363534 549922 363602 549978
rect 363658 549922 394198 549978
rect 394254 549922 394322 549978
rect 394378 549922 424918 549978
rect 424974 549922 425042 549978
rect 425098 549922 455638 549978
rect 455694 549922 455762 549978
rect 455818 549922 486358 549978
rect 486414 549922 486482 549978
rect 486538 549922 517078 549978
rect 517134 549922 517202 549978
rect 517258 549922 547798 549978
rect 547854 549922 547922 549978
rect 547978 549922 562194 549978
rect 562250 549922 562318 549978
rect 562374 549922 562442 549978
rect 562498 549922 562566 549978
rect 562622 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect -1916 549826 597980 549922
rect -1916 544350 597980 544446
rect -1916 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 36234 544350
rect 36290 544294 36358 544350
rect 36414 544294 36482 544350
rect 36538 544294 36606 544350
rect 36662 544294 66954 544350
rect 67010 544294 67078 544350
rect 67134 544294 67202 544350
rect 67258 544294 67326 544350
rect 67382 544294 97674 544350
rect 97730 544294 97798 544350
rect 97854 544294 97922 544350
rect 97978 544294 98046 544350
rect 98102 544294 128394 544350
rect 128450 544294 128518 544350
rect 128574 544294 128642 544350
rect 128698 544294 128766 544350
rect 128822 544294 159114 544350
rect 159170 544294 159238 544350
rect 159294 544294 159362 544350
rect 159418 544294 159486 544350
rect 159542 544294 189834 544350
rect 189890 544294 189958 544350
rect 190014 544294 190082 544350
rect 190138 544294 190206 544350
rect 190262 544294 194518 544350
rect 194574 544294 194642 544350
rect 194698 544294 225238 544350
rect 225294 544294 225362 544350
rect 225418 544294 255958 544350
rect 256014 544294 256082 544350
rect 256138 544294 286678 544350
rect 286734 544294 286802 544350
rect 286858 544294 317398 544350
rect 317454 544294 317522 544350
rect 317578 544294 348118 544350
rect 348174 544294 348242 544350
rect 348298 544294 378838 544350
rect 378894 544294 378962 544350
rect 379018 544294 409558 544350
rect 409614 544294 409682 544350
rect 409738 544294 440278 544350
rect 440334 544294 440402 544350
rect 440458 544294 470998 544350
rect 471054 544294 471122 544350
rect 471178 544294 501718 544350
rect 501774 544294 501842 544350
rect 501898 544294 532438 544350
rect 532494 544294 532562 544350
rect 532618 544294 558474 544350
rect 558530 544294 558598 544350
rect 558654 544294 558722 544350
rect 558778 544294 558846 544350
rect 558902 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597980 544350
rect -1916 544290 597980 544294
rect -1916 544234 100965 544290
rect 101021 544234 101089 544290
rect 101145 544234 101213 544290
rect 101269 544234 101337 544290
rect 101393 544234 101461 544290
rect 101517 544234 101585 544290
rect 101641 544234 101709 544290
rect 101765 544234 101833 544290
rect 101889 544234 101957 544290
rect 102013 544234 102081 544290
rect 102137 544234 102205 544290
rect 102261 544234 102329 544290
rect 102385 544234 102453 544290
rect 102509 544234 102577 544290
rect 102633 544234 102701 544290
rect 102757 544234 102825 544290
rect 102881 544234 102949 544290
rect 103005 544234 103073 544290
rect 103129 544234 103197 544290
rect 103253 544234 103321 544290
rect 103377 544234 103445 544290
rect 103501 544234 103569 544290
rect 103625 544234 103693 544290
rect 103749 544234 103817 544290
rect 103873 544234 103941 544290
rect 103997 544234 104065 544290
rect 104121 544234 104189 544290
rect 104245 544234 104313 544290
rect 104369 544234 104437 544290
rect 104493 544234 104561 544290
rect 104617 544234 104685 544290
rect 104741 544234 104809 544290
rect 104865 544234 104933 544290
rect 104989 544234 105057 544290
rect 105113 544234 105181 544290
rect 105237 544234 105305 544290
rect 105361 544234 105429 544290
rect 105485 544234 105553 544290
rect 105609 544234 105677 544290
rect 105733 544234 105801 544290
rect 105857 544234 105925 544290
rect 105981 544234 106049 544290
rect 106105 544234 106173 544290
rect 106229 544234 106297 544290
rect 106353 544234 106421 544290
rect 106477 544234 106545 544290
rect 106601 544234 106669 544290
rect 106725 544234 106793 544290
rect 106849 544234 106917 544290
rect 106973 544234 107041 544290
rect 107097 544234 107165 544290
rect 107221 544234 107289 544290
rect 107345 544234 107413 544290
rect 107469 544234 107537 544290
rect 107593 544234 107661 544290
rect 107717 544234 107785 544290
rect 107841 544234 107909 544290
rect 107965 544234 108033 544290
rect 108089 544234 108157 544290
rect 108213 544234 108281 544290
rect 108337 544234 108405 544290
rect 108461 544234 108529 544290
rect 108585 544234 108653 544290
rect 108709 544234 108777 544290
rect 108833 544234 108901 544290
rect 108957 544234 109025 544290
rect 109081 544234 109149 544290
rect 109205 544234 109273 544290
rect 109329 544234 109397 544290
rect 109453 544234 109521 544290
rect 109577 544234 109645 544290
rect 109701 544234 109769 544290
rect 109825 544234 109893 544290
rect 109949 544234 110017 544290
rect 110073 544234 110141 544290
rect 110197 544234 110265 544290
rect 110321 544234 110389 544290
rect 110445 544234 110513 544290
rect 110569 544234 110637 544290
rect 110693 544234 110761 544290
rect 110817 544234 110885 544290
rect 110941 544234 111009 544290
rect 111065 544234 111133 544290
rect 111189 544234 111257 544290
rect 111313 544234 111381 544290
rect 111437 544234 111505 544290
rect 111561 544234 111629 544290
rect 111685 544234 111753 544290
rect 111809 544234 111877 544290
rect 111933 544234 112001 544290
rect 112057 544234 112125 544290
rect 112181 544234 112249 544290
rect 112305 544234 112373 544290
rect 112429 544234 112497 544290
rect 112553 544234 112621 544290
rect 112677 544234 112745 544290
rect 112801 544234 112869 544290
rect 112925 544234 112993 544290
rect 113049 544234 113117 544290
rect 113173 544234 113241 544290
rect 113297 544234 113365 544290
rect 113421 544234 113489 544290
rect 113545 544234 113613 544290
rect 113669 544234 113737 544290
rect 113793 544234 113861 544290
rect 113917 544234 113985 544290
rect 114041 544234 114109 544290
rect 114165 544234 114233 544290
rect 114289 544234 114357 544290
rect 114413 544234 114481 544290
rect 114537 544234 114605 544290
rect 114661 544234 114729 544290
rect 114785 544234 114853 544290
rect 114909 544234 114977 544290
rect 115033 544234 115101 544290
rect 115157 544234 115225 544290
rect 115281 544234 115349 544290
rect 115405 544234 115473 544290
rect 115529 544234 115597 544290
rect 115653 544234 115721 544290
rect 115777 544234 115845 544290
rect 115901 544234 115969 544290
rect 116025 544234 116093 544290
rect 116149 544234 116217 544290
rect 116273 544234 116341 544290
rect 116397 544234 116465 544290
rect 116521 544234 116589 544290
rect 116645 544234 116713 544290
rect 116769 544234 116837 544290
rect 116893 544234 116961 544290
rect 117017 544234 117085 544290
rect 117141 544234 117209 544290
rect 117265 544234 117333 544290
rect 117389 544234 117457 544290
rect 117513 544234 117581 544290
rect 117637 544234 117705 544290
rect 117761 544234 117829 544290
rect 117885 544234 597980 544290
rect -1916 544226 597980 544234
rect -1916 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 36234 544226
rect 36290 544170 36358 544226
rect 36414 544170 36482 544226
rect 36538 544170 36606 544226
rect 36662 544170 66954 544226
rect 67010 544170 67078 544226
rect 67134 544170 67202 544226
rect 67258 544170 67326 544226
rect 67382 544170 97674 544226
rect 97730 544170 97798 544226
rect 97854 544170 97922 544226
rect 97978 544170 98046 544226
rect 98102 544170 128394 544226
rect 128450 544170 128518 544226
rect 128574 544170 128642 544226
rect 128698 544170 128766 544226
rect 128822 544170 159114 544226
rect 159170 544170 159238 544226
rect 159294 544170 159362 544226
rect 159418 544170 159486 544226
rect 159542 544170 189834 544226
rect 189890 544170 189958 544226
rect 190014 544170 190082 544226
rect 190138 544170 190206 544226
rect 190262 544170 194518 544226
rect 194574 544170 194642 544226
rect 194698 544170 225238 544226
rect 225294 544170 225362 544226
rect 225418 544170 255958 544226
rect 256014 544170 256082 544226
rect 256138 544170 286678 544226
rect 286734 544170 286802 544226
rect 286858 544170 317398 544226
rect 317454 544170 317522 544226
rect 317578 544170 348118 544226
rect 348174 544170 348242 544226
rect 348298 544170 378838 544226
rect 378894 544170 378962 544226
rect 379018 544170 409558 544226
rect 409614 544170 409682 544226
rect 409738 544170 440278 544226
rect 440334 544170 440402 544226
rect 440458 544170 470998 544226
rect 471054 544170 471122 544226
rect 471178 544170 501718 544226
rect 501774 544170 501842 544226
rect 501898 544170 532438 544226
rect 532494 544170 532562 544226
rect 532618 544170 558474 544226
rect 558530 544170 558598 544226
rect 558654 544170 558722 544226
rect 558778 544170 558846 544226
rect 558902 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597980 544226
rect -1916 544166 597980 544170
rect -1916 544110 100965 544166
rect 101021 544110 101089 544166
rect 101145 544110 101213 544166
rect 101269 544110 101337 544166
rect 101393 544110 101461 544166
rect 101517 544110 101585 544166
rect 101641 544110 101709 544166
rect 101765 544110 101833 544166
rect 101889 544110 101957 544166
rect 102013 544110 102081 544166
rect 102137 544110 102205 544166
rect 102261 544110 102329 544166
rect 102385 544110 102453 544166
rect 102509 544110 102577 544166
rect 102633 544110 102701 544166
rect 102757 544110 102825 544166
rect 102881 544110 102949 544166
rect 103005 544110 103073 544166
rect 103129 544110 103197 544166
rect 103253 544110 103321 544166
rect 103377 544110 103445 544166
rect 103501 544110 103569 544166
rect 103625 544110 103693 544166
rect 103749 544110 103817 544166
rect 103873 544110 103941 544166
rect 103997 544110 104065 544166
rect 104121 544110 104189 544166
rect 104245 544110 104313 544166
rect 104369 544110 104437 544166
rect 104493 544110 104561 544166
rect 104617 544110 104685 544166
rect 104741 544110 104809 544166
rect 104865 544110 104933 544166
rect 104989 544110 105057 544166
rect 105113 544110 105181 544166
rect 105237 544110 105305 544166
rect 105361 544110 105429 544166
rect 105485 544110 105553 544166
rect 105609 544110 105677 544166
rect 105733 544110 105801 544166
rect 105857 544110 105925 544166
rect 105981 544110 106049 544166
rect 106105 544110 106173 544166
rect 106229 544110 106297 544166
rect 106353 544110 106421 544166
rect 106477 544110 106545 544166
rect 106601 544110 106669 544166
rect 106725 544110 106793 544166
rect 106849 544110 106917 544166
rect 106973 544110 107041 544166
rect 107097 544110 107165 544166
rect 107221 544110 107289 544166
rect 107345 544110 107413 544166
rect 107469 544110 107537 544166
rect 107593 544110 107661 544166
rect 107717 544110 107785 544166
rect 107841 544110 107909 544166
rect 107965 544110 108033 544166
rect 108089 544110 108157 544166
rect 108213 544110 108281 544166
rect 108337 544110 108405 544166
rect 108461 544110 108529 544166
rect 108585 544110 108653 544166
rect 108709 544110 108777 544166
rect 108833 544110 108901 544166
rect 108957 544110 109025 544166
rect 109081 544110 109149 544166
rect 109205 544110 109273 544166
rect 109329 544110 109397 544166
rect 109453 544110 109521 544166
rect 109577 544110 109645 544166
rect 109701 544110 109769 544166
rect 109825 544110 109893 544166
rect 109949 544110 110017 544166
rect 110073 544110 110141 544166
rect 110197 544110 110265 544166
rect 110321 544110 110389 544166
rect 110445 544110 110513 544166
rect 110569 544110 110637 544166
rect 110693 544110 110761 544166
rect 110817 544110 110885 544166
rect 110941 544110 111009 544166
rect 111065 544110 111133 544166
rect 111189 544110 111257 544166
rect 111313 544110 111381 544166
rect 111437 544110 111505 544166
rect 111561 544110 111629 544166
rect 111685 544110 111753 544166
rect 111809 544110 111877 544166
rect 111933 544110 112001 544166
rect 112057 544110 112125 544166
rect 112181 544110 112249 544166
rect 112305 544110 112373 544166
rect 112429 544110 112497 544166
rect 112553 544110 112621 544166
rect 112677 544110 112745 544166
rect 112801 544110 112869 544166
rect 112925 544110 112993 544166
rect 113049 544110 113117 544166
rect 113173 544110 113241 544166
rect 113297 544110 113365 544166
rect 113421 544110 113489 544166
rect 113545 544110 113613 544166
rect 113669 544110 113737 544166
rect 113793 544110 113861 544166
rect 113917 544110 113985 544166
rect 114041 544110 114109 544166
rect 114165 544110 114233 544166
rect 114289 544110 114357 544166
rect 114413 544110 114481 544166
rect 114537 544110 114605 544166
rect 114661 544110 114729 544166
rect 114785 544110 114853 544166
rect 114909 544110 114977 544166
rect 115033 544110 115101 544166
rect 115157 544110 115225 544166
rect 115281 544110 115349 544166
rect 115405 544110 115473 544166
rect 115529 544110 115597 544166
rect 115653 544110 115721 544166
rect 115777 544110 115845 544166
rect 115901 544110 115969 544166
rect 116025 544110 116093 544166
rect 116149 544110 116217 544166
rect 116273 544110 116341 544166
rect 116397 544110 116465 544166
rect 116521 544110 116589 544166
rect 116645 544110 116713 544166
rect 116769 544110 116837 544166
rect 116893 544110 116961 544166
rect 117017 544110 117085 544166
rect 117141 544110 117209 544166
rect 117265 544110 117333 544166
rect 117389 544110 117457 544166
rect 117513 544110 117581 544166
rect 117637 544110 117705 544166
rect 117761 544110 117829 544166
rect 117885 544110 597980 544166
rect -1916 544102 597980 544110
rect -1916 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 36234 544102
rect 36290 544046 36358 544102
rect 36414 544046 36482 544102
rect 36538 544046 36606 544102
rect 36662 544046 66954 544102
rect 67010 544046 67078 544102
rect 67134 544046 67202 544102
rect 67258 544046 67326 544102
rect 67382 544046 97674 544102
rect 97730 544046 97798 544102
rect 97854 544046 97922 544102
rect 97978 544046 98046 544102
rect 98102 544046 128394 544102
rect 128450 544046 128518 544102
rect 128574 544046 128642 544102
rect 128698 544046 128766 544102
rect 128822 544046 159114 544102
rect 159170 544046 159238 544102
rect 159294 544046 159362 544102
rect 159418 544046 159486 544102
rect 159542 544046 189834 544102
rect 189890 544046 189958 544102
rect 190014 544046 190082 544102
rect 190138 544046 190206 544102
rect 190262 544046 194518 544102
rect 194574 544046 194642 544102
rect 194698 544046 225238 544102
rect 225294 544046 225362 544102
rect 225418 544046 255958 544102
rect 256014 544046 256082 544102
rect 256138 544046 286678 544102
rect 286734 544046 286802 544102
rect 286858 544046 317398 544102
rect 317454 544046 317522 544102
rect 317578 544046 348118 544102
rect 348174 544046 348242 544102
rect 348298 544046 378838 544102
rect 378894 544046 378962 544102
rect 379018 544046 409558 544102
rect 409614 544046 409682 544102
rect 409738 544046 440278 544102
rect 440334 544046 440402 544102
rect 440458 544046 470998 544102
rect 471054 544046 471122 544102
rect 471178 544046 501718 544102
rect 501774 544046 501842 544102
rect 501898 544046 532438 544102
rect 532494 544046 532562 544102
rect 532618 544046 558474 544102
rect 558530 544046 558598 544102
rect 558654 544046 558722 544102
rect 558778 544046 558846 544102
rect 558902 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597980 544102
rect -1916 543978 597980 544046
rect -1916 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 36234 543978
rect 36290 543922 36358 543978
rect 36414 543922 36482 543978
rect 36538 543922 36606 543978
rect 36662 543922 66954 543978
rect 67010 543922 67078 543978
rect 67134 543922 67202 543978
rect 67258 543922 67326 543978
rect 67382 543922 97674 543978
rect 97730 543922 97798 543978
rect 97854 543922 97922 543978
rect 97978 543922 98046 543978
rect 98102 543922 128394 543978
rect 128450 543922 128518 543978
rect 128574 543922 128642 543978
rect 128698 543922 128766 543978
rect 128822 543922 159114 543978
rect 159170 543922 159238 543978
rect 159294 543922 159362 543978
rect 159418 543922 159486 543978
rect 159542 543922 189834 543978
rect 189890 543922 189958 543978
rect 190014 543922 190082 543978
rect 190138 543922 190206 543978
rect 190262 543922 194518 543978
rect 194574 543922 194642 543978
rect 194698 543922 225238 543978
rect 225294 543922 225362 543978
rect 225418 543922 255958 543978
rect 256014 543922 256082 543978
rect 256138 543922 286678 543978
rect 286734 543922 286802 543978
rect 286858 543922 317398 543978
rect 317454 543922 317522 543978
rect 317578 543922 348118 543978
rect 348174 543922 348242 543978
rect 348298 543922 378838 543978
rect 378894 543922 378962 543978
rect 379018 543922 409558 543978
rect 409614 543922 409682 543978
rect 409738 543922 440278 543978
rect 440334 543922 440402 543978
rect 440458 543922 470998 543978
rect 471054 543922 471122 543978
rect 471178 543922 501718 543978
rect 501774 543922 501842 543978
rect 501898 543922 532438 543978
rect 532494 543922 532562 543978
rect 532618 543922 558474 543978
rect 558530 543922 558598 543978
rect 558654 543922 558722 543978
rect 558778 543922 558846 543978
rect 558902 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597980 543978
rect -1916 543891 597980 543922
rect -1916 543835 100823 543891
rect 100879 543835 100927 543891
rect 100983 543835 101031 543891
rect 101087 543835 101135 543891
rect 101191 543835 101239 543891
rect 101295 543835 101343 543891
rect 101399 543835 101447 543891
rect 101503 543835 101551 543891
rect 101607 543835 101655 543891
rect 101711 543835 101759 543891
rect 101815 543835 101863 543891
rect 101919 543835 101967 543891
rect 102023 543835 102071 543891
rect 102127 543835 102175 543891
rect 102231 543835 102279 543891
rect 102335 543835 102383 543891
rect 102439 543835 102487 543891
rect 102543 543835 102591 543891
rect 102647 543835 102695 543891
rect 102751 543835 102799 543891
rect 102855 543835 102903 543891
rect 102959 543835 103007 543891
rect 103063 543835 103111 543891
rect 103167 543835 103215 543891
rect 103271 543835 103319 543891
rect 103375 543835 103423 543891
rect 103479 543835 103527 543891
rect 103583 543835 103631 543891
rect 103687 543835 103735 543891
rect 103791 543835 103839 543891
rect 103895 543835 103943 543891
rect 103999 543835 104047 543891
rect 104103 543835 104151 543891
rect 104207 543835 104255 543891
rect 104311 543835 104359 543891
rect 104415 543835 104463 543891
rect 104519 543835 104567 543891
rect 104623 543835 104671 543891
rect 104727 543835 104775 543891
rect 104831 543835 104879 543891
rect 104935 543835 104983 543891
rect 105039 543835 105087 543891
rect 105143 543835 105191 543891
rect 105247 543835 105295 543891
rect 105351 543835 105399 543891
rect 105455 543835 105503 543891
rect 105559 543835 105607 543891
rect 105663 543835 105711 543891
rect 105767 543835 105815 543891
rect 105871 543835 105919 543891
rect 105975 543835 106023 543891
rect 106079 543835 106127 543891
rect 106183 543835 106231 543891
rect 106287 543835 106335 543891
rect 106391 543835 106439 543891
rect 106495 543835 106543 543891
rect 106599 543835 106647 543891
rect 106703 543835 106751 543891
rect 106807 543835 106855 543891
rect 106911 543835 106959 543891
rect 107015 543835 107063 543891
rect 107119 543835 107167 543891
rect 107223 543835 107271 543891
rect 107327 543835 107375 543891
rect 107431 543835 107479 543891
rect 107535 543835 107583 543891
rect 107639 543835 107687 543891
rect 107743 543835 107791 543891
rect 107847 543835 107895 543891
rect 107951 543835 107999 543891
rect 108055 543835 108103 543891
rect 108159 543835 108207 543891
rect 108263 543835 108311 543891
rect 108367 543835 108415 543891
rect 108471 543835 108519 543891
rect 108575 543835 108623 543891
rect 108679 543835 108727 543891
rect 108783 543835 108831 543891
rect 108887 543835 108935 543891
rect 108991 543835 109039 543891
rect 109095 543835 109143 543891
rect 109199 543835 109247 543891
rect 109303 543835 109351 543891
rect 109407 543835 109455 543891
rect 109511 543835 109559 543891
rect 109615 543835 109663 543891
rect 109719 543835 109767 543891
rect 109823 543835 109871 543891
rect 109927 543835 109975 543891
rect 110031 543835 110079 543891
rect 110135 543835 110183 543891
rect 110239 543835 110287 543891
rect 110343 543835 110391 543891
rect 110447 543835 110495 543891
rect 110551 543835 110599 543891
rect 110655 543835 110703 543891
rect 110759 543835 110807 543891
rect 110863 543835 110911 543891
rect 110967 543835 111015 543891
rect 111071 543835 111119 543891
rect 111175 543835 111223 543891
rect 111279 543835 111327 543891
rect 111383 543835 111431 543891
rect 111487 543835 111535 543891
rect 111591 543835 111639 543891
rect 111695 543835 111743 543891
rect 111799 543835 111847 543891
rect 111903 543835 111951 543891
rect 112007 543835 112055 543891
rect 112111 543835 112159 543891
rect 112215 543835 112263 543891
rect 112319 543835 112367 543891
rect 112423 543835 112471 543891
rect 112527 543835 112575 543891
rect 112631 543835 112679 543891
rect 112735 543835 112783 543891
rect 112839 543835 112887 543891
rect 112943 543835 112991 543891
rect 113047 543835 113095 543891
rect 113151 543835 113199 543891
rect 113255 543835 113303 543891
rect 113359 543835 113407 543891
rect 113463 543835 113511 543891
rect 113567 543835 113615 543891
rect 113671 543835 113719 543891
rect 113775 543835 113823 543891
rect 113879 543835 113927 543891
rect 113983 543835 114031 543891
rect 114087 543835 114135 543891
rect 114191 543835 114239 543891
rect 114295 543835 114343 543891
rect 114399 543835 114447 543891
rect 114503 543835 114551 543891
rect 114607 543835 114655 543891
rect 114711 543835 114759 543891
rect 114815 543835 114863 543891
rect 114919 543835 114967 543891
rect 115023 543835 115071 543891
rect 115127 543835 115175 543891
rect 115231 543835 115279 543891
rect 115335 543835 115383 543891
rect 115439 543835 115487 543891
rect 115543 543835 115591 543891
rect 115647 543835 115695 543891
rect 115751 543835 115799 543891
rect 115855 543835 115903 543891
rect 115959 543835 116007 543891
rect 116063 543835 116111 543891
rect 116167 543835 116215 543891
rect 116271 543835 116319 543891
rect 116375 543835 116423 543891
rect 116479 543835 116527 543891
rect 116583 543835 116631 543891
rect 116687 543835 116735 543891
rect 116791 543835 116839 543891
rect 116895 543835 116943 543891
rect 116999 543835 117047 543891
rect 117103 543835 117151 543891
rect 117207 543835 117255 543891
rect 117311 543835 117359 543891
rect 117415 543835 117463 543891
rect 117519 543835 117567 543891
rect 117623 543835 117671 543891
rect 117727 543835 597980 543891
rect -1916 543826 597980 543835
rect -1916 532350 597980 532446
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 9234 532350
rect 9290 532294 9358 532350
rect 9414 532294 9482 532350
rect 9538 532294 9606 532350
rect 9662 532294 39954 532350
rect 40010 532294 40078 532350
rect 40134 532294 40202 532350
rect 40258 532294 40326 532350
rect 40382 532303 162834 532350
rect 40382 532294 69507 532303
rect -1916 532247 69507 532294
rect 69563 532247 69631 532303
rect 69687 532247 69755 532303
rect 69811 532247 69879 532303
rect 69935 532247 70003 532303
rect 70059 532247 70127 532303
rect 70183 532247 70251 532303
rect 70307 532247 70375 532303
rect 70431 532247 70499 532303
rect 70555 532247 70623 532303
rect 70679 532247 70747 532303
rect 70803 532247 70871 532303
rect 70927 532247 70995 532303
rect 71051 532247 71119 532303
rect 71175 532247 71243 532303
rect 71299 532247 71367 532303
rect 71423 532247 71491 532303
rect 71547 532247 71615 532303
rect 71671 532247 71739 532303
rect 71795 532247 71863 532303
rect 71919 532247 71987 532303
rect 72043 532247 72111 532303
rect 72167 532247 72235 532303
rect 72291 532247 72359 532303
rect 72415 532247 72483 532303
rect 72539 532247 72607 532303
rect 72663 532247 72731 532303
rect 72787 532247 72855 532303
rect 72911 532247 72979 532303
rect 73035 532247 73103 532303
rect 73159 532247 73227 532303
rect 73283 532247 73351 532303
rect 73407 532247 73475 532303
rect 73531 532247 73599 532303
rect 73655 532247 73723 532303
rect 73779 532247 73847 532303
rect 73903 532247 73971 532303
rect 74027 532247 74095 532303
rect 74151 532247 74219 532303
rect 74275 532247 74343 532303
rect 74399 532247 74467 532303
rect 74523 532247 74591 532303
rect 74647 532247 74715 532303
rect 74771 532247 74839 532303
rect 74895 532247 74963 532303
rect 75019 532247 75087 532303
rect 75143 532247 75211 532303
rect 75267 532247 75335 532303
rect 75391 532247 75459 532303
rect 75515 532247 75583 532303
rect 75639 532247 75707 532303
rect 75763 532247 75831 532303
rect 75887 532247 75955 532303
rect 76011 532247 76079 532303
rect 76135 532247 76203 532303
rect 76259 532247 76327 532303
rect 76383 532247 76451 532303
rect 76507 532247 76575 532303
rect 76631 532247 76699 532303
rect 76755 532247 76823 532303
rect 76879 532247 76947 532303
rect 77003 532247 77071 532303
rect 77127 532247 77195 532303
rect 77251 532247 77319 532303
rect 77375 532247 77443 532303
rect 77499 532247 77567 532303
rect 77623 532247 77691 532303
rect 77747 532247 77815 532303
rect 77871 532247 77939 532303
rect 77995 532247 78063 532303
rect 78119 532247 78187 532303
rect 78243 532294 162834 532303
rect 162890 532294 162958 532350
rect 163014 532294 163082 532350
rect 163138 532294 163206 532350
rect 163262 532294 209878 532350
rect 209934 532294 210002 532350
rect 210058 532294 240598 532350
rect 240654 532294 240722 532350
rect 240778 532294 271318 532350
rect 271374 532294 271442 532350
rect 271498 532294 302038 532350
rect 302094 532294 302162 532350
rect 302218 532294 332758 532350
rect 332814 532294 332882 532350
rect 332938 532294 363478 532350
rect 363534 532294 363602 532350
rect 363658 532294 394198 532350
rect 394254 532294 394322 532350
rect 394378 532294 424918 532350
rect 424974 532294 425042 532350
rect 425098 532294 455638 532350
rect 455694 532294 455762 532350
rect 455818 532294 486358 532350
rect 486414 532294 486482 532350
rect 486538 532294 517078 532350
rect 517134 532294 517202 532350
rect 517258 532294 547798 532350
rect 547854 532294 547922 532350
rect 547978 532294 562194 532350
rect 562250 532294 562318 532350
rect 562374 532294 562442 532350
rect 562498 532294 562566 532350
rect 562622 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect 78243 532247 597980 532294
rect -1916 532226 597980 532247
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 9234 532226
rect 9290 532170 9358 532226
rect 9414 532170 9482 532226
rect 9538 532170 9606 532226
rect 9662 532170 39954 532226
rect 40010 532170 40078 532226
rect 40134 532170 40202 532226
rect 40258 532170 40326 532226
rect 40382 532170 162834 532226
rect 162890 532170 162958 532226
rect 163014 532170 163082 532226
rect 163138 532170 163206 532226
rect 163262 532170 209878 532226
rect 209934 532170 210002 532226
rect 210058 532170 240598 532226
rect 240654 532170 240722 532226
rect 240778 532170 271318 532226
rect 271374 532170 271442 532226
rect 271498 532170 302038 532226
rect 302094 532170 302162 532226
rect 302218 532170 332758 532226
rect 332814 532170 332882 532226
rect 332938 532170 363478 532226
rect 363534 532170 363602 532226
rect 363658 532170 394198 532226
rect 394254 532170 394322 532226
rect 394378 532170 424918 532226
rect 424974 532170 425042 532226
rect 425098 532170 455638 532226
rect 455694 532170 455762 532226
rect 455818 532170 486358 532226
rect 486414 532170 486482 532226
rect 486538 532170 517078 532226
rect 517134 532170 517202 532226
rect 517258 532170 547798 532226
rect 547854 532170 547922 532226
rect 547978 532170 562194 532226
rect 562250 532170 562318 532226
rect 562374 532170 562442 532226
rect 562498 532170 562566 532226
rect 562622 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect -1916 532102 597980 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 9234 532102
rect 9290 532046 9358 532102
rect 9414 532046 9482 532102
rect 9538 532046 9606 532102
rect 9662 532046 39954 532102
rect 40010 532046 40078 532102
rect 40134 532046 40202 532102
rect 40258 532046 40326 532102
rect 40382 532046 162834 532102
rect 162890 532046 162958 532102
rect 163014 532046 163082 532102
rect 163138 532046 163206 532102
rect 163262 532046 209878 532102
rect 209934 532046 210002 532102
rect 210058 532046 240598 532102
rect 240654 532046 240722 532102
rect 240778 532046 271318 532102
rect 271374 532046 271442 532102
rect 271498 532046 302038 532102
rect 302094 532046 302162 532102
rect 302218 532046 332758 532102
rect 332814 532046 332882 532102
rect 332938 532046 363478 532102
rect 363534 532046 363602 532102
rect 363658 532046 394198 532102
rect 394254 532046 394322 532102
rect 394378 532046 424918 532102
rect 424974 532046 425042 532102
rect 425098 532046 455638 532102
rect 455694 532046 455762 532102
rect 455818 532046 486358 532102
rect 486414 532046 486482 532102
rect 486538 532046 517078 532102
rect 517134 532046 517202 532102
rect 517258 532046 547798 532102
rect 547854 532046 547922 532102
rect 547978 532046 562194 532102
rect 562250 532046 562318 532102
rect 562374 532046 562442 532102
rect 562498 532046 562566 532102
rect 562622 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect -1916 532003 597980 532046
rect -1916 531978 69181 532003
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 9234 531978
rect 9290 531922 9358 531978
rect 9414 531922 9482 531978
rect 9538 531922 9606 531978
rect 9662 531922 39954 531978
rect 40010 531922 40078 531978
rect 40134 531922 40202 531978
rect 40258 531922 40326 531978
rect 40382 531947 69181 531978
rect 69237 531947 69305 532003
rect 69361 531947 69429 532003
rect 69485 531947 69553 532003
rect 69609 531947 69677 532003
rect 69733 531947 69801 532003
rect 69857 531947 69925 532003
rect 69981 531947 70049 532003
rect 70105 531947 70173 532003
rect 70229 531947 70297 532003
rect 70353 531947 70421 532003
rect 70477 531947 70545 532003
rect 70601 531947 70669 532003
rect 70725 531947 70793 532003
rect 70849 531947 70917 532003
rect 70973 531947 71041 532003
rect 71097 531947 71165 532003
rect 71221 531947 71289 532003
rect 71345 531947 71413 532003
rect 71469 531947 71537 532003
rect 71593 531947 71661 532003
rect 71717 531947 71785 532003
rect 71841 531947 71909 532003
rect 71965 531947 72033 532003
rect 72089 531947 72157 532003
rect 72213 531947 72281 532003
rect 72337 531947 72405 532003
rect 72461 531947 72529 532003
rect 72585 531947 72653 532003
rect 72709 531947 72777 532003
rect 72833 531947 72901 532003
rect 72957 531947 73025 532003
rect 73081 531947 73149 532003
rect 73205 531947 73273 532003
rect 73329 531947 73397 532003
rect 73453 531947 73521 532003
rect 73577 531947 73645 532003
rect 73701 531947 73769 532003
rect 73825 531947 73893 532003
rect 73949 531947 74017 532003
rect 74073 531947 74141 532003
rect 74197 531947 74265 532003
rect 74321 531947 74389 532003
rect 74445 531947 74513 532003
rect 74569 531947 74637 532003
rect 74693 531947 74761 532003
rect 74817 531947 74885 532003
rect 74941 531947 75009 532003
rect 75065 531947 75133 532003
rect 75189 531947 75257 532003
rect 75313 531947 75381 532003
rect 75437 531947 75505 532003
rect 75561 531947 75629 532003
rect 75685 531947 75753 532003
rect 75809 531947 75877 532003
rect 75933 531947 76001 532003
rect 76057 531947 76125 532003
rect 76181 531947 76249 532003
rect 76305 531947 76373 532003
rect 76429 531947 76497 532003
rect 76553 531947 76621 532003
rect 76677 531947 76745 532003
rect 76801 531947 76869 532003
rect 76925 531947 76993 532003
rect 77049 531947 77117 532003
rect 77173 531947 77241 532003
rect 77297 531947 77365 532003
rect 77421 531947 77489 532003
rect 77545 531947 77613 532003
rect 77669 531978 597980 532003
rect 77669 531947 162834 531978
rect 40382 531922 162834 531947
rect 162890 531922 162958 531978
rect 163014 531922 163082 531978
rect 163138 531922 163206 531978
rect 163262 531922 209878 531978
rect 209934 531922 210002 531978
rect 210058 531922 240598 531978
rect 240654 531922 240722 531978
rect 240778 531922 271318 531978
rect 271374 531922 271442 531978
rect 271498 531922 302038 531978
rect 302094 531922 302162 531978
rect 302218 531922 332758 531978
rect 332814 531922 332882 531978
rect 332938 531922 363478 531978
rect 363534 531922 363602 531978
rect 363658 531922 394198 531978
rect 394254 531922 394322 531978
rect 394378 531922 424918 531978
rect 424974 531922 425042 531978
rect 425098 531922 455638 531978
rect 455694 531922 455762 531978
rect 455818 531922 486358 531978
rect 486414 531922 486482 531978
rect 486538 531922 517078 531978
rect 517134 531922 517202 531978
rect 517258 531922 547798 531978
rect 547854 531922 547922 531978
rect 547978 531922 562194 531978
rect 562250 531922 562318 531978
rect 562374 531922 562442 531978
rect 562498 531922 562566 531978
rect 562622 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect -1916 531826 597980 531922
rect -1916 526350 597980 526446
rect -1916 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 36234 526350
rect 36290 526294 36358 526350
rect 36414 526294 36482 526350
rect 36538 526294 36606 526350
rect 36662 526294 159114 526350
rect 159170 526294 159238 526350
rect 159294 526294 159362 526350
rect 159418 526294 159486 526350
rect 159542 526294 189834 526350
rect 189890 526294 189958 526350
rect 190014 526294 190082 526350
rect 190138 526294 190206 526350
rect 190262 526294 194518 526350
rect 194574 526294 194642 526350
rect 194698 526294 225238 526350
rect 225294 526294 225362 526350
rect 225418 526294 255958 526350
rect 256014 526294 256082 526350
rect 256138 526294 286678 526350
rect 286734 526294 286802 526350
rect 286858 526294 317398 526350
rect 317454 526294 317522 526350
rect 317578 526294 348118 526350
rect 348174 526294 348242 526350
rect 348298 526294 378838 526350
rect 378894 526294 378962 526350
rect 379018 526294 409558 526350
rect 409614 526294 409682 526350
rect 409738 526294 440278 526350
rect 440334 526294 440402 526350
rect 440458 526294 470998 526350
rect 471054 526294 471122 526350
rect 471178 526294 501718 526350
rect 501774 526294 501842 526350
rect 501898 526294 532438 526350
rect 532494 526294 532562 526350
rect 532618 526294 558474 526350
rect 558530 526294 558598 526350
rect 558654 526294 558722 526350
rect 558778 526294 558846 526350
rect 558902 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597980 526350
rect -1916 526226 597980 526294
rect -1916 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 36234 526226
rect 36290 526170 36358 526226
rect 36414 526170 36482 526226
rect 36538 526170 36606 526226
rect 36662 526170 159114 526226
rect 159170 526170 159238 526226
rect 159294 526170 159362 526226
rect 159418 526170 159486 526226
rect 159542 526170 189834 526226
rect 189890 526170 189958 526226
rect 190014 526170 190082 526226
rect 190138 526170 190206 526226
rect 190262 526170 194518 526226
rect 194574 526170 194642 526226
rect 194698 526170 225238 526226
rect 225294 526170 225362 526226
rect 225418 526170 255958 526226
rect 256014 526170 256082 526226
rect 256138 526170 286678 526226
rect 286734 526170 286802 526226
rect 286858 526170 317398 526226
rect 317454 526170 317522 526226
rect 317578 526170 348118 526226
rect 348174 526170 348242 526226
rect 348298 526170 378838 526226
rect 378894 526170 378962 526226
rect 379018 526170 409558 526226
rect 409614 526170 409682 526226
rect 409738 526170 440278 526226
rect 440334 526170 440402 526226
rect 440458 526170 470998 526226
rect 471054 526170 471122 526226
rect 471178 526170 501718 526226
rect 501774 526170 501842 526226
rect 501898 526170 532438 526226
rect 532494 526170 532562 526226
rect 532618 526170 558474 526226
rect 558530 526170 558598 526226
rect 558654 526170 558722 526226
rect 558778 526170 558846 526226
rect 558902 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597980 526226
rect -1916 526153 597980 526170
rect -1916 526102 91381 526153
rect -1916 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 36234 526102
rect 36290 526046 36358 526102
rect 36414 526046 36482 526102
rect 36538 526046 36606 526102
rect 36662 526097 91381 526102
rect 91437 526097 91505 526153
rect 91561 526097 91629 526153
rect 91685 526097 91753 526153
rect 91809 526097 91877 526153
rect 91933 526097 92001 526153
rect 92057 526097 92125 526153
rect 92181 526097 92249 526153
rect 92305 526097 92373 526153
rect 92429 526097 92497 526153
rect 92553 526097 92621 526153
rect 92677 526097 92745 526153
rect 92801 526097 92869 526153
rect 92925 526097 92993 526153
rect 93049 526097 93117 526153
rect 93173 526097 93241 526153
rect 93297 526097 93365 526153
rect 93421 526097 93489 526153
rect 93545 526097 93613 526153
rect 93669 526097 93737 526153
rect 93793 526097 93861 526153
rect 93917 526097 93985 526153
rect 94041 526097 94109 526153
rect 94165 526097 94233 526153
rect 94289 526097 94357 526153
rect 94413 526097 94481 526153
rect 94537 526097 94605 526153
rect 94661 526097 94729 526153
rect 94785 526097 94853 526153
rect 94909 526097 94977 526153
rect 95033 526097 95101 526153
rect 95157 526097 95225 526153
rect 95281 526097 95349 526153
rect 95405 526097 95473 526153
rect 95529 526097 95597 526153
rect 95653 526097 95721 526153
rect 95777 526097 95845 526153
rect 95901 526097 95969 526153
rect 96025 526097 96093 526153
rect 96149 526097 96217 526153
rect 96273 526097 96341 526153
rect 96397 526097 96465 526153
rect 96521 526097 96589 526153
rect 96645 526097 96713 526153
rect 96769 526097 96837 526153
rect 96893 526097 96961 526153
rect 97017 526097 97085 526153
rect 97141 526097 97209 526153
rect 97265 526097 97333 526153
rect 97389 526097 97457 526153
rect 97513 526097 97581 526153
rect 97637 526097 97705 526153
rect 97761 526097 97829 526153
rect 97885 526097 97953 526153
rect 98009 526097 98077 526153
rect 98133 526097 98201 526153
rect 98257 526097 98325 526153
rect 98381 526097 98449 526153
rect 98505 526097 98573 526153
rect 98629 526097 98697 526153
rect 98753 526097 98821 526153
rect 98877 526097 98945 526153
rect 99001 526097 99069 526153
rect 99125 526097 99193 526153
rect 99249 526097 99317 526153
rect 99373 526097 99441 526153
rect 99497 526097 99565 526153
rect 99621 526097 99689 526153
rect 99745 526097 99813 526153
rect 99869 526097 99937 526153
rect 99993 526097 100061 526153
rect 100117 526097 100185 526153
rect 100241 526097 100309 526153
rect 100365 526097 100433 526153
rect 100489 526097 100557 526153
rect 100613 526097 100681 526153
rect 100737 526097 100805 526153
rect 100861 526097 100929 526153
rect 100985 526097 101053 526153
rect 101109 526097 101177 526153
rect 101233 526097 101301 526153
rect 101357 526097 101425 526153
rect 101481 526097 101549 526153
rect 101605 526097 101673 526153
rect 101729 526097 101797 526153
rect 101853 526097 101921 526153
rect 101977 526097 102045 526153
rect 102101 526097 102169 526153
rect 102225 526097 102293 526153
rect 102349 526097 102417 526153
rect 102473 526097 102541 526153
rect 102597 526097 102665 526153
rect 102721 526097 102789 526153
rect 102845 526097 102913 526153
rect 102969 526097 103037 526153
rect 103093 526097 103161 526153
rect 103217 526097 103285 526153
rect 103341 526097 103409 526153
rect 103465 526097 103533 526153
rect 103589 526097 103657 526153
rect 103713 526097 103781 526153
rect 103837 526097 103905 526153
rect 103961 526097 104029 526153
rect 104085 526097 104153 526153
rect 104209 526097 104277 526153
rect 104333 526097 104401 526153
rect 104457 526097 104525 526153
rect 104581 526097 104649 526153
rect 104705 526097 104773 526153
rect 104829 526097 104897 526153
rect 104953 526097 105021 526153
rect 105077 526097 105145 526153
rect 105201 526097 105269 526153
rect 105325 526097 105393 526153
rect 105449 526097 105517 526153
rect 105573 526097 105641 526153
rect 105697 526097 105765 526153
rect 105821 526097 105889 526153
rect 105945 526097 106013 526153
rect 106069 526097 106137 526153
rect 106193 526097 106261 526153
rect 106317 526097 106385 526153
rect 106441 526097 106509 526153
rect 106565 526097 106633 526153
rect 106689 526097 106757 526153
rect 106813 526097 106881 526153
rect 106937 526097 107005 526153
rect 107061 526097 107129 526153
rect 107185 526097 107253 526153
rect 107309 526097 107377 526153
rect 107433 526097 107501 526153
rect 107557 526097 107625 526153
rect 107681 526097 107749 526153
rect 107805 526097 107873 526153
rect 107929 526097 107997 526153
rect 108053 526097 108121 526153
rect 108177 526097 108245 526153
rect 108301 526097 108369 526153
rect 108425 526097 108493 526153
rect 108549 526097 108617 526153
rect 108673 526097 108741 526153
rect 108797 526097 108865 526153
rect 108921 526097 108989 526153
rect 109045 526097 109113 526153
rect 109169 526102 597980 526153
rect 109169 526097 159114 526102
rect 36662 526046 159114 526097
rect 159170 526046 159238 526102
rect 159294 526046 159362 526102
rect 159418 526046 159486 526102
rect 159542 526046 189834 526102
rect 189890 526046 189958 526102
rect 190014 526046 190082 526102
rect 190138 526046 190206 526102
rect 190262 526046 194518 526102
rect 194574 526046 194642 526102
rect 194698 526046 225238 526102
rect 225294 526046 225362 526102
rect 225418 526046 255958 526102
rect 256014 526046 256082 526102
rect 256138 526046 286678 526102
rect 286734 526046 286802 526102
rect 286858 526046 317398 526102
rect 317454 526046 317522 526102
rect 317578 526046 348118 526102
rect 348174 526046 348242 526102
rect 348298 526046 378838 526102
rect 378894 526046 378962 526102
rect 379018 526046 409558 526102
rect 409614 526046 409682 526102
rect 409738 526046 440278 526102
rect 440334 526046 440402 526102
rect 440458 526046 470998 526102
rect 471054 526046 471122 526102
rect 471178 526046 501718 526102
rect 501774 526046 501842 526102
rect 501898 526046 532438 526102
rect 532494 526046 532562 526102
rect 532618 526046 558474 526102
rect 558530 526046 558598 526102
rect 558654 526046 558722 526102
rect 558778 526046 558846 526102
rect 558902 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597980 526102
rect -1916 525978 597980 526046
rect -1916 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 36234 525978
rect 36290 525922 36358 525978
rect 36414 525922 36482 525978
rect 36538 525922 36606 525978
rect 36662 525922 159114 525978
rect 159170 525922 159238 525978
rect 159294 525922 159362 525978
rect 159418 525922 159486 525978
rect 159542 525922 189834 525978
rect 189890 525922 189958 525978
rect 190014 525922 190082 525978
rect 190138 525922 190206 525978
rect 190262 525922 194518 525978
rect 194574 525922 194642 525978
rect 194698 525922 225238 525978
rect 225294 525922 225362 525978
rect 225418 525922 255958 525978
rect 256014 525922 256082 525978
rect 256138 525922 286678 525978
rect 286734 525922 286802 525978
rect 286858 525922 317398 525978
rect 317454 525922 317522 525978
rect 317578 525922 348118 525978
rect 348174 525922 348242 525978
rect 348298 525922 378838 525978
rect 378894 525922 378962 525978
rect 379018 525922 409558 525978
rect 409614 525922 409682 525978
rect 409738 525922 440278 525978
rect 440334 525922 440402 525978
rect 440458 525922 470998 525978
rect 471054 525922 471122 525978
rect 471178 525922 501718 525978
rect 501774 525922 501842 525978
rect 501898 525922 532438 525978
rect 532494 525922 532562 525978
rect 532618 525922 558474 525978
rect 558530 525922 558598 525978
rect 558654 525922 558722 525978
rect 558778 525922 558846 525978
rect 558902 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597980 525978
rect -1916 525891 597980 525922
rect -1916 525835 91234 525891
rect 91290 525835 91338 525891
rect 91394 525835 91442 525891
rect 91498 525835 91546 525891
rect 91602 525835 91650 525891
rect 91706 525835 91754 525891
rect 91810 525835 91858 525891
rect 91914 525835 91962 525891
rect 92018 525835 92066 525891
rect 92122 525835 92170 525891
rect 92226 525835 92274 525891
rect 92330 525835 92378 525891
rect 92434 525835 92482 525891
rect 92538 525835 92586 525891
rect 92642 525835 92690 525891
rect 92746 525835 92794 525891
rect 92850 525835 92898 525891
rect 92954 525835 93002 525891
rect 93058 525835 93106 525891
rect 93162 525835 93210 525891
rect 93266 525835 93314 525891
rect 93370 525835 93418 525891
rect 93474 525835 93522 525891
rect 93578 525835 93626 525891
rect 93682 525835 93730 525891
rect 93786 525835 93834 525891
rect 93890 525835 93938 525891
rect 93994 525835 94042 525891
rect 94098 525835 94146 525891
rect 94202 525835 94250 525891
rect 94306 525835 94354 525891
rect 94410 525835 94458 525891
rect 94514 525835 94562 525891
rect 94618 525835 94666 525891
rect 94722 525835 94770 525891
rect 94826 525835 94874 525891
rect 94930 525835 94978 525891
rect 95034 525835 95082 525891
rect 95138 525835 95186 525891
rect 95242 525835 95290 525891
rect 95346 525835 95394 525891
rect 95450 525835 95498 525891
rect 95554 525835 95602 525891
rect 95658 525835 95706 525891
rect 95762 525835 95810 525891
rect 95866 525835 95914 525891
rect 95970 525835 96018 525891
rect 96074 525835 96122 525891
rect 96178 525835 96226 525891
rect 96282 525835 96330 525891
rect 96386 525835 96434 525891
rect 96490 525835 96538 525891
rect 96594 525835 96642 525891
rect 96698 525835 96746 525891
rect 96802 525835 96850 525891
rect 96906 525835 96954 525891
rect 97010 525835 97058 525891
rect 97114 525835 97162 525891
rect 97218 525835 97266 525891
rect 97322 525835 97370 525891
rect 97426 525835 97474 525891
rect 97530 525835 97578 525891
rect 97634 525835 97682 525891
rect 97738 525835 97786 525891
rect 97842 525835 97890 525891
rect 97946 525835 97994 525891
rect 98050 525835 98098 525891
rect 98154 525835 98202 525891
rect 98258 525835 98306 525891
rect 98362 525835 98410 525891
rect 98466 525835 98514 525891
rect 98570 525835 98618 525891
rect 98674 525835 98722 525891
rect 98778 525835 98826 525891
rect 98882 525835 98930 525891
rect 98986 525835 99034 525891
rect 99090 525835 99138 525891
rect 99194 525835 99242 525891
rect 99298 525835 99346 525891
rect 99402 525835 99450 525891
rect 99506 525835 99554 525891
rect 99610 525835 99658 525891
rect 99714 525835 99762 525891
rect 99818 525835 99866 525891
rect 99922 525835 99970 525891
rect 100026 525835 100074 525891
rect 100130 525835 100178 525891
rect 100234 525835 100282 525891
rect 100338 525835 100386 525891
rect 100442 525835 100490 525891
rect 100546 525835 100594 525891
rect 100650 525835 100698 525891
rect 100754 525835 100802 525891
rect 100858 525835 100906 525891
rect 100962 525835 101010 525891
rect 101066 525835 101114 525891
rect 101170 525835 101218 525891
rect 101274 525835 101322 525891
rect 101378 525835 101426 525891
rect 101482 525835 101530 525891
rect 101586 525835 101634 525891
rect 101690 525835 101738 525891
rect 101794 525835 101842 525891
rect 101898 525835 101946 525891
rect 102002 525835 102050 525891
rect 102106 525835 102154 525891
rect 102210 525835 102258 525891
rect 102314 525835 102362 525891
rect 102418 525835 102466 525891
rect 102522 525835 102570 525891
rect 102626 525835 102674 525891
rect 102730 525835 102778 525891
rect 102834 525835 102882 525891
rect 102938 525835 102986 525891
rect 103042 525835 103090 525891
rect 103146 525835 103194 525891
rect 103250 525835 103298 525891
rect 103354 525835 103402 525891
rect 103458 525835 103506 525891
rect 103562 525835 103610 525891
rect 103666 525835 103714 525891
rect 103770 525835 103818 525891
rect 103874 525835 103922 525891
rect 103978 525835 104026 525891
rect 104082 525835 104130 525891
rect 104186 525835 104234 525891
rect 104290 525835 104338 525891
rect 104394 525835 104442 525891
rect 104498 525835 104546 525891
rect 104602 525835 104650 525891
rect 104706 525835 104754 525891
rect 104810 525835 104858 525891
rect 104914 525835 104962 525891
rect 105018 525835 105066 525891
rect 105122 525835 105170 525891
rect 105226 525835 105274 525891
rect 105330 525835 105378 525891
rect 105434 525835 105482 525891
rect 105538 525835 105586 525891
rect 105642 525835 105690 525891
rect 105746 525835 105794 525891
rect 105850 525835 105898 525891
rect 105954 525835 106002 525891
rect 106058 525835 106106 525891
rect 106162 525835 106210 525891
rect 106266 525835 106314 525891
rect 106370 525835 106418 525891
rect 106474 525835 106522 525891
rect 106578 525835 106626 525891
rect 106682 525835 106730 525891
rect 106786 525835 106834 525891
rect 106890 525835 106938 525891
rect 106994 525835 107042 525891
rect 107098 525835 107146 525891
rect 107202 525835 107250 525891
rect 107306 525835 107354 525891
rect 107410 525835 107458 525891
rect 107514 525835 107562 525891
rect 107618 525835 107666 525891
rect 107722 525835 107770 525891
rect 107826 525835 107874 525891
rect 107930 525835 107978 525891
rect 108034 525835 108082 525891
rect 108138 525835 108186 525891
rect 108242 525835 108290 525891
rect 108346 525835 108394 525891
rect 108450 525835 108498 525891
rect 108554 525835 108602 525891
rect 108658 525835 108706 525891
rect 108762 525835 108810 525891
rect 108866 525835 597980 525891
rect -1916 525826 597980 525835
rect -1916 514412 597980 514446
rect -1916 514356 60355 514412
rect 60411 514356 60479 514412
rect 60535 514356 60603 514412
rect 60659 514356 60727 514412
rect 60783 514356 60851 514412
rect 60907 514356 60975 514412
rect 61031 514356 61099 514412
rect 61155 514356 61223 514412
rect 61279 514356 61347 514412
rect 61403 514356 61471 514412
rect 61527 514356 61595 514412
rect 61651 514356 61719 514412
rect 61775 514356 61843 514412
rect 61899 514356 61967 514412
rect 62023 514356 62091 514412
rect 62147 514356 62215 514412
rect 62271 514356 62339 514412
rect 62395 514356 62463 514412
rect 62519 514356 62587 514412
rect 62643 514356 62711 514412
rect 62767 514356 62835 514412
rect 62891 514356 62959 514412
rect 63015 514356 63083 514412
rect 63139 514356 63207 514412
rect 63263 514356 63331 514412
rect 63387 514356 63455 514412
rect 63511 514356 63579 514412
rect 63635 514356 63703 514412
rect 63759 514356 63827 514412
rect 63883 514356 63951 514412
rect 64007 514356 64075 514412
rect 64131 514356 64199 514412
rect 64255 514356 64323 514412
rect 64379 514356 64447 514412
rect 64503 514356 64571 514412
rect 64627 514356 64695 514412
rect 64751 514356 64819 514412
rect 64875 514356 64943 514412
rect 64999 514356 65067 514412
rect 65123 514356 65191 514412
rect 65247 514356 65315 514412
rect 65371 514356 65439 514412
rect 65495 514356 597980 514412
rect -1916 514350 597980 514356
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 9234 514350
rect 9290 514294 9358 514350
rect 9414 514294 9482 514350
rect 9538 514294 9606 514350
rect 9662 514294 39954 514350
rect 40010 514294 40078 514350
rect 40134 514294 40202 514350
rect 40258 514294 40326 514350
rect 40382 514294 162834 514350
rect 162890 514294 162958 514350
rect 163014 514294 163082 514350
rect 163138 514294 163206 514350
rect 163262 514294 209878 514350
rect 209934 514294 210002 514350
rect 210058 514294 240598 514350
rect 240654 514294 240722 514350
rect 240778 514294 271318 514350
rect 271374 514294 271442 514350
rect 271498 514294 302038 514350
rect 302094 514294 302162 514350
rect 302218 514294 332758 514350
rect 332814 514294 332882 514350
rect 332938 514294 363478 514350
rect 363534 514294 363602 514350
rect 363658 514294 394198 514350
rect 394254 514294 394322 514350
rect 394378 514294 424918 514350
rect 424974 514294 425042 514350
rect 425098 514294 455638 514350
rect 455694 514294 455762 514350
rect 455818 514294 486358 514350
rect 486414 514294 486482 514350
rect 486538 514294 517078 514350
rect 517134 514294 517202 514350
rect 517258 514294 547798 514350
rect 547854 514294 547922 514350
rect 547978 514294 562194 514350
rect 562250 514294 562318 514350
rect 562374 514294 562442 514350
rect 562498 514294 562566 514350
rect 562622 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect -1916 514288 597980 514294
rect -1916 514232 60355 514288
rect 60411 514232 60479 514288
rect 60535 514232 60603 514288
rect 60659 514232 60727 514288
rect 60783 514232 60851 514288
rect 60907 514232 60975 514288
rect 61031 514232 61099 514288
rect 61155 514232 61223 514288
rect 61279 514232 61347 514288
rect 61403 514232 61471 514288
rect 61527 514232 61595 514288
rect 61651 514232 61719 514288
rect 61775 514232 61843 514288
rect 61899 514232 61967 514288
rect 62023 514232 62091 514288
rect 62147 514232 62215 514288
rect 62271 514232 62339 514288
rect 62395 514232 62463 514288
rect 62519 514232 62587 514288
rect 62643 514232 62711 514288
rect 62767 514232 62835 514288
rect 62891 514232 62959 514288
rect 63015 514232 63083 514288
rect 63139 514232 63207 514288
rect 63263 514232 63331 514288
rect 63387 514232 63455 514288
rect 63511 514232 63579 514288
rect 63635 514232 63703 514288
rect 63759 514232 63827 514288
rect 63883 514232 63951 514288
rect 64007 514232 64075 514288
rect 64131 514232 64199 514288
rect 64255 514232 64323 514288
rect 64379 514232 64447 514288
rect 64503 514232 64571 514288
rect 64627 514232 64695 514288
rect 64751 514232 64819 514288
rect 64875 514232 64943 514288
rect 64999 514232 65067 514288
rect 65123 514232 65191 514288
rect 65247 514232 65315 514288
rect 65371 514232 65439 514288
rect 65495 514232 597980 514288
rect -1916 514226 597980 514232
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 9234 514226
rect 9290 514170 9358 514226
rect 9414 514170 9482 514226
rect 9538 514170 9606 514226
rect 9662 514170 39954 514226
rect 40010 514170 40078 514226
rect 40134 514170 40202 514226
rect 40258 514170 40326 514226
rect 40382 514170 162834 514226
rect 162890 514170 162958 514226
rect 163014 514170 163082 514226
rect 163138 514170 163206 514226
rect 163262 514170 209878 514226
rect 209934 514170 210002 514226
rect 210058 514170 240598 514226
rect 240654 514170 240722 514226
rect 240778 514170 271318 514226
rect 271374 514170 271442 514226
rect 271498 514170 302038 514226
rect 302094 514170 302162 514226
rect 302218 514170 332758 514226
rect 332814 514170 332882 514226
rect 332938 514170 363478 514226
rect 363534 514170 363602 514226
rect 363658 514170 394198 514226
rect 394254 514170 394322 514226
rect 394378 514170 424918 514226
rect 424974 514170 425042 514226
rect 425098 514170 455638 514226
rect 455694 514170 455762 514226
rect 455818 514170 486358 514226
rect 486414 514170 486482 514226
rect 486538 514170 517078 514226
rect 517134 514170 517202 514226
rect 517258 514170 547798 514226
rect 547854 514170 547922 514226
rect 547978 514170 562194 514226
rect 562250 514170 562318 514226
rect 562374 514170 562442 514226
rect 562498 514170 562566 514226
rect 562622 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect -1916 514164 597980 514170
rect -1916 514108 60355 514164
rect 60411 514108 60479 514164
rect 60535 514108 60603 514164
rect 60659 514108 60727 514164
rect 60783 514108 60851 514164
rect 60907 514108 60975 514164
rect 61031 514108 61099 514164
rect 61155 514108 61223 514164
rect 61279 514108 61347 514164
rect 61403 514108 61471 514164
rect 61527 514108 61595 514164
rect 61651 514108 61719 514164
rect 61775 514108 61843 514164
rect 61899 514108 61967 514164
rect 62023 514108 62091 514164
rect 62147 514108 62215 514164
rect 62271 514108 62339 514164
rect 62395 514108 62463 514164
rect 62519 514108 62587 514164
rect 62643 514108 62711 514164
rect 62767 514108 62835 514164
rect 62891 514108 62959 514164
rect 63015 514108 63083 514164
rect 63139 514108 63207 514164
rect 63263 514108 63331 514164
rect 63387 514108 63455 514164
rect 63511 514108 63579 514164
rect 63635 514108 63703 514164
rect 63759 514108 63827 514164
rect 63883 514108 63951 514164
rect 64007 514108 64075 514164
rect 64131 514108 64199 514164
rect 64255 514108 64323 514164
rect 64379 514108 64447 514164
rect 64503 514108 64571 514164
rect 64627 514108 64695 514164
rect 64751 514108 64819 514164
rect 64875 514108 64943 514164
rect 64999 514108 65067 514164
rect 65123 514108 65191 514164
rect 65247 514108 65315 514164
rect 65371 514108 65439 514164
rect 65495 514108 597980 514164
rect -1916 514102 597980 514108
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 9234 514102
rect 9290 514046 9358 514102
rect 9414 514046 9482 514102
rect 9538 514046 9606 514102
rect 9662 514046 39954 514102
rect 40010 514046 40078 514102
rect 40134 514046 40202 514102
rect 40258 514046 40326 514102
rect 40382 514046 162834 514102
rect 162890 514046 162958 514102
rect 163014 514046 163082 514102
rect 163138 514046 163206 514102
rect 163262 514046 209878 514102
rect 209934 514046 210002 514102
rect 210058 514046 240598 514102
rect 240654 514046 240722 514102
rect 240778 514046 271318 514102
rect 271374 514046 271442 514102
rect 271498 514046 302038 514102
rect 302094 514046 302162 514102
rect 302218 514046 332758 514102
rect 332814 514046 332882 514102
rect 332938 514046 363478 514102
rect 363534 514046 363602 514102
rect 363658 514046 394198 514102
rect 394254 514046 394322 514102
rect 394378 514046 424918 514102
rect 424974 514046 425042 514102
rect 425098 514046 455638 514102
rect 455694 514046 455762 514102
rect 455818 514046 486358 514102
rect 486414 514046 486482 514102
rect 486538 514046 517078 514102
rect 517134 514046 517202 514102
rect 517258 514046 547798 514102
rect 547854 514046 547922 514102
rect 547978 514046 562194 514102
rect 562250 514046 562318 514102
rect 562374 514046 562442 514102
rect 562498 514046 562566 514102
rect 562622 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect -1916 514040 597980 514046
rect -1916 513984 60355 514040
rect 60411 513984 60479 514040
rect 60535 513984 60603 514040
rect 60659 513984 60727 514040
rect 60783 513984 60851 514040
rect 60907 513984 60975 514040
rect 61031 513984 61099 514040
rect 61155 513984 61223 514040
rect 61279 513984 61347 514040
rect 61403 513984 61471 514040
rect 61527 513984 61595 514040
rect 61651 513984 61719 514040
rect 61775 513984 61843 514040
rect 61899 513984 61967 514040
rect 62023 513984 62091 514040
rect 62147 513984 62215 514040
rect 62271 513984 62339 514040
rect 62395 513984 62463 514040
rect 62519 513984 62587 514040
rect 62643 513984 62711 514040
rect 62767 513984 62835 514040
rect 62891 513984 62959 514040
rect 63015 513984 63083 514040
rect 63139 513984 63207 514040
rect 63263 513984 63331 514040
rect 63387 513984 63455 514040
rect 63511 513984 63579 514040
rect 63635 513984 63703 514040
rect 63759 513984 63827 514040
rect 63883 513984 63951 514040
rect 64007 513984 64075 514040
rect 64131 513984 64199 514040
rect 64255 513984 64323 514040
rect 64379 513984 64447 514040
rect 64503 513984 64571 514040
rect 64627 513984 64695 514040
rect 64751 513984 64819 514040
rect 64875 513984 64943 514040
rect 64999 513984 65067 514040
rect 65123 513984 65191 514040
rect 65247 513984 65315 514040
rect 65371 513984 65439 514040
rect 65495 513984 597980 514040
rect -1916 513978 597980 513984
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 9234 513978
rect 9290 513922 9358 513978
rect 9414 513922 9482 513978
rect 9538 513922 9606 513978
rect 9662 513922 39954 513978
rect 40010 513922 40078 513978
rect 40134 513922 40202 513978
rect 40258 513922 40326 513978
rect 40382 513922 162834 513978
rect 162890 513922 162958 513978
rect 163014 513922 163082 513978
rect 163138 513922 163206 513978
rect 163262 513922 209878 513978
rect 209934 513922 210002 513978
rect 210058 513922 240598 513978
rect 240654 513922 240722 513978
rect 240778 513922 271318 513978
rect 271374 513922 271442 513978
rect 271498 513922 302038 513978
rect 302094 513922 302162 513978
rect 302218 513922 332758 513978
rect 332814 513922 332882 513978
rect 332938 513922 363478 513978
rect 363534 513922 363602 513978
rect 363658 513922 394198 513978
rect 394254 513922 394322 513978
rect 394378 513922 424918 513978
rect 424974 513922 425042 513978
rect 425098 513922 455638 513978
rect 455694 513922 455762 513978
rect 455818 513922 486358 513978
rect 486414 513922 486482 513978
rect 486538 513922 517078 513978
rect 517134 513922 517202 513978
rect 517258 513922 547798 513978
rect 547854 513922 547922 513978
rect 547978 513922 562194 513978
rect 562250 513922 562318 513978
rect 562374 513922 562442 513978
rect 562498 513922 562566 513978
rect 562622 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect -1916 513916 597980 513922
rect -1916 513860 60355 513916
rect 60411 513860 60479 513916
rect 60535 513860 60603 513916
rect 60659 513860 60727 513916
rect 60783 513860 60851 513916
rect 60907 513860 60975 513916
rect 61031 513860 61099 513916
rect 61155 513860 61223 513916
rect 61279 513860 61347 513916
rect 61403 513860 61471 513916
rect 61527 513860 61595 513916
rect 61651 513860 61719 513916
rect 61775 513860 61843 513916
rect 61899 513860 61967 513916
rect 62023 513860 62091 513916
rect 62147 513860 62215 513916
rect 62271 513860 62339 513916
rect 62395 513860 62463 513916
rect 62519 513860 62587 513916
rect 62643 513860 62711 513916
rect 62767 513860 62835 513916
rect 62891 513860 62959 513916
rect 63015 513860 63083 513916
rect 63139 513860 63207 513916
rect 63263 513860 63331 513916
rect 63387 513860 63455 513916
rect 63511 513860 63579 513916
rect 63635 513860 63703 513916
rect 63759 513860 63827 513916
rect 63883 513860 63951 513916
rect 64007 513860 64075 513916
rect 64131 513860 64199 513916
rect 64255 513860 64323 513916
rect 64379 513860 64447 513916
rect 64503 513860 64571 513916
rect 64627 513860 64695 513916
rect 64751 513860 64819 513916
rect 64875 513860 64943 513916
rect 64999 513860 65067 513916
rect 65123 513860 65191 513916
rect 65247 513860 65315 513916
rect 65371 513860 65439 513916
rect 65495 513860 597980 513916
rect -1916 513826 597980 513860
rect -1916 508350 597980 508446
rect -1916 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 36234 508350
rect 36290 508294 36358 508350
rect 36414 508294 36482 508350
rect 36538 508294 36606 508350
rect 36662 508294 159114 508350
rect 159170 508294 159238 508350
rect 159294 508294 159362 508350
rect 159418 508294 159486 508350
rect 159542 508294 189834 508350
rect 189890 508294 189958 508350
rect 190014 508294 190082 508350
rect 190138 508294 190206 508350
rect 190262 508294 194518 508350
rect 194574 508294 194642 508350
rect 194698 508294 225238 508350
rect 225294 508294 225362 508350
rect 225418 508294 255958 508350
rect 256014 508294 256082 508350
rect 256138 508294 286678 508350
rect 286734 508294 286802 508350
rect 286858 508294 317398 508350
rect 317454 508294 317522 508350
rect 317578 508294 348118 508350
rect 348174 508294 348242 508350
rect 348298 508294 378838 508350
rect 378894 508294 378962 508350
rect 379018 508294 409558 508350
rect 409614 508294 409682 508350
rect 409738 508294 440278 508350
rect 440334 508294 440402 508350
rect 440458 508294 470998 508350
rect 471054 508294 471122 508350
rect 471178 508294 501718 508350
rect 501774 508294 501842 508350
rect 501898 508294 532438 508350
rect 532494 508294 532562 508350
rect 532618 508294 558474 508350
rect 558530 508294 558598 508350
rect 558654 508294 558722 508350
rect 558778 508294 558846 508350
rect 558902 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597980 508350
rect -1916 508290 597980 508294
rect -1916 508234 85231 508290
rect 85287 508234 85355 508290
rect 85411 508234 85479 508290
rect 85535 508234 85603 508290
rect 85659 508234 85727 508290
rect 85783 508234 85851 508290
rect 85907 508234 85975 508290
rect 86031 508234 86099 508290
rect 86155 508234 86223 508290
rect 86279 508234 86347 508290
rect 86403 508234 86471 508290
rect 86527 508234 86595 508290
rect 86651 508234 86719 508290
rect 86775 508234 86843 508290
rect 86899 508234 86967 508290
rect 87023 508234 87091 508290
rect 87147 508234 87215 508290
rect 87271 508234 87339 508290
rect 87395 508234 87463 508290
rect 87519 508234 87587 508290
rect 87643 508234 87711 508290
rect 87767 508234 87835 508290
rect 87891 508234 87959 508290
rect 88015 508234 88083 508290
rect 88139 508234 88207 508290
rect 88263 508234 88331 508290
rect 88387 508234 88455 508290
rect 88511 508234 88579 508290
rect 88635 508234 88703 508290
rect 88759 508234 88827 508290
rect 88883 508234 88951 508290
rect 89007 508234 89075 508290
rect 89131 508234 89199 508290
rect 89255 508234 89323 508290
rect 89379 508234 89447 508290
rect 89503 508234 89571 508290
rect 89627 508234 89695 508290
rect 89751 508234 89819 508290
rect 89875 508234 89943 508290
rect 89999 508234 90067 508290
rect 90123 508234 90191 508290
rect 90247 508234 90315 508290
rect 90371 508234 90439 508290
rect 90495 508234 90563 508290
rect 90619 508234 90687 508290
rect 90743 508234 90811 508290
rect 90867 508234 90935 508290
rect 90991 508234 91059 508290
rect 91115 508234 91183 508290
rect 91239 508234 91307 508290
rect 91363 508234 91431 508290
rect 91487 508234 91555 508290
rect 91611 508234 91679 508290
rect 91735 508234 91803 508290
rect 91859 508234 91927 508290
rect 91983 508234 92051 508290
rect 92107 508234 92175 508290
rect 92231 508234 92299 508290
rect 92355 508234 92423 508290
rect 92479 508234 92547 508290
rect 92603 508234 92671 508290
rect 92727 508234 92795 508290
rect 92851 508234 92919 508290
rect 92975 508234 93043 508290
rect 93099 508234 93167 508290
rect 93223 508234 93291 508290
rect 93347 508234 93415 508290
rect 93471 508234 93539 508290
rect 93595 508234 93663 508290
rect 93719 508234 597980 508290
rect -1916 508226 597980 508234
rect -1916 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 36234 508226
rect 36290 508170 36358 508226
rect 36414 508170 36482 508226
rect 36538 508170 36606 508226
rect 36662 508170 159114 508226
rect 159170 508170 159238 508226
rect 159294 508170 159362 508226
rect 159418 508170 159486 508226
rect 159542 508170 189834 508226
rect 189890 508170 189958 508226
rect 190014 508170 190082 508226
rect 190138 508170 190206 508226
rect 190262 508170 194518 508226
rect 194574 508170 194642 508226
rect 194698 508170 225238 508226
rect 225294 508170 225362 508226
rect 225418 508170 255958 508226
rect 256014 508170 256082 508226
rect 256138 508170 286678 508226
rect 286734 508170 286802 508226
rect 286858 508170 317398 508226
rect 317454 508170 317522 508226
rect 317578 508170 348118 508226
rect 348174 508170 348242 508226
rect 348298 508170 378838 508226
rect 378894 508170 378962 508226
rect 379018 508170 409558 508226
rect 409614 508170 409682 508226
rect 409738 508170 440278 508226
rect 440334 508170 440402 508226
rect 440458 508170 470998 508226
rect 471054 508170 471122 508226
rect 471178 508170 501718 508226
rect 501774 508170 501842 508226
rect 501898 508170 532438 508226
rect 532494 508170 532562 508226
rect 532618 508170 558474 508226
rect 558530 508170 558598 508226
rect 558654 508170 558722 508226
rect 558778 508170 558846 508226
rect 558902 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597980 508226
rect -1916 508166 597980 508170
rect -1916 508110 85231 508166
rect 85287 508110 85355 508166
rect 85411 508110 85479 508166
rect 85535 508110 85603 508166
rect 85659 508110 85727 508166
rect 85783 508110 85851 508166
rect 85907 508110 85975 508166
rect 86031 508110 86099 508166
rect 86155 508110 86223 508166
rect 86279 508110 86347 508166
rect 86403 508110 86471 508166
rect 86527 508110 86595 508166
rect 86651 508110 86719 508166
rect 86775 508110 86843 508166
rect 86899 508110 86967 508166
rect 87023 508110 87091 508166
rect 87147 508110 87215 508166
rect 87271 508110 87339 508166
rect 87395 508110 87463 508166
rect 87519 508110 87587 508166
rect 87643 508110 87711 508166
rect 87767 508110 87835 508166
rect 87891 508110 87959 508166
rect 88015 508110 88083 508166
rect 88139 508110 88207 508166
rect 88263 508110 88331 508166
rect 88387 508110 88455 508166
rect 88511 508110 88579 508166
rect 88635 508110 88703 508166
rect 88759 508110 88827 508166
rect 88883 508110 88951 508166
rect 89007 508110 89075 508166
rect 89131 508110 89199 508166
rect 89255 508110 89323 508166
rect 89379 508110 89447 508166
rect 89503 508110 89571 508166
rect 89627 508110 89695 508166
rect 89751 508110 89819 508166
rect 89875 508110 89943 508166
rect 89999 508110 90067 508166
rect 90123 508110 90191 508166
rect 90247 508110 90315 508166
rect 90371 508110 90439 508166
rect 90495 508110 90563 508166
rect 90619 508110 90687 508166
rect 90743 508110 90811 508166
rect 90867 508110 90935 508166
rect 90991 508110 91059 508166
rect 91115 508110 91183 508166
rect 91239 508110 91307 508166
rect 91363 508110 91431 508166
rect 91487 508110 91555 508166
rect 91611 508110 91679 508166
rect 91735 508110 91803 508166
rect 91859 508110 91927 508166
rect 91983 508110 92051 508166
rect 92107 508110 92175 508166
rect 92231 508110 92299 508166
rect 92355 508110 92423 508166
rect 92479 508110 92547 508166
rect 92603 508110 92671 508166
rect 92727 508110 92795 508166
rect 92851 508110 92919 508166
rect 92975 508110 93043 508166
rect 93099 508110 93167 508166
rect 93223 508110 93291 508166
rect 93347 508110 93415 508166
rect 93471 508110 93539 508166
rect 93595 508110 93663 508166
rect 93719 508110 597980 508166
rect -1916 508102 597980 508110
rect -1916 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 36234 508102
rect 36290 508046 36358 508102
rect 36414 508046 36482 508102
rect 36538 508046 36606 508102
rect 36662 508046 159114 508102
rect 159170 508046 159238 508102
rect 159294 508046 159362 508102
rect 159418 508046 159486 508102
rect 159542 508046 189834 508102
rect 189890 508046 189958 508102
rect 190014 508046 190082 508102
rect 190138 508046 190206 508102
rect 190262 508046 194518 508102
rect 194574 508046 194642 508102
rect 194698 508046 225238 508102
rect 225294 508046 225362 508102
rect 225418 508046 255958 508102
rect 256014 508046 256082 508102
rect 256138 508046 286678 508102
rect 286734 508046 286802 508102
rect 286858 508046 317398 508102
rect 317454 508046 317522 508102
rect 317578 508046 348118 508102
rect 348174 508046 348242 508102
rect 348298 508046 378838 508102
rect 378894 508046 378962 508102
rect 379018 508046 409558 508102
rect 409614 508046 409682 508102
rect 409738 508046 440278 508102
rect 440334 508046 440402 508102
rect 440458 508046 470998 508102
rect 471054 508046 471122 508102
rect 471178 508046 501718 508102
rect 501774 508046 501842 508102
rect 501898 508046 532438 508102
rect 532494 508046 532562 508102
rect 532618 508046 558474 508102
rect 558530 508046 558598 508102
rect 558654 508046 558722 508102
rect 558778 508046 558846 508102
rect 558902 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597980 508102
rect -1916 507978 597980 508046
rect -1916 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 36234 507978
rect 36290 507922 36358 507978
rect 36414 507922 36482 507978
rect 36538 507922 36606 507978
rect 36662 507922 159114 507978
rect 159170 507922 159238 507978
rect 159294 507922 159362 507978
rect 159418 507922 159486 507978
rect 159542 507922 189834 507978
rect 189890 507922 189958 507978
rect 190014 507922 190082 507978
rect 190138 507922 190206 507978
rect 190262 507922 194518 507978
rect 194574 507922 194642 507978
rect 194698 507922 225238 507978
rect 225294 507922 225362 507978
rect 225418 507922 255958 507978
rect 256014 507922 256082 507978
rect 256138 507922 286678 507978
rect 286734 507922 286802 507978
rect 286858 507922 317398 507978
rect 317454 507922 317522 507978
rect 317578 507922 348118 507978
rect 348174 507922 348242 507978
rect 348298 507922 378838 507978
rect 378894 507922 378962 507978
rect 379018 507922 409558 507978
rect 409614 507922 409682 507978
rect 409738 507922 440278 507978
rect 440334 507922 440402 507978
rect 440458 507922 470998 507978
rect 471054 507922 471122 507978
rect 471178 507922 501718 507978
rect 501774 507922 501842 507978
rect 501898 507922 532438 507978
rect 532494 507922 532562 507978
rect 532618 507922 558474 507978
rect 558530 507922 558598 507978
rect 558654 507922 558722 507978
rect 558778 507922 558846 507978
rect 558902 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597980 507978
rect -1916 507891 597980 507922
rect -1916 507835 85062 507891
rect 85118 507835 85166 507891
rect 85222 507835 85270 507891
rect 85326 507835 85374 507891
rect 85430 507835 85478 507891
rect 85534 507835 85582 507891
rect 85638 507835 85686 507891
rect 85742 507835 85790 507891
rect 85846 507835 85894 507891
rect 85950 507835 85998 507891
rect 86054 507835 86102 507891
rect 86158 507835 86206 507891
rect 86262 507835 86310 507891
rect 86366 507835 86414 507891
rect 86470 507835 86518 507891
rect 86574 507835 86622 507891
rect 86678 507835 86726 507891
rect 86782 507835 86830 507891
rect 86886 507835 86934 507891
rect 86990 507835 87038 507891
rect 87094 507835 87142 507891
rect 87198 507835 87246 507891
rect 87302 507835 87350 507891
rect 87406 507835 87454 507891
rect 87510 507835 87558 507891
rect 87614 507835 87662 507891
rect 87718 507835 87766 507891
rect 87822 507835 87870 507891
rect 87926 507835 87974 507891
rect 88030 507835 88078 507891
rect 88134 507835 88182 507891
rect 88238 507835 88286 507891
rect 88342 507835 88390 507891
rect 88446 507835 88494 507891
rect 88550 507835 88598 507891
rect 88654 507835 88702 507891
rect 88758 507835 88806 507891
rect 88862 507835 88910 507891
rect 88966 507835 89014 507891
rect 89070 507835 89118 507891
rect 89174 507835 89222 507891
rect 89278 507835 89326 507891
rect 89382 507835 89430 507891
rect 89486 507835 89534 507891
rect 89590 507835 89638 507891
rect 89694 507835 89742 507891
rect 89798 507835 89846 507891
rect 89902 507835 89950 507891
rect 90006 507835 90054 507891
rect 90110 507835 90158 507891
rect 90214 507835 90262 507891
rect 90318 507835 90366 507891
rect 90422 507835 90470 507891
rect 90526 507835 90574 507891
rect 90630 507835 90678 507891
rect 90734 507835 90782 507891
rect 90838 507835 90886 507891
rect 90942 507835 90990 507891
rect 91046 507835 91094 507891
rect 91150 507835 91198 507891
rect 91254 507835 91302 507891
rect 91358 507835 91406 507891
rect 91462 507835 91510 507891
rect 91566 507835 91614 507891
rect 91670 507835 91718 507891
rect 91774 507835 91822 507891
rect 91878 507835 91926 507891
rect 91982 507835 92030 507891
rect 92086 507835 92134 507891
rect 92190 507835 92238 507891
rect 92294 507835 92342 507891
rect 92398 507835 92446 507891
rect 92502 507835 92550 507891
rect 92606 507835 92654 507891
rect 92710 507835 92758 507891
rect 92814 507835 92862 507891
rect 92918 507835 92966 507891
rect 93022 507835 93070 507891
rect 93126 507835 93174 507891
rect 93230 507835 93278 507891
rect 93334 507835 93382 507891
rect 93438 507835 597980 507891
rect -1916 507826 597980 507835
rect -1916 496413 597980 496446
rect -1916 496357 63508 496413
rect 63564 496357 63632 496413
rect 63688 496357 63756 496413
rect 63812 496357 63880 496413
rect 63936 496357 64004 496413
rect 64060 496357 64128 496413
rect 64184 496357 64252 496413
rect 64308 496357 64376 496413
rect 64432 496357 64500 496413
rect 64556 496357 64624 496413
rect 64680 496357 64748 496413
rect 64804 496357 64872 496413
rect 64928 496357 64996 496413
rect 65052 496357 65120 496413
rect 65176 496357 65244 496413
rect 65300 496357 65368 496413
rect 65424 496357 65492 496413
rect 65548 496357 65616 496413
rect 65672 496357 65740 496413
rect 65796 496357 65864 496413
rect 65920 496357 65988 496413
rect 66044 496357 66112 496413
rect 66168 496357 66236 496413
rect 66292 496357 66360 496413
rect 66416 496357 66484 496413
rect 66540 496357 66608 496413
rect 66664 496357 66732 496413
rect 66788 496357 66856 496413
rect 66912 496357 66980 496413
rect 67036 496357 67104 496413
rect 67160 496357 67228 496413
rect 67284 496357 67352 496413
rect 67408 496357 67476 496413
rect 67532 496357 67600 496413
rect 67656 496357 67724 496413
rect 67780 496357 67848 496413
rect 67904 496357 67972 496413
rect 68028 496357 68096 496413
rect 68152 496357 68220 496413
rect 68276 496357 68344 496413
rect 68400 496357 68468 496413
rect 68524 496357 68592 496413
rect 68648 496357 68716 496413
rect 68772 496357 68840 496413
rect 68896 496357 68964 496413
rect 69020 496357 69088 496413
rect 69144 496357 69212 496413
rect 69268 496357 69336 496413
rect 69392 496357 597980 496413
rect -1916 496350 597980 496357
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 9234 496350
rect 9290 496294 9358 496350
rect 9414 496294 9482 496350
rect 9538 496294 9606 496350
rect 9662 496294 39954 496350
rect 40010 496294 40078 496350
rect 40134 496294 40202 496350
rect 40258 496294 40326 496350
rect 40382 496294 132114 496350
rect 132170 496294 132238 496350
rect 132294 496294 132362 496350
rect 132418 496294 132486 496350
rect 132542 496294 162834 496350
rect 162890 496294 162958 496350
rect 163014 496294 163082 496350
rect 163138 496294 163206 496350
rect 163262 496294 209878 496350
rect 209934 496294 210002 496350
rect 210058 496294 240598 496350
rect 240654 496294 240722 496350
rect 240778 496294 271318 496350
rect 271374 496294 271442 496350
rect 271498 496294 302038 496350
rect 302094 496294 302162 496350
rect 302218 496294 332758 496350
rect 332814 496294 332882 496350
rect 332938 496294 363478 496350
rect 363534 496294 363602 496350
rect 363658 496294 394198 496350
rect 394254 496294 394322 496350
rect 394378 496294 424918 496350
rect 424974 496294 425042 496350
rect 425098 496294 455638 496350
rect 455694 496294 455762 496350
rect 455818 496294 486358 496350
rect 486414 496294 486482 496350
rect 486538 496294 517078 496350
rect 517134 496294 517202 496350
rect 517258 496294 547798 496350
rect 547854 496294 547922 496350
rect 547978 496294 562194 496350
rect 562250 496294 562318 496350
rect 562374 496294 562442 496350
rect 562498 496294 562566 496350
rect 562622 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect -1916 496289 597980 496294
rect -1916 496233 63508 496289
rect 63564 496233 63632 496289
rect 63688 496233 63756 496289
rect 63812 496233 63880 496289
rect 63936 496233 64004 496289
rect 64060 496233 64128 496289
rect 64184 496233 64252 496289
rect 64308 496233 64376 496289
rect 64432 496233 64500 496289
rect 64556 496233 64624 496289
rect 64680 496233 64748 496289
rect 64804 496233 64872 496289
rect 64928 496233 64996 496289
rect 65052 496233 65120 496289
rect 65176 496233 65244 496289
rect 65300 496233 65368 496289
rect 65424 496233 65492 496289
rect 65548 496233 65616 496289
rect 65672 496233 65740 496289
rect 65796 496233 65864 496289
rect 65920 496233 65988 496289
rect 66044 496233 66112 496289
rect 66168 496233 66236 496289
rect 66292 496233 66360 496289
rect 66416 496233 66484 496289
rect 66540 496233 66608 496289
rect 66664 496233 66732 496289
rect 66788 496233 66856 496289
rect 66912 496233 66980 496289
rect 67036 496233 67104 496289
rect 67160 496233 67228 496289
rect 67284 496233 67352 496289
rect 67408 496233 67476 496289
rect 67532 496233 67600 496289
rect 67656 496233 67724 496289
rect 67780 496233 67848 496289
rect 67904 496233 67972 496289
rect 68028 496233 68096 496289
rect 68152 496233 68220 496289
rect 68276 496233 68344 496289
rect 68400 496233 68468 496289
rect 68524 496233 68592 496289
rect 68648 496233 68716 496289
rect 68772 496233 68840 496289
rect 68896 496233 68964 496289
rect 69020 496233 69088 496289
rect 69144 496233 69212 496289
rect 69268 496233 69336 496289
rect 69392 496233 597980 496289
rect -1916 496226 597980 496233
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 9234 496226
rect 9290 496170 9358 496226
rect 9414 496170 9482 496226
rect 9538 496170 9606 496226
rect 9662 496170 39954 496226
rect 40010 496170 40078 496226
rect 40134 496170 40202 496226
rect 40258 496170 40326 496226
rect 40382 496170 132114 496226
rect 132170 496170 132238 496226
rect 132294 496170 132362 496226
rect 132418 496170 132486 496226
rect 132542 496170 162834 496226
rect 162890 496170 162958 496226
rect 163014 496170 163082 496226
rect 163138 496170 163206 496226
rect 163262 496170 209878 496226
rect 209934 496170 210002 496226
rect 210058 496170 240598 496226
rect 240654 496170 240722 496226
rect 240778 496170 271318 496226
rect 271374 496170 271442 496226
rect 271498 496170 302038 496226
rect 302094 496170 302162 496226
rect 302218 496170 332758 496226
rect 332814 496170 332882 496226
rect 332938 496170 363478 496226
rect 363534 496170 363602 496226
rect 363658 496170 394198 496226
rect 394254 496170 394322 496226
rect 394378 496170 424918 496226
rect 424974 496170 425042 496226
rect 425098 496170 455638 496226
rect 455694 496170 455762 496226
rect 455818 496170 486358 496226
rect 486414 496170 486482 496226
rect 486538 496170 517078 496226
rect 517134 496170 517202 496226
rect 517258 496170 547798 496226
rect 547854 496170 547922 496226
rect 547978 496170 562194 496226
rect 562250 496170 562318 496226
rect 562374 496170 562442 496226
rect 562498 496170 562566 496226
rect 562622 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect -1916 496102 597980 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 9234 496102
rect 9290 496046 9358 496102
rect 9414 496046 9482 496102
rect 9538 496046 9606 496102
rect 9662 496046 39954 496102
rect 40010 496046 40078 496102
rect 40134 496046 40202 496102
rect 40258 496046 40326 496102
rect 40382 496046 132114 496102
rect 132170 496046 132238 496102
rect 132294 496046 132362 496102
rect 132418 496046 132486 496102
rect 132542 496046 162834 496102
rect 162890 496046 162958 496102
rect 163014 496046 163082 496102
rect 163138 496046 163206 496102
rect 163262 496046 209878 496102
rect 209934 496046 210002 496102
rect 210058 496046 240598 496102
rect 240654 496046 240722 496102
rect 240778 496046 271318 496102
rect 271374 496046 271442 496102
rect 271498 496046 302038 496102
rect 302094 496046 302162 496102
rect 302218 496046 332758 496102
rect 332814 496046 332882 496102
rect 332938 496046 363478 496102
rect 363534 496046 363602 496102
rect 363658 496046 394198 496102
rect 394254 496046 394322 496102
rect 394378 496046 424918 496102
rect 424974 496046 425042 496102
rect 425098 496046 455638 496102
rect 455694 496046 455762 496102
rect 455818 496046 486358 496102
rect 486414 496046 486482 496102
rect 486538 496046 517078 496102
rect 517134 496046 517202 496102
rect 517258 496046 547798 496102
rect 547854 496046 547922 496102
rect 547978 496046 562194 496102
rect 562250 496046 562318 496102
rect 562374 496046 562442 496102
rect 562498 496046 562566 496102
rect 562622 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect -1916 496003 597980 496046
rect -1916 495978 63671 496003
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 9234 495978
rect 9290 495922 9358 495978
rect 9414 495922 9482 495978
rect 9538 495922 9606 495978
rect 9662 495922 39954 495978
rect 40010 495922 40078 495978
rect 40134 495922 40202 495978
rect 40258 495922 40326 495978
rect 40382 495947 63671 495978
rect 63727 495947 63795 496003
rect 63851 495947 63919 496003
rect 63975 495947 64043 496003
rect 64099 495947 64167 496003
rect 64223 495947 64291 496003
rect 64347 495947 64415 496003
rect 64471 495947 64539 496003
rect 64595 495947 64663 496003
rect 64719 495947 64787 496003
rect 64843 495947 64911 496003
rect 64967 495947 65035 496003
rect 65091 495947 65159 496003
rect 65215 495947 65283 496003
rect 65339 495947 65407 496003
rect 65463 495947 65531 496003
rect 65587 495947 65655 496003
rect 65711 495947 65779 496003
rect 65835 495947 65903 496003
rect 65959 495947 66027 496003
rect 66083 495947 66151 496003
rect 66207 495947 66275 496003
rect 66331 495947 66399 496003
rect 66455 495947 66523 496003
rect 66579 495947 66647 496003
rect 66703 495947 66771 496003
rect 66827 495947 66895 496003
rect 66951 495947 67019 496003
rect 67075 495947 67143 496003
rect 67199 495947 67267 496003
rect 67323 495947 67391 496003
rect 67447 495947 67515 496003
rect 67571 495947 67639 496003
rect 67695 495947 67763 496003
rect 67819 495947 67887 496003
rect 67943 495947 68011 496003
rect 68067 495947 68135 496003
rect 68191 495947 68259 496003
rect 68315 495947 68383 496003
rect 68439 495947 68507 496003
rect 68563 495947 68631 496003
rect 68687 495947 68755 496003
rect 68811 495947 68879 496003
rect 68935 495947 69003 496003
rect 69059 495947 69127 496003
rect 69183 495947 69251 496003
rect 69307 495947 69375 496003
rect 69431 495947 69499 496003
rect 69555 495947 69623 496003
rect 69679 495978 597980 496003
rect 69679 495947 132114 495978
rect 40382 495922 132114 495947
rect 132170 495922 132238 495978
rect 132294 495922 132362 495978
rect 132418 495922 132486 495978
rect 132542 495922 162834 495978
rect 162890 495922 162958 495978
rect 163014 495922 163082 495978
rect 163138 495922 163206 495978
rect 163262 495922 209878 495978
rect 209934 495922 210002 495978
rect 210058 495922 240598 495978
rect 240654 495922 240722 495978
rect 240778 495922 271318 495978
rect 271374 495922 271442 495978
rect 271498 495922 302038 495978
rect 302094 495922 302162 495978
rect 302218 495922 332758 495978
rect 332814 495922 332882 495978
rect 332938 495922 363478 495978
rect 363534 495922 363602 495978
rect 363658 495922 394198 495978
rect 394254 495922 394322 495978
rect 394378 495922 424918 495978
rect 424974 495922 425042 495978
rect 425098 495922 455638 495978
rect 455694 495922 455762 495978
rect 455818 495922 486358 495978
rect 486414 495922 486482 495978
rect 486538 495922 517078 495978
rect 517134 495922 517202 495978
rect 517258 495922 547798 495978
rect 547854 495922 547922 495978
rect 547978 495922 562194 495978
rect 562250 495922 562318 495978
rect 562374 495922 562442 495978
rect 562498 495922 562566 495978
rect 562622 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect -1916 495826 597980 495922
rect -1916 490350 597980 490446
rect -1916 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 36234 490350
rect 36290 490294 36358 490350
rect 36414 490294 36482 490350
rect 36538 490294 36606 490350
rect 36662 490294 128394 490350
rect 128450 490294 128518 490350
rect 128574 490294 128642 490350
rect 128698 490294 128766 490350
rect 128822 490294 159114 490350
rect 159170 490294 159238 490350
rect 159294 490294 159362 490350
rect 159418 490294 159486 490350
rect 159542 490294 189834 490350
rect 189890 490294 189958 490350
rect 190014 490294 190082 490350
rect 190138 490294 190206 490350
rect 190262 490294 194518 490350
rect 194574 490294 194642 490350
rect 194698 490294 225238 490350
rect 225294 490294 225362 490350
rect 225418 490294 255958 490350
rect 256014 490294 256082 490350
rect 256138 490294 286678 490350
rect 286734 490294 286802 490350
rect 286858 490294 317398 490350
rect 317454 490294 317522 490350
rect 317578 490294 348118 490350
rect 348174 490294 348242 490350
rect 348298 490294 378838 490350
rect 378894 490294 378962 490350
rect 379018 490294 409558 490350
rect 409614 490294 409682 490350
rect 409738 490294 440278 490350
rect 440334 490294 440402 490350
rect 440458 490294 470998 490350
rect 471054 490294 471122 490350
rect 471178 490294 501718 490350
rect 501774 490294 501842 490350
rect 501898 490294 532438 490350
rect 532494 490294 532562 490350
rect 532618 490294 558474 490350
rect 558530 490294 558598 490350
rect 558654 490294 558722 490350
rect 558778 490294 558846 490350
rect 558902 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597980 490350
rect -1916 490290 597980 490294
rect -1916 490234 80593 490290
rect 80649 490234 80717 490290
rect 80773 490234 80841 490290
rect 80897 490234 80965 490290
rect 81021 490234 81089 490290
rect 81145 490234 81213 490290
rect 81269 490234 81337 490290
rect 81393 490234 81461 490290
rect 81517 490234 81585 490290
rect 81641 490234 81709 490290
rect 81765 490234 81833 490290
rect 81889 490234 81957 490290
rect 82013 490234 82081 490290
rect 82137 490234 82205 490290
rect 82261 490234 82329 490290
rect 82385 490234 82453 490290
rect 82509 490234 82577 490290
rect 82633 490234 82701 490290
rect 82757 490234 597980 490290
rect -1916 490226 597980 490234
rect -1916 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 36234 490226
rect 36290 490170 36358 490226
rect 36414 490170 36482 490226
rect 36538 490170 36606 490226
rect 36662 490170 128394 490226
rect 128450 490170 128518 490226
rect 128574 490170 128642 490226
rect 128698 490170 128766 490226
rect 128822 490170 159114 490226
rect 159170 490170 159238 490226
rect 159294 490170 159362 490226
rect 159418 490170 159486 490226
rect 159542 490170 189834 490226
rect 189890 490170 189958 490226
rect 190014 490170 190082 490226
rect 190138 490170 190206 490226
rect 190262 490170 194518 490226
rect 194574 490170 194642 490226
rect 194698 490170 225238 490226
rect 225294 490170 225362 490226
rect 225418 490170 255958 490226
rect 256014 490170 256082 490226
rect 256138 490170 286678 490226
rect 286734 490170 286802 490226
rect 286858 490170 317398 490226
rect 317454 490170 317522 490226
rect 317578 490170 348118 490226
rect 348174 490170 348242 490226
rect 348298 490170 378838 490226
rect 378894 490170 378962 490226
rect 379018 490170 409558 490226
rect 409614 490170 409682 490226
rect 409738 490170 440278 490226
rect 440334 490170 440402 490226
rect 440458 490170 470998 490226
rect 471054 490170 471122 490226
rect 471178 490170 501718 490226
rect 501774 490170 501842 490226
rect 501898 490170 532438 490226
rect 532494 490170 532562 490226
rect 532618 490170 558474 490226
rect 558530 490170 558598 490226
rect 558654 490170 558722 490226
rect 558778 490170 558846 490226
rect 558902 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597980 490226
rect -1916 490166 597980 490170
rect -1916 490110 80593 490166
rect 80649 490110 80717 490166
rect 80773 490110 80841 490166
rect 80897 490110 80965 490166
rect 81021 490110 81089 490166
rect 81145 490110 81213 490166
rect 81269 490110 81337 490166
rect 81393 490110 81461 490166
rect 81517 490110 81585 490166
rect 81641 490110 81709 490166
rect 81765 490110 81833 490166
rect 81889 490110 81957 490166
rect 82013 490110 82081 490166
rect 82137 490110 82205 490166
rect 82261 490110 82329 490166
rect 82385 490110 82453 490166
rect 82509 490110 82577 490166
rect 82633 490110 82701 490166
rect 82757 490110 597980 490166
rect -1916 490102 597980 490110
rect -1916 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 36234 490102
rect 36290 490046 36358 490102
rect 36414 490046 36482 490102
rect 36538 490046 36606 490102
rect 36662 490046 128394 490102
rect 128450 490046 128518 490102
rect 128574 490046 128642 490102
rect 128698 490046 128766 490102
rect 128822 490046 159114 490102
rect 159170 490046 159238 490102
rect 159294 490046 159362 490102
rect 159418 490046 159486 490102
rect 159542 490046 189834 490102
rect 189890 490046 189958 490102
rect 190014 490046 190082 490102
rect 190138 490046 190206 490102
rect 190262 490046 194518 490102
rect 194574 490046 194642 490102
rect 194698 490046 225238 490102
rect 225294 490046 225362 490102
rect 225418 490046 255958 490102
rect 256014 490046 256082 490102
rect 256138 490046 286678 490102
rect 286734 490046 286802 490102
rect 286858 490046 317398 490102
rect 317454 490046 317522 490102
rect 317578 490046 348118 490102
rect 348174 490046 348242 490102
rect 348298 490046 378838 490102
rect 378894 490046 378962 490102
rect 379018 490046 409558 490102
rect 409614 490046 409682 490102
rect 409738 490046 440278 490102
rect 440334 490046 440402 490102
rect 440458 490046 470998 490102
rect 471054 490046 471122 490102
rect 471178 490046 501718 490102
rect 501774 490046 501842 490102
rect 501898 490046 532438 490102
rect 532494 490046 532562 490102
rect 532618 490046 558474 490102
rect 558530 490046 558598 490102
rect 558654 490046 558722 490102
rect 558778 490046 558846 490102
rect 558902 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597980 490102
rect -1916 489978 597980 490046
rect -1916 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 36234 489978
rect 36290 489922 36358 489978
rect 36414 489922 36482 489978
rect 36538 489922 36606 489978
rect 36662 489922 128394 489978
rect 128450 489922 128518 489978
rect 128574 489922 128642 489978
rect 128698 489922 128766 489978
rect 128822 489922 159114 489978
rect 159170 489922 159238 489978
rect 159294 489922 159362 489978
rect 159418 489922 159486 489978
rect 159542 489922 189834 489978
rect 189890 489922 189958 489978
rect 190014 489922 190082 489978
rect 190138 489922 190206 489978
rect 190262 489922 194518 489978
rect 194574 489922 194642 489978
rect 194698 489922 225238 489978
rect 225294 489922 225362 489978
rect 225418 489922 255958 489978
rect 256014 489922 256082 489978
rect 256138 489922 286678 489978
rect 286734 489922 286802 489978
rect 286858 489922 317398 489978
rect 317454 489922 317522 489978
rect 317578 489922 348118 489978
rect 348174 489922 348242 489978
rect 348298 489922 378838 489978
rect 378894 489922 378962 489978
rect 379018 489922 409558 489978
rect 409614 489922 409682 489978
rect 409738 489922 440278 489978
rect 440334 489922 440402 489978
rect 440458 489922 470998 489978
rect 471054 489922 471122 489978
rect 471178 489922 501718 489978
rect 501774 489922 501842 489978
rect 501898 489922 532438 489978
rect 532494 489922 532562 489978
rect 532618 489922 558474 489978
rect 558530 489922 558598 489978
rect 558654 489922 558722 489978
rect 558778 489922 558846 489978
rect 558902 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597980 489978
rect -1916 489891 597980 489922
rect -1916 489835 80457 489891
rect 80513 489835 80561 489891
rect 80617 489835 80665 489891
rect 80721 489835 80769 489891
rect 80825 489835 80873 489891
rect 80929 489835 80977 489891
rect 81033 489835 81081 489891
rect 81137 489835 81185 489891
rect 81241 489835 81289 489891
rect 81345 489835 81393 489891
rect 81449 489835 81497 489891
rect 81553 489835 81601 489891
rect 81657 489835 81705 489891
rect 81761 489835 81809 489891
rect 81865 489835 81913 489891
rect 81969 489835 82017 489891
rect 82073 489835 82121 489891
rect 82177 489835 82225 489891
rect 82281 489835 82329 489891
rect 82385 489835 82433 489891
rect 82489 489835 82537 489891
rect 82593 489835 597980 489891
rect -1916 489826 597980 489835
rect -1916 478350 597980 478446
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 9234 478350
rect 9290 478294 9358 478350
rect 9414 478294 9482 478350
rect 9538 478294 9606 478350
rect 9662 478294 39954 478350
rect 40010 478294 40078 478350
rect 40134 478294 40202 478350
rect 40258 478294 40326 478350
rect 40382 478294 70674 478350
rect 70730 478294 70798 478350
rect 70854 478294 70922 478350
rect 70978 478294 71046 478350
rect 71102 478294 101394 478350
rect 101450 478294 101518 478350
rect 101574 478294 101642 478350
rect 101698 478294 101766 478350
rect 101822 478294 132114 478350
rect 132170 478294 132238 478350
rect 132294 478294 132362 478350
rect 132418 478294 132486 478350
rect 132542 478294 162834 478350
rect 162890 478294 162958 478350
rect 163014 478294 163082 478350
rect 163138 478294 163206 478350
rect 163262 478294 209878 478350
rect 209934 478294 210002 478350
rect 210058 478294 240598 478350
rect 240654 478294 240722 478350
rect 240778 478294 271318 478350
rect 271374 478294 271442 478350
rect 271498 478294 302038 478350
rect 302094 478294 302162 478350
rect 302218 478294 332758 478350
rect 332814 478294 332882 478350
rect 332938 478294 363478 478350
rect 363534 478294 363602 478350
rect 363658 478294 394198 478350
rect 394254 478294 394322 478350
rect 394378 478294 424918 478350
rect 424974 478294 425042 478350
rect 425098 478294 455638 478350
rect 455694 478294 455762 478350
rect 455818 478294 486358 478350
rect 486414 478294 486482 478350
rect 486538 478294 517078 478350
rect 517134 478294 517202 478350
rect 517258 478294 547798 478350
rect 547854 478294 547922 478350
rect 547978 478294 562194 478350
rect 562250 478294 562318 478350
rect 562374 478294 562442 478350
rect 562498 478294 562566 478350
rect 562622 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect -1916 478226 597980 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 9234 478226
rect 9290 478170 9358 478226
rect 9414 478170 9482 478226
rect 9538 478170 9606 478226
rect 9662 478170 39954 478226
rect 40010 478170 40078 478226
rect 40134 478170 40202 478226
rect 40258 478170 40326 478226
rect 40382 478170 70674 478226
rect 70730 478170 70798 478226
rect 70854 478170 70922 478226
rect 70978 478170 71046 478226
rect 71102 478170 101394 478226
rect 101450 478170 101518 478226
rect 101574 478170 101642 478226
rect 101698 478170 101766 478226
rect 101822 478170 132114 478226
rect 132170 478170 132238 478226
rect 132294 478170 132362 478226
rect 132418 478170 132486 478226
rect 132542 478170 162834 478226
rect 162890 478170 162958 478226
rect 163014 478170 163082 478226
rect 163138 478170 163206 478226
rect 163262 478170 209878 478226
rect 209934 478170 210002 478226
rect 210058 478170 240598 478226
rect 240654 478170 240722 478226
rect 240778 478170 271318 478226
rect 271374 478170 271442 478226
rect 271498 478170 302038 478226
rect 302094 478170 302162 478226
rect 302218 478170 332758 478226
rect 332814 478170 332882 478226
rect 332938 478170 363478 478226
rect 363534 478170 363602 478226
rect 363658 478170 394198 478226
rect 394254 478170 394322 478226
rect 394378 478170 424918 478226
rect 424974 478170 425042 478226
rect 425098 478170 455638 478226
rect 455694 478170 455762 478226
rect 455818 478170 486358 478226
rect 486414 478170 486482 478226
rect 486538 478170 517078 478226
rect 517134 478170 517202 478226
rect 517258 478170 547798 478226
rect 547854 478170 547922 478226
rect 547978 478170 562194 478226
rect 562250 478170 562318 478226
rect 562374 478170 562442 478226
rect 562498 478170 562566 478226
rect 562622 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect -1916 478102 597980 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 9234 478102
rect 9290 478046 9358 478102
rect 9414 478046 9482 478102
rect 9538 478046 9606 478102
rect 9662 478046 39954 478102
rect 40010 478046 40078 478102
rect 40134 478046 40202 478102
rect 40258 478046 40326 478102
rect 40382 478046 70674 478102
rect 70730 478046 70798 478102
rect 70854 478046 70922 478102
rect 70978 478046 71046 478102
rect 71102 478046 101394 478102
rect 101450 478046 101518 478102
rect 101574 478046 101642 478102
rect 101698 478046 101766 478102
rect 101822 478046 132114 478102
rect 132170 478046 132238 478102
rect 132294 478046 132362 478102
rect 132418 478046 132486 478102
rect 132542 478046 162834 478102
rect 162890 478046 162958 478102
rect 163014 478046 163082 478102
rect 163138 478046 163206 478102
rect 163262 478046 209878 478102
rect 209934 478046 210002 478102
rect 210058 478046 240598 478102
rect 240654 478046 240722 478102
rect 240778 478046 271318 478102
rect 271374 478046 271442 478102
rect 271498 478046 302038 478102
rect 302094 478046 302162 478102
rect 302218 478046 332758 478102
rect 332814 478046 332882 478102
rect 332938 478046 363478 478102
rect 363534 478046 363602 478102
rect 363658 478046 394198 478102
rect 394254 478046 394322 478102
rect 394378 478046 424918 478102
rect 424974 478046 425042 478102
rect 425098 478046 455638 478102
rect 455694 478046 455762 478102
rect 455818 478046 486358 478102
rect 486414 478046 486482 478102
rect 486538 478046 517078 478102
rect 517134 478046 517202 478102
rect 517258 478046 547798 478102
rect 547854 478046 547922 478102
rect 547978 478046 562194 478102
rect 562250 478046 562318 478102
rect 562374 478046 562442 478102
rect 562498 478046 562566 478102
rect 562622 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect -1916 477978 597980 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 9234 477978
rect 9290 477922 9358 477978
rect 9414 477922 9482 477978
rect 9538 477922 9606 477978
rect 9662 477922 39954 477978
rect 40010 477922 40078 477978
rect 40134 477922 40202 477978
rect 40258 477922 40326 477978
rect 40382 477922 70674 477978
rect 70730 477922 70798 477978
rect 70854 477922 70922 477978
rect 70978 477922 71046 477978
rect 71102 477922 101394 477978
rect 101450 477922 101518 477978
rect 101574 477922 101642 477978
rect 101698 477922 101766 477978
rect 101822 477922 132114 477978
rect 132170 477922 132238 477978
rect 132294 477922 132362 477978
rect 132418 477922 132486 477978
rect 132542 477922 162834 477978
rect 162890 477922 162958 477978
rect 163014 477922 163082 477978
rect 163138 477922 163206 477978
rect 163262 477922 209878 477978
rect 209934 477922 210002 477978
rect 210058 477922 240598 477978
rect 240654 477922 240722 477978
rect 240778 477922 271318 477978
rect 271374 477922 271442 477978
rect 271498 477922 302038 477978
rect 302094 477922 302162 477978
rect 302218 477922 332758 477978
rect 332814 477922 332882 477978
rect 332938 477922 363478 477978
rect 363534 477922 363602 477978
rect 363658 477922 394198 477978
rect 394254 477922 394322 477978
rect 394378 477922 424918 477978
rect 424974 477922 425042 477978
rect 425098 477922 455638 477978
rect 455694 477922 455762 477978
rect 455818 477922 486358 477978
rect 486414 477922 486482 477978
rect 486538 477922 517078 477978
rect 517134 477922 517202 477978
rect 517258 477922 547798 477978
rect 547854 477922 547922 477978
rect 547978 477922 562194 477978
rect 562250 477922 562318 477978
rect 562374 477922 562442 477978
rect 562498 477922 562566 477978
rect 562622 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect -1916 477826 597980 477922
rect -1916 472350 597980 472446
rect -1916 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 36234 472350
rect 36290 472294 36358 472350
rect 36414 472294 36482 472350
rect 36538 472294 36606 472350
rect 36662 472294 66954 472350
rect 67010 472294 67078 472350
rect 67134 472294 67202 472350
rect 67258 472294 67326 472350
rect 67382 472294 97674 472350
rect 97730 472294 97798 472350
rect 97854 472294 97922 472350
rect 97978 472294 98046 472350
rect 98102 472294 128394 472350
rect 128450 472294 128518 472350
rect 128574 472294 128642 472350
rect 128698 472294 128766 472350
rect 128822 472294 159114 472350
rect 159170 472294 159238 472350
rect 159294 472294 159362 472350
rect 159418 472294 159486 472350
rect 159542 472294 189834 472350
rect 189890 472294 189958 472350
rect 190014 472294 190082 472350
rect 190138 472294 190206 472350
rect 190262 472294 194518 472350
rect 194574 472294 194642 472350
rect 194698 472294 225238 472350
rect 225294 472294 225362 472350
rect 225418 472294 255958 472350
rect 256014 472294 256082 472350
rect 256138 472294 286678 472350
rect 286734 472294 286802 472350
rect 286858 472294 317398 472350
rect 317454 472294 317522 472350
rect 317578 472294 348118 472350
rect 348174 472294 348242 472350
rect 348298 472294 378838 472350
rect 378894 472294 378962 472350
rect 379018 472294 409558 472350
rect 409614 472294 409682 472350
rect 409738 472294 440278 472350
rect 440334 472294 440402 472350
rect 440458 472294 470998 472350
rect 471054 472294 471122 472350
rect 471178 472294 501718 472350
rect 501774 472294 501842 472350
rect 501898 472294 532438 472350
rect 532494 472294 532562 472350
rect 532618 472294 558474 472350
rect 558530 472294 558598 472350
rect 558654 472294 558722 472350
rect 558778 472294 558846 472350
rect 558902 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597980 472350
rect -1916 472226 597980 472294
rect -1916 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 36234 472226
rect 36290 472170 36358 472226
rect 36414 472170 36482 472226
rect 36538 472170 36606 472226
rect 36662 472170 66954 472226
rect 67010 472170 67078 472226
rect 67134 472170 67202 472226
rect 67258 472170 67326 472226
rect 67382 472170 97674 472226
rect 97730 472170 97798 472226
rect 97854 472170 97922 472226
rect 97978 472170 98046 472226
rect 98102 472170 128394 472226
rect 128450 472170 128518 472226
rect 128574 472170 128642 472226
rect 128698 472170 128766 472226
rect 128822 472170 159114 472226
rect 159170 472170 159238 472226
rect 159294 472170 159362 472226
rect 159418 472170 159486 472226
rect 159542 472170 189834 472226
rect 189890 472170 189958 472226
rect 190014 472170 190082 472226
rect 190138 472170 190206 472226
rect 190262 472170 194518 472226
rect 194574 472170 194642 472226
rect 194698 472170 225238 472226
rect 225294 472170 225362 472226
rect 225418 472170 255958 472226
rect 256014 472170 256082 472226
rect 256138 472170 286678 472226
rect 286734 472170 286802 472226
rect 286858 472170 317398 472226
rect 317454 472170 317522 472226
rect 317578 472170 348118 472226
rect 348174 472170 348242 472226
rect 348298 472170 378838 472226
rect 378894 472170 378962 472226
rect 379018 472170 409558 472226
rect 409614 472170 409682 472226
rect 409738 472170 440278 472226
rect 440334 472170 440402 472226
rect 440458 472170 470998 472226
rect 471054 472170 471122 472226
rect 471178 472170 501718 472226
rect 501774 472170 501842 472226
rect 501898 472170 532438 472226
rect 532494 472170 532562 472226
rect 532618 472170 558474 472226
rect 558530 472170 558598 472226
rect 558654 472170 558722 472226
rect 558778 472170 558846 472226
rect 558902 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597980 472226
rect -1916 472102 597980 472170
rect -1916 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 36234 472102
rect 36290 472046 36358 472102
rect 36414 472046 36482 472102
rect 36538 472046 36606 472102
rect 36662 472046 66954 472102
rect 67010 472046 67078 472102
rect 67134 472046 67202 472102
rect 67258 472046 67326 472102
rect 67382 472046 97674 472102
rect 97730 472046 97798 472102
rect 97854 472046 97922 472102
rect 97978 472046 98046 472102
rect 98102 472046 128394 472102
rect 128450 472046 128518 472102
rect 128574 472046 128642 472102
rect 128698 472046 128766 472102
rect 128822 472046 159114 472102
rect 159170 472046 159238 472102
rect 159294 472046 159362 472102
rect 159418 472046 159486 472102
rect 159542 472046 189834 472102
rect 189890 472046 189958 472102
rect 190014 472046 190082 472102
rect 190138 472046 190206 472102
rect 190262 472046 194518 472102
rect 194574 472046 194642 472102
rect 194698 472046 225238 472102
rect 225294 472046 225362 472102
rect 225418 472046 255958 472102
rect 256014 472046 256082 472102
rect 256138 472046 286678 472102
rect 286734 472046 286802 472102
rect 286858 472046 317398 472102
rect 317454 472046 317522 472102
rect 317578 472046 348118 472102
rect 348174 472046 348242 472102
rect 348298 472046 378838 472102
rect 378894 472046 378962 472102
rect 379018 472046 409558 472102
rect 409614 472046 409682 472102
rect 409738 472046 440278 472102
rect 440334 472046 440402 472102
rect 440458 472046 470998 472102
rect 471054 472046 471122 472102
rect 471178 472046 501718 472102
rect 501774 472046 501842 472102
rect 501898 472046 532438 472102
rect 532494 472046 532562 472102
rect 532618 472046 558474 472102
rect 558530 472046 558598 472102
rect 558654 472046 558722 472102
rect 558778 472046 558846 472102
rect 558902 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597980 472102
rect -1916 471978 597980 472046
rect -1916 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 36234 471978
rect 36290 471922 36358 471978
rect 36414 471922 36482 471978
rect 36538 471922 36606 471978
rect 36662 471922 66954 471978
rect 67010 471922 67078 471978
rect 67134 471922 67202 471978
rect 67258 471922 67326 471978
rect 67382 471922 97674 471978
rect 97730 471922 97798 471978
rect 97854 471922 97922 471978
rect 97978 471922 98046 471978
rect 98102 471922 128394 471978
rect 128450 471922 128518 471978
rect 128574 471922 128642 471978
rect 128698 471922 128766 471978
rect 128822 471922 159114 471978
rect 159170 471922 159238 471978
rect 159294 471922 159362 471978
rect 159418 471922 159486 471978
rect 159542 471922 189834 471978
rect 189890 471922 189958 471978
rect 190014 471922 190082 471978
rect 190138 471922 190206 471978
rect 190262 471922 194518 471978
rect 194574 471922 194642 471978
rect 194698 471922 225238 471978
rect 225294 471922 225362 471978
rect 225418 471922 255958 471978
rect 256014 471922 256082 471978
rect 256138 471922 286678 471978
rect 286734 471922 286802 471978
rect 286858 471922 317398 471978
rect 317454 471922 317522 471978
rect 317578 471922 348118 471978
rect 348174 471922 348242 471978
rect 348298 471922 378838 471978
rect 378894 471922 378962 471978
rect 379018 471922 409558 471978
rect 409614 471922 409682 471978
rect 409738 471922 440278 471978
rect 440334 471922 440402 471978
rect 440458 471922 470998 471978
rect 471054 471922 471122 471978
rect 471178 471922 501718 471978
rect 501774 471922 501842 471978
rect 501898 471922 532438 471978
rect 532494 471922 532562 471978
rect 532618 471922 558474 471978
rect 558530 471922 558598 471978
rect 558654 471922 558722 471978
rect 558778 471922 558846 471978
rect 558902 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597980 471978
rect -1916 471826 597980 471922
rect -1916 460350 597980 460446
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 9234 460350
rect 9290 460294 9358 460350
rect 9414 460294 9482 460350
rect 9538 460294 9606 460350
rect 9662 460294 39954 460350
rect 40010 460294 40078 460350
rect 40134 460294 40202 460350
rect 40258 460294 40326 460350
rect 40382 460294 70674 460350
rect 70730 460294 70798 460350
rect 70854 460294 70922 460350
rect 70978 460294 71046 460350
rect 71102 460294 101394 460350
rect 101450 460294 101518 460350
rect 101574 460294 101642 460350
rect 101698 460294 101766 460350
rect 101822 460294 132114 460350
rect 132170 460294 132238 460350
rect 132294 460294 132362 460350
rect 132418 460294 132486 460350
rect 132542 460294 162834 460350
rect 162890 460294 162958 460350
rect 163014 460294 163082 460350
rect 163138 460294 163206 460350
rect 163262 460294 209878 460350
rect 209934 460294 210002 460350
rect 210058 460294 240598 460350
rect 240654 460294 240722 460350
rect 240778 460294 271318 460350
rect 271374 460294 271442 460350
rect 271498 460294 302038 460350
rect 302094 460294 302162 460350
rect 302218 460294 332758 460350
rect 332814 460294 332882 460350
rect 332938 460294 363478 460350
rect 363534 460294 363602 460350
rect 363658 460294 394198 460350
rect 394254 460294 394322 460350
rect 394378 460294 424918 460350
rect 424974 460294 425042 460350
rect 425098 460294 455638 460350
rect 455694 460294 455762 460350
rect 455818 460294 486358 460350
rect 486414 460294 486482 460350
rect 486538 460294 517078 460350
rect 517134 460294 517202 460350
rect 517258 460294 547798 460350
rect 547854 460294 547922 460350
rect 547978 460294 562194 460350
rect 562250 460294 562318 460350
rect 562374 460294 562442 460350
rect 562498 460294 562566 460350
rect 562622 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect -1916 460226 597980 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 9234 460226
rect 9290 460170 9358 460226
rect 9414 460170 9482 460226
rect 9538 460170 9606 460226
rect 9662 460170 39954 460226
rect 40010 460170 40078 460226
rect 40134 460170 40202 460226
rect 40258 460170 40326 460226
rect 40382 460170 70674 460226
rect 70730 460170 70798 460226
rect 70854 460170 70922 460226
rect 70978 460170 71046 460226
rect 71102 460170 101394 460226
rect 101450 460170 101518 460226
rect 101574 460170 101642 460226
rect 101698 460170 101766 460226
rect 101822 460170 132114 460226
rect 132170 460170 132238 460226
rect 132294 460170 132362 460226
rect 132418 460170 132486 460226
rect 132542 460170 162834 460226
rect 162890 460170 162958 460226
rect 163014 460170 163082 460226
rect 163138 460170 163206 460226
rect 163262 460170 209878 460226
rect 209934 460170 210002 460226
rect 210058 460170 240598 460226
rect 240654 460170 240722 460226
rect 240778 460170 271318 460226
rect 271374 460170 271442 460226
rect 271498 460170 302038 460226
rect 302094 460170 302162 460226
rect 302218 460170 332758 460226
rect 332814 460170 332882 460226
rect 332938 460170 363478 460226
rect 363534 460170 363602 460226
rect 363658 460170 394198 460226
rect 394254 460170 394322 460226
rect 394378 460170 424918 460226
rect 424974 460170 425042 460226
rect 425098 460170 455638 460226
rect 455694 460170 455762 460226
rect 455818 460170 486358 460226
rect 486414 460170 486482 460226
rect 486538 460170 517078 460226
rect 517134 460170 517202 460226
rect 517258 460170 547798 460226
rect 547854 460170 547922 460226
rect 547978 460170 562194 460226
rect 562250 460170 562318 460226
rect 562374 460170 562442 460226
rect 562498 460170 562566 460226
rect 562622 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect -1916 460102 597980 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 9234 460102
rect 9290 460046 9358 460102
rect 9414 460046 9482 460102
rect 9538 460046 9606 460102
rect 9662 460046 39954 460102
rect 40010 460046 40078 460102
rect 40134 460046 40202 460102
rect 40258 460046 40326 460102
rect 40382 460046 70674 460102
rect 70730 460046 70798 460102
rect 70854 460046 70922 460102
rect 70978 460046 71046 460102
rect 71102 460046 101394 460102
rect 101450 460046 101518 460102
rect 101574 460046 101642 460102
rect 101698 460046 101766 460102
rect 101822 460046 132114 460102
rect 132170 460046 132238 460102
rect 132294 460046 132362 460102
rect 132418 460046 132486 460102
rect 132542 460046 162834 460102
rect 162890 460046 162958 460102
rect 163014 460046 163082 460102
rect 163138 460046 163206 460102
rect 163262 460046 209878 460102
rect 209934 460046 210002 460102
rect 210058 460046 240598 460102
rect 240654 460046 240722 460102
rect 240778 460046 271318 460102
rect 271374 460046 271442 460102
rect 271498 460046 302038 460102
rect 302094 460046 302162 460102
rect 302218 460046 332758 460102
rect 332814 460046 332882 460102
rect 332938 460046 363478 460102
rect 363534 460046 363602 460102
rect 363658 460046 394198 460102
rect 394254 460046 394322 460102
rect 394378 460046 424918 460102
rect 424974 460046 425042 460102
rect 425098 460046 455638 460102
rect 455694 460046 455762 460102
rect 455818 460046 486358 460102
rect 486414 460046 486482 460102
rect 486538 460046 517078 460102
rect 517134 460046 517202 460102
rect 517258 460046 547798 460102
rect 547854 460046 547922 460102
rect 547978 460046 562194 460102
rect 562250 460046 562318 460102
rect 562374 460046 562442 460102
rect 562498 460046 562566 460102
rect 562622 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect -1916 459978 597980 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 9234 459978
rect 9290 459922 9358 459978
rect 9414 459922 9482 459978
rect 9538 459922 9606 459978
rect 9662 459922 39954 459978
rect 40010 459922 40078 459978
rect 40134 459922 40202 459978
rect 40258 459922 40326 459978
rect 40382 459922 70674 459978
rect 70730 459922 70798 459978
rect 70854 459922 70922 459978
rect 70978 459922 71046 459978
rect 71102 459922 101394 459978
rect 101450 459922 101518 459978
rect 101574 459922 101642 459978
rect 101698 459922 101766 459978
rect 101822 459922 132114 459978
rect 132170 459922 132238 459978
rect 132294 459922 132362 459978
rect 132418 459922 132486 459978
rect 132542 459922 162834 459978
rect 162890 459922 162958 459978
rect 163014 459922 163082 459978
rect 163138 459922 163206 459978
rect 163262 459922 209878 459978
rect 209934 459922 210002 459978
rect 210058 459922 240598 459978
rect 240654 459922 240722 459978
rect 240778 459922 271318 459978
rect 271374 459922 271442 459978
rect 271498 459922 302038 459978
rect 302094 459922 302162 459978
rect 302218 459922 332758 459978
rect 332814 459922 332882 459978
rect 332938 459922 363478 459978
rect 363534 459922 363602 459978
rect 363658 459922 394198 459978
rect 394254 459922 394322 459978
rect 394378 459922 424918 459978
rect 424974 459922 425042 459978
rect 425098 459922 455638 459978
rect 455694 459922 455762 459978
rect 455818 459922 486358 459978
rect 486414 459922 486482 459978
rect 486538 459922 517078 459978
rect 517134 459922 517202 459978
rect 517258 459922 547798 459978
rect 547854 459922 547922 459978
rect 547978 459922 562194 459978
rect 562250 459922 562318 459978
rect 562374 459922 562442 459978
rect 562498 459922 562566 459978
rect 562622 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect -1916 459826 597980 459922
rect -1916 454350 597980 454446
rect -1916 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 36234 454350
rect 36290 454294 36358 454350
rect 36414 454294 36482 454350
rect 36538 454294 36606 454350
rect 36662 454294 66954 454350
rect 67010 454294 67078 454350
rect 67134 454294 67202 454350
rect 67258 454294 67326 454350
rect 67382 454294 97674 454350
rect 97730 454294 97798 454350
rect 97854 454294 97922 454350
rect 97978 454294 98046 454350
rect 98102 454294 128394 454350
rect 128450 454294 128518 454350
rect 128574 454294 128642 454350
rect 128698 454294 128766 454350
rect 128822 454294 159114 454350
rect 159170 454294 159238 454350
rect 159294 454294 159362 454350
rect 159418 454294 159486 454350
rect 159542 454294 189834 454350
rect 189890 454294 189958 454350
rect 190014 454294 190082 454350
rect 190138 454294 190206 454350
rect 190262 454294 194518 454350
rect 194574 454294 194642 454350
rect 194698 454294 225238 454350
rect 225294 454294 225362 454350
rect 225418 454294 255958 454350
rect 256014 454294 256082 454350
rect 256138 454294 286678 454350
rect 286734 454294 286802 454350
rect 286858 454294 317398 454350
rect 317454 454294 317522 454350
rect 317578 454294 348118 454350
rect 348174 454294 348242 454350
rect 348298 454294 378838 454350
rect 378894 454294 378962 454350
rect 379018 454294 409558 454350
rect 409614 454294 409682 454350
rect 409738 454294 440278 454350
rect 440334 454294 440402 454350
rect 440458 454294 470998 454350
rect 471054 454294 471122 454350
rect 471178 454294 501718 454350
rect 501774 454294 501842 454350
rect 501898 454294 532438 454350
rect 532494 454294 532562 454350
rect 532618 454294 558474 454350
rect 558530 454294 558598 454350
rect 558654 454294 558722 454350
rect 558778 454294 558846 454350
rect 558902 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597980 454350
rect -1916 454226 597980 454294
rect -1916 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 36234 454226
rect 36290 454170 36358 454226
rect 36414 454170 36482 454226
rect 36538 454170 36606 454226
rect 36662 454170 66954 454226
rect 67010 454170 67078 454226
rect 67134 454170 67202 454226
rect 67258 454170 67326 454226
rect 67382 454170 97674 454226
rect 97730 454170 97798 454226
rect 97854 454170 97922 454226
rect 97978 454170 98046 454226
rect 98102 454170 128394 454226
rect 128450 454170 128518 454226
rect 128574 454170 128642 454226
rect 128698 454170 128766 454226
rect 128822 454170 159114 454226
rect 159170 454170 159238 454226
rect 159294 454170 159362 454226
rect 159418 454170 159486 454226
rect 159542 454170 189834 454226
rect 189890 454170 189958 454226
rect 190014 454170 190082 454226
rect 190138 454170 190206 454226
rect 190262 454170 194518 454226
rect 194574 454170 194642 454226
rect 194698 454170 225238 454226
rect 225294 454170 225362 454226
rect 225418 454170 255958 454226
rect 256014 454170 256082 454226
rect 256138 454170 286678 454226
rect 286734 454170 286802 454226
rect 286858 454170 317398 454226
rect 317454 454170 317522 454226
rect 317578 454170 348118 454226
rect 348174 454170 348242 454226
rect 348298 454170 378838 454226
rect 378894 454170 378962 454226
rect 379018 454170 409558 454226
rect 409614 454170 409682 454226
rect 409738 454170 440278 454226
rect 440334 454170 440402 454226
rect 440458 454170 470998 454226
rect 471054 454170 471122 454226
rect 471178 454170 501718 454226
rect 501774 454170 501842 454226
rect 501898 454170 532438 454226
rect 532494 454170 532562 454226
rect 532618 454170 558474 454226
rect 558530 454170 558598 454226
rect 558654 454170 558722 454226
rect 558778 454170 558846 454226
rect 558902 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597980 454226
rect -1916 454102 597980 454170
rect -1916 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 36234 454102
rect 36290 454046 36358 454102
rect 36414 454046 36482 454102
rect 36538 454046 36606 454102
rect 36662 454046 66954 454102
rect 67010 454046 67078 454102
rect 67134 454046 67202 454102
rect 67258 454046 67326 454102
rect 67382 454046 97674 454102
rect 97730 454046 97798 454102
rect 97854 454046 97922 454102
rect 97978 454046 98046 454102
rect 98102 454046 128394 454102
rect 128450 454046 128518 454102
rect 128574 454046 128642 454102
rect 128698 454046 128766 454102
rect 128822 454046 159114 454102
rect 159170 454046 159238 454102
rect 159294 454046 159362 454102
rect 159418 454046 159486 454102
rect 159542 454046 189834 454102
rect 189890 454046 189958 454102
rect 190014 454046 190082 454102
rect 190138 454046 190206 454102
rect 190262 454046 194518 454102
rect 194574 454046 194642 454102
rect 194698 454046 225238 454102
rect 225294 454046 225362 454102
rect 225418 454046 255958 454102
rect 256014 454046 256082 454102
rect 256138 454046 286678 454102
rect 286734 454046 286802 454102
rect 286858 454046 317398 454102
rect 317454 454046 317522 454102
rect 317578 454046 348118 454102
rect 348174 454046 348242 454102
rect 348298 454046 378838 454102
rect 378894 454046 378962 454102
rect 379018 454046 409558 454102
rect 409614 454046 409682 454102
rect 409738 454046 440278 454102
rect 440334 454046 440402 454102
rect 440458 454046 470998 454102
rect 471054 454046 471122 454102
rect 471178 454046 501718 454102
rect 501774 454046 501842 454102
rect 501898 454046 532438 454102
rect 532494 454046 532562 454102
rect 532618 454046 558474 454102
rect 558530 454046 558598 454102
rect 558654 454046 558722 454102
rect 558778 454046 558846 454102
rect 558902 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597980 454102
rect -1916 453978 597980 454046
rect -1916 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 36234 453978
rect 36290 453922 36358 453978
rect 36414 453922 36482 453978
rect 36538 453922 36606 453978
rect 36662 453922 66954 453978
rect 67010 453922 67078 453978
rect 67134 453922 67202 453978
rect 67258 453922 67326 453978
rect 67382 453922 97674 453978
rect 97730 453922 97798 453978
rect 97854 453922 97922 453978
rect 97978 453922 98046 453978
rect 98102 453922 128394 453978
rect 128450 453922 128518 453978
rect 128574 453922 128642 453978
rect 128698 453922 128766 453978
rect 128822 453922 159114 453978
rect 159170 453922 159238 453978
rect 159294 453922 159362 453978
rect 159418 453922 159486 453978
rect 159542 453922 189834 453978
rect 189890 453922 189958 453978
rect 190014 453922 190082 453978
rect 190138 453922 190206 453978
rect 190262 453922 194518 453978
rect 194574 453922 194642 453978
rect 194698 453922 225238 453978
rect 225294 453922 225362 453978
rect 225418 453922 255958 453978
rect 256014 453922 256082 453978
rect 256138 453922 286678 453978
rect 286734 453922 286802 453978
rect 286858 453922 317398 453978
rect 317454 453922 317522 453978
rect 317578 453922 348118 453978
rect 348174 453922 348242 453978
rect 348298 453922 378838 453978
rect 378894 453922 378962 453978
rect 379018 453922 409558 453978
rect 409614 453922 409682 453978
rect 409738 453922 440278 453978
rect 440334 453922 440402 453978
rect 440458 453922 470998 453978
rect 471054 453922 471122 453978
rect 471178 453922 501718 453978
rect 501774 453922 501842 453978
rect 501898 453922 532438 453978
rect 532494 453922 532562 453978
rect 532618 453922 558474 453978
rect 558530 453922 558598 453978
rect 558654 453922 558722 453978
rect 558778 453922 558846 453978
rect 558902 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597980 453978
rect -1916 453826 597980 453922
rect -1916 442350 597980 442446
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 9234 442350
rect 9290 442294 9358 442350
rect 9414 442294 9482 442350
rect 9538 442294 9606 442350
rect 9662 442294 39954 442350
rect 40010 442294 40078 442350
rect 40134 442294 40202 442350
rect 40258 442294 40326 442350
rect 40382 442294 70674 442350
rect 70730 442294 70798 442350
rect 70854 442294 70922 442350
rect 70978 442294 71046 442350
rect 71102 442294 101394 442350
rect 101450 442294 101518 442350
rect 101574 442294 101642 442350
rect 101698 442294 101766 442350
rect 101822 442294 132114 442350
rect 132170 442294 132238 442350
rect 132294 442294 132362 442350
rect 132418 442294 132486 442350
rect 132542 442294 162834 442350
rect 162890 442294 162958 442350
rect 163014 442294 163082 442350
rect 163138 442294 163206 442350
rect 163262 442294 209878 442350
rect 209934 442294 210002 442350
rect 210058 442294 240598 442350
rect 240654 442294 240722 442350
rect 240778 442294 271318 442350
rect 271374 442294 271442 442350
rect 271498 442294 302038 442350
rect 302094 442294 302162 442350
rect 302218 442294 332758 442350
rect 332814 442294 332882 442350
rect 332938 442294 363478 442350
rect 363534 442294 363602 442350
rect 363658 442294 394198 442350
rect 394254 442294 394322 442350
rect 394378 442294 424918 442350
rect 424974 442294 425042 442350
rect 425098 442294 455638 442350
rect 455694 442294 455762 442350
rect 455818 442294 486358 442350
rect 486414 442294 486482 442350
rect 486538 442294 517078 442350
rect 517134 442294 517202 442350
rect 517258 442294 547798 442350
rect 547854 442294 547922 442350
rect 547978 442294 562194 442350
rect 562250 442294 562318 442350
rect 562374 442294 562442 442350
rect 562498 442294 562566 442350
rect 562622 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect -1916 442226 597980 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 9234 442226
rect 9290 442170 9358 442226
rect 9414 442170 9482 442226
rect 9538 442170 9606 442226
rect 9662 442170 39954 442226
rect 40010 442170 40078 442226
rect 40134 442170 40202 442226
rect 40258 442170 40326 442226
rect 40382 442170 70674 442226
rect 70730 442170 70798 442226
rect 70854 442170 70922 442226
rect 70978 442170 71046 442226
rect 71102 442170 101394 442226
rect 101450 442170 101518 442226
rect 101574 442170 101642 442226
rect 101698 442170 101766 442226
rect 101822 442170 132114 442226
rect 132170 442170 132238 442226
rect 132294 442170 132362 442226
rect 132418 442170 132486 442226
rect 132542 442170 162834 442226
rect 162890 442170 162958 442226
rect 163014 442170 163082 442226
rect 163138 442170 163206 442226
rect 163262 442170 209878 442226
rect 209934 442170 210002 442226
rect 210058 442170 240598 442226
rect 240654 442170 240722 442226
rect 240778 442170 271318 442226
rect 271374 442170 271442 442226
rect 271498 442170 302038 442226
rect 302094 442170 302162 442226
rect 302218 442170 332758 442226
rect 332814 442170 332882 442226
rect 332938 442170 363478 442226
rect 363534 442170 363602 442226
rect 363658 442170 394198 442226
rect 394254 442170 394322 442226
rect 394378 442170 424918 442226
rect 424974 442170 425042 442226
rect 425098 442170 455638 442226
rect 455694 442170 455762 442226
rect 455818 442170 486358 442226
rect 486414 442170 486482 442226
rect 486538 442170 517078 442226
rect 517134 442170 517202 442226
rect 517258 442170 547798 442226
rect 547854 442170 547922 442226
rect 547978 442170 562194 442226
rect 562250 442170 562318 442226
rect 562374 442170 562442 442226
rect 562498 442170 562566 442226
rect 562622 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect -1916 442102 597980 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 9234 442102
rect 9290 442046 9358 442102
rect 9414 442046 9482 442102
rect 9538 442046 9606 442102
rect 9662 442046 39954 442102
rect 40010 442046 40078 442102
rect 40134 442046 40202 442102
rect 40258 442046 40326 442102
rect 40382 442046 70674 442102
rect 70730 442046 70798 442102
rect 70854 442046 70922 442102
rect 70978 442046 71046 442102
rect 71102 442046 101394 442102
rect 101450 442046 101518 442102
rect 101574 442046 101642 442102
rect 101698 442046 101766 442102
rect 101822 442046 132114 442102
rect 132170 442046 132238 442102
rect 132294 442046 132362 442102
rect 132418 442046 132486 442102
rect 132542 442046 162834 442102
rect 162890 442046 162958 442102
rect 163014 442046 163082 442102
rect 163138 442046 163206 442102
rect 163262 442046 209878 442102
rect 209934 442046 210002 442102
rect 210058 442046 240598 442102
rect 240654 442046 240722 442102
rect 240778 442046 271318 442102
rect 271374 442046 271442 442102
rect 271498 442046 302038 442102
rect 302094 442046 302162 442102
rect 302218 442046 332758 442102
rect 332814 442046 332882 442102
rect 332938 442046 363478 442102
rect 363534 442046 363602 442102
rect 363658 442046 394198 442102
rect 394254 442046 394322 442102
rect 394378 442046 424918 442102
rect 424974 442046 425042 442102
rect 425098 442046 455638 442102
rect 455694 442046 455762 442102
rect 455818 442046 486358 442102
rect 486414 442046 486482 442102
rect 486538 442046 517078 442102
rect 517134 442046 517202 442102
rect 517258 442046 547798 442102
rect 547854 442046 547922 442102
rect 547978 442046 562194 442102
rect 562250 442046 562318 442102
rect 562374 442046 562442 442102
rect 562498 442046 562566 442102
rect 562622 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect -1916 441978 597980 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 9234 441978
rect 9290 441922 9358 441978
rect 9414 441922 9482 441978
rect 9538 441922 9606 441978
rect 9662 441922 39954 441978
rect 40010 441922 40078 441978
rect 40134 441922 40202 441978
rect 40258 441922 40326 441978
rect 40382 441922 70674 441978
rect 70730 441922 70798 441978
rect 70854 441922 70922 441978
rect 70978 441922 71046 441978
rect 71102 441922 101394 441978
rect 101450 441922 101518 441978
rect 101574 441922 101642 441978
rect 101698 441922 101766 441978
rect 101822 441922 132114 441978
rect 132170 441922 132238 441978
rect 132294 441922 132362 441978
rect 132418 441922 132486 441978
rect 132542 441922 162834 441978
rect 162890 441922 162958 441978
rect 163014 441922 163082 441978
rect 163138 441922 163206 441978
rect 163262 441922 209878 441978
rect 209934 441922 210002 441978
rect 210058 441922 240598 441978
rect 240654 441922 240722 441978
rect 240778 441922 271318 441978
rect 271374 441922 271442 441978
rect 271498 441922 302038 441978
rect 302094 441922 302162 441978
rect 302218 441922 332758 441978
rect 332814 441922 332882 441978
rect 332938 441922 363478 441978
rect 363534 441922 363602 441978
rect 363658 441922 394198 441978
rect 394254 441922 394322 441978
rect 394378 441922 424918 441978
rect 424974 441922 425042 441978
rect 425098 441922 455638 441978
rect 455694 441922 455762 441978
rect 455818 441922 486358 441978
rect 486414 441922 486482 441978
rect 486538 441922 517078 441978
rect 517134 441922 517202 441978
rect 517258 441922 547798 441978
rect 547854 441922 547922 441978
rect 547978 441922 562194 441978
rect 562250 441922 562318 441978
rect 562374 441922 562442 441978
rect 562498 441922 562566 441978
rect 562622 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect -1916 441826 597980 441922
rect -1916 436350 597980 436446
rect -1916 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 36234 436350
rect 36290 436294 36358 436350
rect 36414 436294 36482 436350
rect 36538 436294 36606 436350
rect 36662 436294 66954 436350
rect 67010 436294 67078 436350
rect 67134 436294 67202 436350
rect 67258 436294 67326 436350
rect 67382 436294 97674 436350
rect 97730 436294 97798 436350
rect 97854 436294 97922 436350
rect 97978 436294 98046 436350
rect 98102 436294 128394 436350
rect 128450 436294 128518 436350
rect 128574 436294 128642 436350
rect 128698 436294 128766 436350
rect 128822 436294 159114 436350
rect 159170 436294 159238 436350
rect 159294 436294 159362 436350
rect 159418 436294 159486 436350
rect 159542 436294 189834 436350
rect 189890 436294 189958 436350
rect 190014 436294 190082 436350
rect 190138 436294 190206 436350
rect 190262 436294 194518 436350
rect 194574 436294 194642 436350
rect 194698 436294 225238 436350
rect 225294 436294 225362 436350
rect 225418 436294 255958 436350
rect 256014 436294 256082 436350
rect 256138 436294 286678 436350
rect 286734 436294 286802 436350
rect 286858 436294 317398 436350
rect 317454 436294 317522 436350
rect 317578 436294 348118 436350
rect 348174 436294 348242 436350
rect 348298 436294 378838 436350
rect 378894 436294 378962 436350
rect 379018 436294 409558 436350
rect 409614 436294 409682 436350
rect 409738 436294 440278 436350
rect 440334 436294 440402 436350
rect 440458 436294 470998 436350
rect 471054 436294 471122 436350
rect 471178 436294 501718 436350
rect 501774 436294 501842 436350
rect 501898 436294 532438 436350
rect 532494 436294 532562 436350
rect 532618 436294 558474 436350
rect 558530 436294 558598 436350
rect 558654 436294 558722 436350
rect 558778 436294 558846 436350
rect 558902 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597980 436350
rect -1916 436226 597980 436294
rect -1916 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 36234 436226
rect 36290 436170 36358 436226
rect 36414 436170 36482 436226
rect 36538 436170 36606 436226
rect 36662 436170 66954 436226
rect 67010 436170 67078 436226
rect 67134 436170 67202 436226
rect 67258 436170 67326 436226
rect 67382 436170 97674 436226
rect 97730 436170 97798 436226
rect 97854 436170 97922 436226
rect 97978 436170 98046 436226
rect 98102 436170 128394 436226
rect 128450 436170 128518 436226
rect 128574 436170 128642 436226
rect 128698 436170 128766 436226
rect 128822 436170 159114 436226
rect 159170 436170 159238 436226
rect 159294 436170 159362 436226
rect 159418 436170 159486 436226
rect 159542 436170 189834 436226
rect 189890 436170 189958 436226
rect 190014 436170 190082 436226
rect 190138 436170 190206 436226
rect 190262 436170 194518 436226
rect 194574 436170 194642 436226
rect 194698 436170 225238 436226
rect 225294 436170 225362 436226
rect 225418 436170 255958 436226
rect 256014 436170 256082 436226
rect 256138 436170 286678 436226
rect 286734 436170 286802 436226
rect 286858 436170 317398 436226
rect 317454 436170 317522 436226
rect 317578 436170 348118 436226
rect 348174 436170 348242 436226
rect 348298 436170 378838 436226
rect 378894 436170 378962 436226
rect 379018 436170 409558 436226
rect 409614 436170 409682 436226
rect 409738 436170 440278 436226
rect 440334 436170 440402 436226
rect 440458 436170 470998 436226
rect 471054 436170 471122 436226
rect 471178 436170 501718 436226
rect 501774 436170 501842 436226
rect 501898 436170 532438 436226
rect 532494 436170 532562 436226
rect 532618 436170 558474 436226
rect 558530 436170 558598 436226
rect 558654 436170 558722 436226
rect 558778 436170 558846 436226
rect 558902 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597980 436226
rect -1916 436102 597980 436170
rect -1916 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 36234 436102
rect 36290 436046 36358 436102
rect 36414 436046 36482 436102
rect 36538 436046 36606 436102
rect 36662 436046 66954 436102
rect 67010 436046 67078 436102
rect 67134 436046 67202 436102
rect 67258 436046 67326 436102
rect 67382 436046 97674 436102
rect 97730 436046 97798 436102
rect 97854 436046 97922 436102
rect 97978 436046 98046 436102
rect 98102 436046 128394 436102
rect 128450 436046 128518 436102
rect 128574 436046 128642 436102
rect 128698 436046 128766 436102
rect 128822 436046 159114 436102
rect 159170 436046 159238 436102
rect 159294 436046 159362 436102
rect 159418 436046 159486 436102
rect 159542 436046 189834 436102
rect 189890 436046 189958 436102
rect 190014 436046 190082 436102
rect 190138 436046 190206 436102
rect 190262 436046 194518 436102
rect 194574 436046 194642 436102
rect 194698 436046 225238 436102
rect 225294 436046 225362 436102
rect 225418 436046 255958 436102
rect 256014 436046 256082 436102
rect 256138 436046 286678 436102
rect 286734 436046 286802 436102
rect 286858 436046 317398 436102
rect 317454 436046 317522 436102
rect 317578 436046 348118 436102
rect 348174 436046 348242 436102
rect 348298 436046 378838 436102
rect 378894 436046 378962 436102
rect 379018 436046 409558 436102
rect 409614 436046 409682 436102
rect 409738 436046 440278 436102
rect 440334 436046 440402 436102
rect 440458 436046 470998 436102
rect 471054 436046 471122 436102
rect 471178 436046 501718 436102
rect 501774 436046 501842 436102
rect 501898 436046 532438 436102
rect 532494 436046 532562 436102
rect 532618 436046 558474 436102
rect 558530 436046 558598 436102
rect 558654 436046 558722 436102
rect 558778 436046 558846 436102
rect 558902 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597980 436102
rect -1916 435978 597980 436046
rect -1916 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 36234 435978
rect 36290 435922 36358 435978
rect 36414 435922 36482 435978
rect 36538 435922 36606 435978
rect 36662 435922 66954 435978
rect 67010 435922 67078 435978
rect 67134 435922 67202 435978
rect 67258 435922 67326 435978
rect 67382 435922 97674 435978
rect 97730 435922 97798 435978
rect 97854 435922 97922 435978
rect 97978 435922 98046 435978
rect 98102 435922 128394 435978
rect 128450 435922 128518 435978
rect 128574 435922 128642 435978
rect 128698 435922 128766 435978
rect 128822 435922 159114 435978
rect 159170 435922 159238 435978
rect 159294 435922 159362 435978
rect 159418 435922 159486 435978
rect 159542 435922 189834 435978
rect 189890 435922 189958 435978
rect 190014 435922 190082 435978
rect 190138 435922 190206 435978
rect 190262 435922 194518 435978
rect 194574 435922 194642 435978
rect 194698 435922 225238 435978
rect 225294 435922 225362 435978
rect 225418 435922 255958 435978
rect 256014 435922 256082 435978
rect 256138 435922 286678 435978
rect 286734 435922 286802 435978
rect 286858 435922 317398 435978
rect 317454 435922 317522 435978
rect 317578 435922 348118 435978
rect 348174 435922 348242 435978
rect 348298 435922 378838 435978
rect 378894 435922 378962 435978
rect 379018 435922 409558 435978
rect 409614 435922 409682 435978
rect 409738 435922 440278 435978
rect 440334 435922 440402 435978
rect 440458 435922 470998 435978
rect 471054 435922 471122 435978
rect 471178 435922 501718 435978
rect 501774 435922 501842 435978
rect 501898 435922 532438 435978
rect 532494 435922 532562 435978
rect 532618 435922 558474 435978
rect 558530 435922 558598 435978
rect 558654 435922 558722 435978
rect 558778 435922 558846 435978
rect 558902 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597980 435978
rect -1916 435826 597980 435922
rect -1916 424350 597980 424446
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 9234 424350
rect 9290 424294 9358 424350
rect 9414 424294 9482 424350
rect 9538 424294 9606 424350
rect 9662 424294 39954 424350
rect 40010 424294 40078 424350
rect 40134 424294 40202 424350
rect 40258 424294 40326 424350
rect 40382 424294 70674 424350
rect 70730 424294 70798 424350
rect 70854 424294 70922 424350
rect 70978 424294 71046 424350
rect 71102 424294 101394 424350
rect 101450 424294 101518 424350
rect 101574 424294 101642 424350
rect 101698 424294 101766 424350
rect 101822 424294 132114 424350
rect 132170 424294 132238 424350
rect 132294 424294 132362 424350
rect 132418 424294 132486 424350
rect 132542 424294 162834 424350
rect 162890 424294 162958 424350
rect 163014 424294 163082 424350
rect 163138 424294 163206 424350
rect 163262 424294 209878 424350
rect 209934 424294 210002 424350
rect 210058 424294 240598 424350
rect 240654 424294 240722 424350
rect 240778 424294 271318 424350
rect 271374 424294 271442 424350
rect 271498 424294 302038 424350
rect 302094 424294 302162 424350
rect 302218 424294 332758 424350
rect 332814 424294 332882 424350
rect 332938 424294 363478 424350
rect 363534 424294 363602 424350
rect 363658 424294 394198 424350
rect 394254 424294 394322 424350
rect 394378 424294 424918 424350
rect 424974 424294 425042 424350
rect 425098 424294 455638 424350
rect 455694 424294 455762 424350
rect 455818 424294 486358 424350
rect 486414 424294 486482 424350
rect 486538 424294 517078 424350
rect 517134 424294 517202 424350
rect 517258 424294 547798 424350
rect 547854 424294 547922 424350
rect 547978 424294 562194 424350
rect 562250 424294 562318 424350
rect 562374 424294 562442 424350
rect 562498 424294 562566 424350
rect 562622 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect -1916 424226 597980 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 9234 424226
rect 9290 424170 9358 424226
rect 9414 424170 9482 424226
rect 9538 424170 9606 424226
rect 9662 424170 39954 424226
rect 40010 424170 40078 424226
rect 40134 424170 40202 424226
rect 40258 424170 40326 424226
rect 40382 424170 70674 424226
rect 70730 424170 70798 424226
rect 70854 424170 70922 424226
rect 70978 424170 71046 424226
rect 71102 424170 101394 424226
rect 101450 424170 101518 424226
rect 101574 424170 101642 424226
rect 101698 424170 101766 424226
rect 101822 424170 132114 424226
rect 132170 424170 132238 424226
rect 132294 424170 132362 424226
rect 132418 424170 132486 424226
rect 132542 424170 162834 424226
rect 162890 424170 162958 424226
rect 163014 424170 163082 424226
rect 163138 424170 163206 424226
rect 163262 424170 209878 424226
rect 209934 424170 210002 424226
rect 210058 424170 240598 424226
rect 240654 424170 240722 424226
rect 240778 424170 271318 424226
rect 271374 424170 271442 424226
rect 271498 424170 302038 424226
rect 302094 424170 302162 424226
rect 302218 424170 332758 424226
rect 332814 424170 332882 424226
rect 332938 424170 363478 424226
rect 363534 424170 363602 424226
rect 363658 424170 394198 424226
rect 394254 424170 394322 424226
rect 394378 424170 424918 424226
rect 424974 424170 425042 424226
rect 425098 424170 455638 424226
rect 455694 424170 455762 424226
rect 455818 424170 486358 424226
rect 486414 424170 486482 424226
rect 486538 424170 517078 424226
rect 517134 424170 517202 424226
rect 517258 424170 547798 424226
rect 547854 424170 547922 424226
rect 547978 424170 562194 424226
rect 562250 424170 562318 424226
rect 562374 424170 562442 424226
rect 562498 424170 562566 424226
rect 562622 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect -1916 424102 597980 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 9234 424102
rect 9290 424046 9358 424102
rect 9414 424046 9482 424102
rect 9538 424046 9606 424102
rect 9662 424046 39954 424102
rect 40010 424046 40078 424102
rect 40134 424046 40202 424102
rect 40258 424046 40326 424102
rect 40382 424046 70674 424102
rect 70730 424046 70798 424102
rect 70854 424046 70922 424102
rect 70978 424046 71046 424102
rect 71102 424046 101394 424102
rect 101450 424046 101518 424102
rect 101574 424046 101642 424102
rect 101698 424046 101766 424102
rect 101822 424046 132114 424102
rect 132170 424046 132238 424102
rect 132294 424046 132362 424102
rect 132418 424046 132486 424102
rect 132542 424046 162834 424102
rect 162890 424046 162958 424102
rect 163014 424046 163082 424102
rect 163138 424046 163206 424102
rect 163262 424046 209878 424102
rect 209934 424046 210002 424102
rect 210058 424046 240598 424102
rect 240654 424046 240722 424102
rect 240778 424046 271318 424102
rect 271374 424046 271442 424102
rect 271498 424046 302038 424102
rect 302094 424046 302162 424102
rect 302218 424046 332758 424102
rect 332814 424046 332882 424102
rect 332938 424046 363478 424102
rect 363534 424046 363602 424102
rect 363658 424046 394198 424102
rect 394254 424046 394322 424102
rect 394378 424046 424918 424102
rect 424974 424046 425042 424102
rect 425098 424046 455638 424102
rect 455694 424046 455762 424102
rect 455818 424046 486358 424102
rect 486414 424046 486482 424102
rect 486538 424046 517078 424102
rect 517134 424046 517202 424102
rect 517258 424046 547798 424102
rect 547854 424046 547922 424102
rect 547978 424046 562194 424102
rect 562250 424046 562318 424102
rect 562374 424046 562442 424102
rect 562498 424046 562566 424102
rect 562622 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect -1916 423978 597980 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 9234 423978
rect 9290 423922 9358 423978
rect 9414 423922 9482 423978
rect 9538 423922 9606 423978
rect 9662 423922 39954 423978
rect 40010 423922 40078 423978
rect 40134 423922 40202 423978
rect 40258 423922 40326 423978
rect 40382 423922 70674 423978
rect 70730 423922 70798 423978
rect 70854 423922 70922 423978
rect 70978 423922 71046 423978
rect 71102 423922 101394 423978
rect 101450 423922 101518 423978
rect 101574 423922 101642 423978
rect 101698 423922 101766 423978
rect 101822 423922 132114 423978
rect 132170 423922 132238 423978
rect 132294 423922 132362 423978
rect 132418 423922 132486 423978
rect 132542 423922 162834 423978
rect 162890 423922 162958 423978
rect 163014 423922 163082 423978
rect 163138 423922 163206 423978
rect 163262 423922 209878 423978
rect 209934 423922 210002 423978
rect 210058 423922 240598 423978
rect 240654 423922 240722 423978
rect 240778 423922 271318 423978
rect 271374 423922 271442 423978
rect 271498 423922 302038 423978
rect 302094 423922 302162 423978
rect 302218 423922 332758 423978
rect 332814 423922 332882 423978
rect 332938 423922 363478 423978
rect 363534 423922 363602 423978
rect 363658 423922 394198 423978
rect 394254 423922 394322 423978
rect 394378 423922 424918 423978
rect 424974 423922 425042 423978
rect 425098 423922 455638 423978
rect 455694 423922 455762 423978
rect 455818 423922 486358 423978
rect 486414 423922 486482 423978
rect 486538 423922 517078 423978
rect 517134 423922 517202 423978
rect 517258 423922 547798 423978
rect 547854 423922 547922 423978
rect 547978 423922 562194 423978
rect 562250 423922 562318 423978
rect 562374 423922 562442 423978
rect 562498 423922 562566 423978
rect 562622 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect -1916 423826 597980 423922
rect -1916 418350 597980 418446
rect -1916 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 36234 418350
rect 36290 418294 36358 418350
rect 36414 418294 36482 418350
rect 36538 418294 36606 418350
rect 36662 418294 66954 418350
rect 67010 418294 67078 418350
rect 67134 418294 67202 418350
rect 67258 418294 67326 418350
rect 67382 418294 97674 418350
rect 97730 418294 97798 418350
rect 97854 418294 97922 418350
rect 97978 418294 98046 418350
rect 98102 418294 128394 418350
rect 128450 418294 128518 418350
rect 128574 418294 128642 418350
rect 128698 418294 128766 418350
rect 128822 418294 159114 418350
rect 159170 418294 159238 418350
rect 159294 418294 159362 418350
rect 159418 418294 159486 418350
rect 159542 418294 189834 418350
rect 189890 418294 189958 418350
rect 190014 418294 190082 418350
rect 190138 418294 190206 418350
rect 190262 418294 194518 418350
rect 194574 418294 194642 418350
rect 194698 418294 225238 418350
rect 225294 418294 225362 418350
rect 225418 418294 255958 418350
rect 256014 418294 256082 418350
rect 256138 418294 286678 418350
rect 286734 418294 286802 418350
rect 286858 418294 317398 418350
rect 317454 418294 317522 418350
rect 317578 418294 348118 418350
rect 348174 418294 348242 418350
rect 348298 418294 378838 418350
rect 378894 418294 378962 418350
rect 379018 418294 409558 418350
rect 409614 418294 409682 418350
rect 409738 418294 440278 418350
rect 440334 418294 440402 418350
rect 440458 418294 470998 418350
rect 471054 418294 471122 418350
rect 471178 418294 501718 418350
rect 501774 418294 501842 418350
rect 501898 418294 532438 418350
rect 532494 418294 532562 418350
rect 532618 418294 558474 418350
rect 558530 418294 558598 418350
rect 558654 418294 558722 418350
rect 558778 418294 558846 418350
rect 558902 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597980 418350
rect -1916 418226 597980 418294
rect -1916 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 36234 418226
rect 36290 418170 36358 418226
rect 36414 418170 36482 418226
rect 36538 418170 36606 418226
rect 36662 418170 66954 418226
rect 67010 418170 67078 418226
rect 67134 418170 67202 418226
rect 67258 418170 67326 418226
rect 67382 418170 97674 418226
rect 97730 418170 97798 418226
rect 97854 418170 97922 418226
rect 97978 418170 98046 418226
rect 98102 418170 128394 418226
rect 128450 418170 128518 418226
rect 128574 418170 128642 418226
rect 128698 418170 128766 418226
rect 128822 418170 159114 418226
rect 159170 418170 159238 418226
rect 159294 418170 159362 418226
rect 159418 418170 159486 418226
rect 159542 418170 189834 418226
rect 189890 418170 189958 418226
rect 190014 418170 190082 418226
rect 190138 418170 190206 418226
rect 190262 418170 194518 418226
rect 194574 418170 194642 418226
rect 194698 418170 225238 418226
rect 225294 418170 225362 418226
rect 225418 418170 255958 418226
rect 256014 418170 256082 418226
rect 256138 418170 286678 418226
rect 286734 418170 286802 418226
rect 286858 418170 317398 418226
rect 317454 418170 317522 418226
rect 317578 418170 348118 418226
rect 348174 418170 348242 418226
rect 348298 418170 378838 418226
rect 378894 418170 378962 418226
rect 379018 418170 409558 418226
rect 409614 418170 409682 418226
rect 409738 418170 440278 418226
rect 440334 418170 440402 418226
rect 440458 418170 470998 418226
rect 471054 418170 471122 418226
rect 471178 418170 501718 418226
rect 501774 418170 501842 418226
rect 501898 418170 532438 418226
rect 532494 418170 532562 418226
rect 532618 418170 558474 418226
rect 558530 418170 558598 418226
rect 558654 418170 558722 418226
rect 558778 418170 558846 418226
rect 558902 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597980 418226
rect -1916 418102 597980 418170
rect -1916 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 36234 418102
rect 36290 418046 36358 418102
rect 36414 418046 36482 418102
rect 36538 418046 36606 418102
rect 36662 418046 66954 418102
rect 67010 418046 67078 418102
rect 67134 418046 67202 418102
rect 67258 418046 67326 418102
rect 67382 418046 97674 418102
rect 97730 418046 97798 418102
rect 97854 418046 97922 418102
rect 97978 418046 98046 418102
rect 98102 418046 128394 418102
rect 128450 418046 128518 418102
rect 128574 418046 128642 418102
rect 128698 418046 128766 418102
rect 128822 418046 159114 418102
rect 159170 418046 159238 418102
rect 159294 418046 159362 418102
rect 159418 418046 159486 418102
rect 159542 418046 189834 418102
rect 189890 418046 189958 418102
rect 190014 418046 190082 418102
rect 190138 418046 190206 418102
rect 190262 418046 194518 418102
rect 194574 418046 194642 418102
rect 194698 418046 225238 418102
rect 225294 418046 225362 418102
rect 225418 418046 255958 418102
rect 256014 418046 256082 418102
rect 256138 418046 286678 418102
rect 286734 418046 286802 418102
rect 286858 418046 317398 418102
rect 317454 418046 317522 418102
rect 317578 418046 348118 418102
rect 348174 418046 348242 418102
rect 348298 418046 378838 418102
rect 378894 418046 378962 418102
rect 379018 418046 409558 418102
rect 409614 418046 409682 418102
rect 409738 418046 440278 418102
rect 440334 418046 440402 418102
rect 440458 418046 470998 418102
rect 471054 418046 471122 418102
rect 471178 418046 501718 418102
rect 501774 418046 501842 418102
rect 501898 418046 532438 418102
rect 532494 418046 532562 418102
rect 532618 418046 558474 418102
rect 558530 418046 558598 418102
rect 558654 418046 558722 418102
rect 558778 418046 558846 418102
rect 558902 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597980 418102
rect -1916 417978 597980 418046
rect -1916 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 36234 417978
rect 36290 417922 36358 417978
rect 36414 417922 36482 417978
rect 36538 417922 36606 417978
rect 36662 417922 66954 417978
rect 67010 417922 67078 417978
rect 67134 417922 67202 417978
rect 67258 417922 67326 417978
rect 67382 417922 97674 417978
rect 97730 417922 97798 417978
rect 97854 417922 97922 417978
rect 97978 417922 98046 417978
rect 98102 417922 128394 417978
rect 128450 417922 128518 417978
rect 128574 417922 128642 417978
rect 128698 417922 128766 417978
rect 128822 417922 159114 417978
rect 159170 417922 159238 417978
rect 159294 417922 159362 417978
rect 159418 417922 159486 417978
rect 159542 417922 189834 417978
rect 189890 417922 189958 417978
rect 190014 417922 190082 417978
rect 190138 417922 190206 417978
rect 190262 417922 194518 417978
rect 194574 417922 194642 417978
rect 194698 417922 225238 417978
rect 225294 417922 225362 417978
rect 225418 417922 255958 417978
rect 256014 417922 256082 417978
rect 256138 417922 286678 417978
rect 286734 417922 286802 417978
rect 286858 417922 317398 417978
rect 317454 417922 317522 417978
rect 317578 417922 348118 417978
rect 348174 417922 348242 417978
rect 348298 417922 378838 417978
rect 378894 417922 378962 417978
rect 379018 417922 409558 417978
rect 409614 417922 409682 417978
rect 409738 417922 440278 417978
rect 440334 417922 440402 417978
rect 440458 417922 470998 417978
rect 471054 417922 471122 417978
rect 471178 417922 501718 417978
rect 501774 417922 501842 417978
rect 501898 417922 532438 417978
rect 532494 417922 532562 417978
rect 532618 417922 558474 417978
rect 558530 417922 558598 417978
rect 558654 417922 558722 417978
rect 558778 417922 558846 417978
rect 558902 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597980 417978
rect -1916 417826 597980 417922
rect 57916 409258 308100 409274
rect 57916 409202 57932 409258
rect 57988 409202 308028 409258
rect 308084 409202 308100 409258
rect 57916 409186 308100 409202
rect 7516 409078 302724 409094
rect 7516 409022 7532 409078
rect 7588 409022 302652 409078
rect 302708 409022 302724 409078
rect 7516 409006 302724 409022
rect 245180 407638 477220 407654
rect 245180 407582 245196 407638
rect 245252 407582 477148 407638
rect 477204 407582 477220 407638
rect 245180 407566 477220 407582
rect 238124 407458 475540 407474
rect 238124 407402 238140 407458
rect 238196 407402 475468 407458
rect 475524 407402 475540 407458
rect 238124 407386 475540 407402
rect -1916 406350 597980 406446
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 9234 406350
rect 9290 406294 9358 406350
rect 9414 406294 9482 406350
rect 9538 406294 9606 406350
rect 9662 406294 39954 406350
rect 40010 406294 40078 406350
rect 40134 406294 40202 406350
rect 40258 406294 40326 406350
rect 40382 406294 70674 406350
rect 70730 406294 70798 406350
rect 70854 406294 70922 406350
rect 70978 406294 71046 406350
rect 71102 406294 101394 406350
rect 101450 406294 101518 406350
rect 101574 406294 101642 406350
rect 101698 406294 101766 406350
rect 101822 406294 132114 406350
rect 132170 406294 132238 406350
rect 132294 406294 132362 406350
rect 132418 406294 132486 406350
rect 132542 406294 162834 406350
rect 162890 406294 162958 406350
rect 163014 406294 163082 406350
rect 163138 406294 163206 406350
rect 163262 406294 193554 406350
rect 193610 406294 193678 406350
rect 193734 406294 193802 406350
rect 193858 406294 193926 406350
rect 193982 406294 224274 406350
rect 224330 406294 224398 406350
rect 224454 406294 224522 406350
rect 224578 406294 224646 406350
rect 224702 406294 254994 406350
rect 255050 406294 255118 406350
rect 255174 406294 255242 406350
rect 255298 406294 255366 406350
rect 255422 406294 285714 406350
rect 285770 406294 285838 406350
rect 285894 406294 285962 406350
rect 286018 406294 286086 406350
rect 286142 406294 316434 406350
rect 316490 406294 316558 406350
rect 316614 406294 316682 406350
rect 316738 406294 316806 406350
rect 316862 406294 347154 406350
rect 347210 406294 347278 406350
rect 347334 406294 347402 406350
rect 347458 406294 347526 406350
rect 347582 406294 377874 406350
rect 377930 406294 377998 406350
rect 378054 406294 378122 406350
rect 378178 406294 378246 406350
rect 378302 406294 408594 406350
rect 408650 406294 408718 406350
rect 408774 406294 408842 406350
rect 408898 406294 408966 406350
rect 409022 406294 439314 406350
rect 439370 406294 439438 406350
rect 439494 406294 439562 406350
rect 439618 406294 439686 406350
rect 439742 406294 470034 406350
rect 470090 406294 470158 406350
rect 470214 406294 470282 406350
rect 470338 406294 470406 406350
rect 470462 406294 500754 406350
rect 500810 406294 500878 406350
rect 500934 406294 501002 406350
rect 501058 406294 501126 406350
rect 501182 406294 531474 406350
rect 531530 406294 531598 406350
rect 531654 406294 531722 406350
rect 531778 406294 531846 406350
rect 531902 406294 562194 406350
rect 562250 406294 562318 406350
rect 562374 406294 562442 406350
rect 562498 406294 562566 406350
rect 562622 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect -1916 406226 597980 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 9234 406226
rect 9290 406170 9358 406226
rect 9414 406170 9482 406226
rect 9538 406170 9606 406226
rect 9662 406170 39954 406226
rect 40010 406170 40078 406226
rect 40134 406170 40202 406226
rect 40258 406170 40326 406226
rect 40382 406170 70674 406226
rect 70730 406170 70798 406226
rect 70854 406170 70922 406226
rect 70978 406170 71046 406226
rect 71102 406170 101394 406226
rect 101450 406170 101518 406226
rect 101574 406170 101642 406226
rect 101698 406170 101766 406226
rect 101822 406170 132114 406226
rect 132170 406170 132238 406226
rect 132294 406170 132362 406226
rect 132418 406170 132486 406226
rect 132542 406170 162834 406226
rect 162890 406170 162958 406226
rect 163014 406170 163082 406226
rect 163138 406170 163206 406226
rect 163262 406170 193554 406226
rect 193610 406170 193678 406226
rect 193734 406170 193802 406226
rect 193858 406170 193926 406226
rect 193982 406170 224274 406226
rect 224330 406170 224398 406226
rect 224454 406170 224522 406226
rect 224578 406170 224646 406226
rect 224702 406170 254994 406226
rect 255050 406170 255118 406226
rect 255174 406170 255242 406226
rect 255298 406170 255366 406226
rect 255422 406170 285714 406226
rect 285770 406170 285838 406226
rect 285894 406170 285962 406226
rect 286018 406170 286086 406226
rect 286142 406170 316434 406226
rect 316490 406170 316558 406226
rect 316614 406170 316682 406226
rect 316738 406170 316806 406226
rect 316862 406170 347154 406226
rect 347210 406170 347278 406226
rect 347334 406170 347402 406226
rect 347458 406170 347526 406226
rect 347582 406170 377874 406226
rect 377930 406170 377998 406226
rect 378054 406170 378122 406226
rect 378178 406170 378246 406226
rect 378302 406170 408594 406226
rect 408650 406170 408718 406226
rect 408774 406170 408842 406226
rect 408898 406170 408966 406226
rect 409022 406170 439314 406226
rect 439370 406170 439438 406226
rect 439494 406170 439562 406226
rect 439618 406170 439686 406226
rect 439742 406170 470034 406226
rect 470090 406170 470158 406226
rect 470214 406170 470282 406226
rect 470338 406170 470406 406226
rect 470462 406170 500754 406226
rect 500810 406170 500878 406226
rect 500934 406170 501002 406226
rect 501058 406170 501126 406226
rect 501182 406170 531474 406226
rect 531530 406170 531598 406226
rect 531654 406170 531722 406226
rect 531778 406170 531846 406226
rect 531902 406170 562194 406226
rect 562250 406170 562318 406226
rect 562374 406170 562442 406226
rect 562498 406170 562566 406226
rect 562622 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect -1916 406102 597980 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 9234 406102
rect 9290 406046 9358 406102
rect 9414 406046 9482 406102
rect 9538 406046 9606 406102
rect 9662 406046 39954 406102
rect 40010 406046 40078 406102
rect 40134 406046 40202 406102
rect 40258 406046 40326 406102
rect 40382 406046 70674 406102
rect 70730 406046 70798 406102
rect 70854 406046 70922 406102
rect 70978 406046 71046 406102
rect 71102 406046 101394 406102
rect 101450 406046 101518 406102
rect 101574 406046 101642 406102
rect 101698 406046 101766 406102
rect 101822 406046 132114 406102
rect 132170 406046 132238 406102
rect 132294 406046 132362 406102
rect 132418 406046 132486 406102
rect 132542 406046 162834 406102
rect 162890 406046 162958 406102
rect 163014 406046 163082 406102
rect 163138 406046 163206 406102
rect 163262 406046 193554 406102
rect 193610 406046 193678 406102
rect 193734 406046 193802 406102
rect 193858 406046 193926 406102
rect 193982 406046 224274 406102
rect 224330 406046 224398 406102
rect 224454 406046 224522 406102
rect 224578 406046 224646 406102
rect 224702 406046 254994 406102
rect 255050 406046 255118 406102
rect 255174 406046 255242 406102
rect 255298 406046 255366 406102
rect 255422 406046 285714 406102
rect 285770 406046 285838 406102
rect 285894 406046 285962 406102
rect 286018 406046 286086 406102
rect 286142 406046 316434 406102
rect 316490 406046 316558 406102
rect 316614 406046 316682 406102
rect 316738 406046 316806 406102
rect 316862 406046 347154 406102
rect 347210 406046 347278 406102
rect 347334 406046 347402 406102
rect 347458 406046 347526 406102
rect 347582 406046 377874 406102
rect 377930 406046 377998 406102
rect 378054 406046 378122 406102
rect 378178 406046 378246 406102
rect 378302 406046 408594 406102
rect 408650 406046 408718 406102
rect 408774 406046 408842 406102
rect 408898 406046 408966 406102
rect 409022 406046 439314 406102
rect 439370 406046 439438 406102
rect 439494 406046 439562 406102
rect 439618 406046 439686 406102
rect 439742 406046 470034 406102
rect 470090 406046 470158 406102
rect 470214 406046 470282 406102
rect 470338 406046 470406 406102
rect 470462 406046 500754 406102
rect 500810 406046 500878 406102
rect 500934 406046 501002 406102
rect 501058 406046 501126 406102
rect 501182 406046 531474 406102
rect 531530 406046 531598 406102
rect 531654 406046 531722 406102
rect 531778 406046 531846 406102
rect 531902 406046 562194 406102
rect 562250 406046 562318 406102
rect 562374 406046 562442 406102
rect 562498 406046 562566 406102
rect 562622 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect -1916 405978 597980 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 9234 405978
rect 9290 405922 9358 405978
rect 9414 405922 9482 405978
rect 9538 405922 9606 405978
rect 9662 405922 39954 405978
rect 40010 405922 40078 405978
rect 40134 405922 40202 405978
rect 40258 405922 40326 405978
rect 40382 405922 70674 405978
rect 70730 405922 70798 405978
rect 70854 405922 70922 405978
rect 70978 405922 71046 405978
rect 71102 405922 101394 405978
rect 101450 405922 101518 405978
rect 101574 405922 101642 405978
rect 101698 405922 101766 405978
rect 101822 405922 132114 405978
rect 132170 405922 132238 405978
rect 132294 405922 132362 405978
rect 132418 405922 132486 405978
rect 132542 405922 162834 405978
rect 162890 405922 162958 405978
rect 163014 405922 163082 405978
rect 163138 405922 163206 405978
rect 163262 405922 193554 405978
rect 193610 405922 193678 405978
rect 193734 405922 193802 405978
rect 193858 405922 193926 405978
rect 193982 405922 224274 405978
rect 224330 405922 224398 405978
rect 224454 405922 224522 405978
rect 224578 405922 224646 405978
rect 224702 405922 254994 405978
rect 255050 405922 255118 405978
rect 255174 405922 255242 405978
rect 255298 405922 255366 405978
rect 255422 405922 285714 405978
rect 285770 405922 285838 405978
rect 285894 405922 285962 405978
rect 286018 405922 286086 405978
rect 286142 405922 316434 405978
rect 316490 405922 316558 405978
rect 316614 405922 316682 405978
rect 316738 405922 316806 405978
rect 316862 405922 347154 405978
rect 347210 405922 347278 405978
rect 347334 405922 347402 405978
rect 347458 405922 347526 405978
rect 347582 405922 377874 405978
rect 377930 405922 377998 405978
rect 378054 405922 378122 405978
rect 378178 405922 378246 405978
rect 378302 405922 408594 405978
rect 408650 405922 408718 405978
rect 408774 405922 408842 405978
rect 408898 405922 408966 405978
rect 409022 405922 439314 405978
rect 439370 405922 439438 405978
rect 439494 405922 439562 405978
rect 439618 405922 439686 405978
rect 439742 405922 470034 405978
rect 470090 405922 470158 405978
rect 470214 405922 470282 405978
rect 470338 405922 470406 405978
rect 470462 405922 500754 405978
rect 500810 405922 500878 405978
rect 500934 405922 501002 405978
rect 501058 405922 501126 405978
rect 501182 405922 531474 405978
rect 531530 405922 531598 405978
rect 531654 405922 531722 405978
rect 531778 405922 531846 405978
rect 531902 405922 562194 405978
rect 562250 405922 562318 405978
rect 562374 405922 562442 405978
rect 562498 405922 562566 405978
rect 562622 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect -1916 405826 597980 405922
rect 231740 404038 590900 404054
rect 231740 403982 231756 404038
rect 231812 403982 590828 404038
rect 590884 403982 590900 404038
rect 231740 403966 590900 403982
rect -1916 400350 597980 400446
rect -1916 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 36234 400350
rect 36290 400294 36358 400350
rect 36414 400294 36482 400350
rect 36538 400294 36606 400350
rect 36662 400294 66954 400350
rect 67010 400294 67078 400350
rect 67134 400294 67202 400350
rect 67258 400294 67326 400350
rect 67382 400294 97674 400350
rect 97730 400294 97798 400350
rect 97854 400294 97922 400350
rect 97978 400294 98046 400350
rect 98102 400294 128394 400350
rect 128450 400294 128518 400350
rect 128574 400294 128642 400350
rect 128698 400294 128766 400350
rect 128822 400294 159114 400350
rect 159170 400294 159238 400350
rect 159294 400294 159362 400350
rect 159418 400294 159486 400350
rect 159542 400294 189834 400350
rect 189890 400294 189958 400350
rect 190014 400294 190082 400350
rect 190138 400294 190206 400350
rect 190262 400294 220554 400350
rect 220610 400294 220678 400350
rect 220734 400294 220802 400350
rect 220858 400294 220926 400350
rect 220982 400294 404874 400350
rect 404930 400294 404998 400350
rect 405054 400294 405122 400350
rect 405178 400294 405246 400350
rect 405302 400294 435594 400350
rect 435650 400294 435718 400350
rect 435774 400294 435842 400350
rect 435898 400294 435966 400350
rect 436022 400294 466314 400350
rect 466370 400294 466438 400350
rect 466494 400294 466562 400350
rect 466618 400294 466686 400350
rect 466742 400294 497034 400350
rect 497090 400294 497158 400350
rect 497214 400294 497282 400350
rect 497338 400294 497406 400350
rect 497462 400294 527754 400350
rect 527810 400294 527878 400350
rect 527934 400294 528002 400350
rect 528058 400294 528126 400350
rect 528182 400294 558474 400350
rect 558530 400294 558598 400350
rect 558654 400294 558722 400350
rect 558778 400294 558846 400350
rect 558902 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597980 400350
rect -1916 400226 597980 400294
rect -1916 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 36234 400226
rect 36290 400170 36358 400226
rect 36414 400170 36482 400226
rect 36538 400170 36606 400226
rect 36662 400170 66954 400226
rect 67010 400170 67078 400226
rect 67134 400170 67202 400226
rect 67258 400170 67326 400226
rect 67382 400170 97674 400226
rect 97730 400170 97798 400226
rect 97854 400170 97922 400226
rect 97978 400170 98046 400226
rect 98102 400170 128394 400226
rect 128450 400170 128518 400226
rect 128574 400170 128642 400226
rect 128698 400170 128766 400226
rect 128822 400170 159114 400226
rect 159170 400170 159238 400226
rect 159294 400170 159362 400226
rect 159418 400170 159486 400226
rect 159542 400170 189834 400226
rect 189890 400170 189958 400226
rect 190014 400170 190082 400226
rect 190138 400170 190206 400226
rect 190262 400170 220554 400226
rect 220610 400170 220678 400226
rect 220734 400170 220802 400226
rect 220858 400170 220926 400226
rect 220982 400170 404874 400226
rect 404930 400170 404998 400226
rect 405054 400170 405122 400226
rect 405178 400170 405246 400226
rect 405302 400170 435594 400226
rect 435650 400170 435718 400226
rect 435774 400170 435842 400226
rect 435898 400170 435966 400226
rect 436022 400170 466314 400226
rect 466370 400170 466438 400226
rect 466494 400170 466562 400226
rect 466618 400170 466686 400226
rect 466742 400170 497034 400226
rect 497090 400170 497158 400226
rect 497214 400170 497282 400226
rect 497338 400170 497406 400226
rect 497462 400170 527754 400226
rect 527810 400170 527878 400226
rect 527934 400170 528002 400226
rect 528058 400170 528126 400226
rect 528182 400170 558474 400226
rect 558530 400170 558598 400226
rect 558654 400170 558722 400226
rect 558778 400170 558846 400226
rect 558902 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597980 400226
rect -1916 400102 597980 400170
rect -1916 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 36234 400102
rect 36290 400046 36358 400102
rect 36414 400046 36482 400102
rect 36538 400046 36606 400102
rect 36662 400046 66954 400102
rect 67010 400046 67078 400102
rect 67134 400046 67202 400102
rect 67258 400046 67326 400102
rect 67382 400046 97674 400102
rect 97730 400046 97798 400102
rect 97854 400046 97922 400102
rect 97978 400046 98046 400102
rect 98102 400046 128394 400102
rect 128450 400046 128518 400102
rect 128574 400046 128642 400102
rect 128698 400046 128766 400102
rect 128822 400046 159114 400102
rect 159170 400046 159238 400102
rect 159294 400046 159362 400102
rect 159418 400046 159486 400102
rect 159542 400046 189834 400102
rect 189890 400046 189958 400102
rect 190014 400046 190082 400102
rect 190138 400046 190206 400102
rect 190262 400046 220554 400102
rect 220610 400046 220678 400102
rect 220734 400046 220802 400102
rect 220858 400046 220926 400102
rect 220982 400046 404874 400102
rect 404930 400046 404998 400102
rect 405054 400046 405122 400102
rect 405178 400046 405246 400102
rect 405302 400046 435594 400102
rect 435650 400046 435718 400102
rect 435774 400046 435842 400102
rect 435898 400046 435966 400102
rect 436022 400046 466314 400102
rect 466370 400046 466438 400102
rect 466494 400046 466562 400102
rect 466618 400046 466686 400102
rect 466742 400046 497034 400102
rect 497090 400046 497158 400102
rect 497214 400046 497282 400102
rect 497338 400046 497406 400102
rect 497462 400046 527754 400102
rect 527810 400046 527878 400102
rect 527934 400046 528002 400102
rect 528058 400046 528126 400102
rect 528182 400046 558474 400102
rect 558530 400046 558598 400102
rect 558654 400046 558722 400102
rect 558778 400046 558846 400102
rect 558902 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597980 400102
rect -1916 399978 597980 400046
rect -1916 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 36234 399978
rect 36290 399922 36358 399978
rect 36414 399922 36482 399978
rect 36538 399922 36606 399978
rect 36662 399922 66954 399978
rect 67010 399922 67078 399978
rect 67134 399922 67202 399978
rect 67258 399922 67326 399978
rect 67382 399922 97674 399978
rect 97730 399922 97798 399978
rect 97854 399922 97922 399978
rect 97978 399922 98046 399978
rect 98102 399922 128394 399978
rect 128450 399922 128518 399978
rect 128574 399922 128642 399978
rect 128698 399922 128766 399978
rect 128822 399922 159114 399978
rect 159170 399922 159238 399978
rect 159294 399922 159362 399978
rect 159418 399922 159486 399978
rect 159542 399922 189834 399978
rect 189890 399922 189958 399978
rect 190014 399922 190082 399978
rect 190138 399922 190206 399978
rect 190262 399922 220554 399978
rect 220610 399922 220678 399978
rect 220734 399922 220802 399978
rect 220858 399922 220926 399978
rect 220982 399922 404874 399978
rect 404930 399922 404998 399978
rect 405054 399922 405122 399978
rect 405178 399922 405246 399978
rect 405302 399922 435594 399978
rect 435650 399922 435718 399978
rect 435774 399922 435842 399978
rect 435898 399922 435966 399978
rect 436022 399922 466314 399978
rect 466370 399922 466438 399978
rect 466494 399922 466562 399978
rect 466618 399922 466686 399978
rect 466742 399922 497034 399978
rect 497090 399922 497158 399978
rect 497214 399922 497282 399978
rect 497338 399922 497406 399978
rect 497462 399922 527754 399978
rect 527810 399922 527878 399978
rect 527934 399922 528002 399978
rect 528058 399922 528126 399978
rect 528182 399922 558474 399978
rect 558530 399922 558598 399978
rect 558654 399922 558722 399978
rect 558778 399922 558846 399978
rect 558902 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597980 399978
rect -1916 399826 597980 399922
rect 238236 389818 577124 389834
rect 238236 389762 238252 389818
rect 238308 389762 577052 389818
rect 577108 389762 577124 389818
rect 238236 389746 577124 389762
rect 212476 388918 297460 388934
rect 212476 388862 212492 388918
rect 212548 388862 297388 388918
rect 297444 388862 297460 388918
rect 212476 388846 297460 388862
rect 282140 388738 384036 388754
rect 282140 388682 282156 388738
rect 282212 388682 383964 388738
rect 384020 388682 384036 388738
rect 282140 388666 384036 388682
rect -1916 388350 597980 388446
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 9234 388350
rect 9290 388294 9358 388350
rect 9414 388294 9482 388350
rect 9538 388294 9606 388350
rect 9662 388294 39954 388350
rect 40010 388294 40078 388350
rect 40134 388294 40202 388350
rect 40258 388294 40326 388350
rect 40382 388294 70674 388350
rect 70730 388294 70798 388350
rect 70854 388294 70922 388350
rect 70978 388294 71046 388350
rect 71102 388294 101394 388350
rect 101450 388294 101518 388350
rect 101574 388294 101642 388350
rect 101698 388294 101766 388350
rect 101822 388294 132114 388350
rect 132170 388294 132238 388350
rect 132294 388294 132362 388350
rect 132418 388294 132486 388350
rect 132542 388294 162834 388350
rect 162890 388294 162958 388350
rect 163014 388294 163082 388350
rect 163138 388294 163206 388350
rect 163262 388294 193554 388350
rect 193610 388294 193678 388350
rect 193734 388294 193802 388350
rect 193858 388294 193926 388350
rect 193982 388294 224274 388350
rect 224330 388294 224398 388350
rect 224454 388294 224522 388350
rect 224578 388294 224646 388350
rect 224702 388294 254994 388350
rect 255050 388294 255118 388350
rect 255174 388294 255242 388350
rect 255298 388294 255366 388350
rect 255422 388294 285714 388350
rect 285770 388294 285838 388350
rect 285894 388294 285962 388350
rect 286018 388294 286086 388350
rect 286142 388294 316434 388350
rect 316490 388294 316558 388350
rect 316614 388294 316682 388350
rect 316738 388294 316806 388350
rect 316862 388294 347154 388350
rect 347210 388294 347278 388350
rect 347334 388294 347402 388350
rect 347458 388294 347526 388350
rect 347582 388294 377874 388350
rect 377930 388294 377998 388350
rect 378054 388294 378122 388350
rect 378178 388294 378246 388350
rect 378302 388294 408594 388350
rect 408650 388294 408718 388350
rect 408774 388294 408842 388350
rect 408898 388294 408966 388350
rect 409022 388294 439314 388350
rect 439370 388294 439438 388350
rect 439494 388294 439562 388350
rect 439618 388294 439686 388350
rect 439742 388294 470034 388350
rect 470090 388294 470158 388350
rect 470214 388294 470282 388350
rect 470338 388294 470406 388350
rect 470462 388294 500754 388350
rect 500810 388294 500878 388350
rect 500934 388294 501002 388350
rect 501058 388294 501126 388350
rect 501182 388294 531474 388350
rect 531530 388294 531598 388350
rect 531654 388294 531722 388350
rect 531778 388294 531846 388350
rect 531902 388294 562194 388350
rect 562250 388294 562318 388350
rect 562374 388294 562442 388350
rect 562498 388294 562566 388350
rect 562622 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect -1916 388226 597980 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 9234 388226
rect 9290 388170 9358 388226
rect 9414 388170 9482 388226
rect 9538 388170 9606 388226
rect 9662 388170 39954 388226
rect 40010 388170 40078 388226
rect 40134 388170 40202 388226
rect 40258 388170 40326 388226
rect 40382 388170 70674 388226
rect 70730 388170 70798 388226
rect 70854 388170 70922 388226
rect 70978 388170 71046 388226
rect 71102 388170 101394 388226
rect 101450 388170 101518 388226
rect 101574 388170 101642 388226
rect 101698 388170 101766 388226
rect 101822 388170 132114 388226
rect 132170 388170 132238 388226
rect 132294 388170 132362 388226
rect 132418 388170 132486 388226
rect 132542 388170 162834 388226
rect 162890 388170 162958 388226
rect 163014 388170 163082 388226
rect 163138 388170 163206 388226
rect 163262 388170 193554 388226
rect 193610 388170 193678 388226
rect 193734 388170 193802 388226
rect 193858 388170 193926 388226
rect 193982 388170 224274 388226
rect 224330 388170 224398 388226
rect 224454 388170 224522 388226
rect 224578 388170 224646 388226
rect 224702 388170 254994 388226
rect 255050 388170 255118 388226
rect 255174 388170 255242 388226
rect 255298 388170 255366 388226
rect 255422 388170 285714 388226
rect 285770 388170 285838 388226
rect 285894 388170 285962 388226
rect 286018 388170 286086 388226
rect 286142 388170 316434 388226
rect 316490 388170 316558 388226
rect 316614 388170 316682 388226
rect 316738 388170 316806 388226
rect 316862 388170 347154 388226
rect 347210 388170 347278 388226
rect 347334 388170 347402 388226
rect 347458 388170 347526 388226
rect 347582 388170 377874 388226
rect 377930 388170 377998 388226
rect 378054 388170 378122 388226
rect 378178 388170 378246 388226
rect 378302 388170 408594 388226
rect 408650 388170 408718 388226
rect 408774 388170 408842 388226
rect 408898 388170 408966 388226
rect 409022 388170 439314 388226
rect 439370 388170 439438 388226
rect 439494 388170 439562 388226
rect 439618 388170 439686 388226
rect 439742 388170 470034 388226
rect 470090 388170 470158 388226
rect 470214 388170 470282 388226
rect 470338 388170 470406 388226
rect 470462 388170 500754 388226
rect 500810 388170 500878 388226
rect 500934 388170 501002 388226
rect 501058 388170 501126 388226
rect 501182 388170 531474 388226
rect 531530 388170 531598 388226
rect 531654 388170 531722 388226
rect 531778 388170 531846 388226
rect 531902 388170 562194 388226
rect 562250 388170 562318 388226
rect 562374 388170 562442 388226
rect 562498 388170 562566 388226
rect 562622 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect -1916 388102 597980 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 9234 388102
rect 9290 388046 9358 388102
rect 9414 388046 9482 388102
rect 9538 388046 9606 388102
rect 9662 388046 39954 388102
rect 40010 388046 40078 388102
rect 40134 388046 40202 388102
rect 40258 388046 40326 388102
rect 40382 388046 70674 388102
rect 70730 388046 70798 388102
rect 70854 388046 70922 388102
rect 70978 388046 71046 388102
rect 71102 388046 101394 388102
rect 101450 388046 101518 388102
rect 101574 388046 101642 388102
rect 101698 388046 101766 388102
rect 101822 388046 132114 388102
rect 132170 388046 132238 388102
rect 132294 388046 132362 388102
rect 132418 388046 132486 388102
rect 132542 388046 162834 388102
rect 162890 388046 162958 388102
rect 163014 388046 163082 388102
rect 163138 388046 163206 388102
rect 163262 388046 193554 388102
rect 193610 388046 193678 388102
rect 193734 388046 193802 388102
rect 193858 388046 193926 388102
rect 193982 388046 224274 388102
rect 224330 388046 224398 388102
rect 224454 388046 224522 388102
rect 224578 388046 224646 388102
rect 224702 388046 254994 388102
rect 255050 388046 255118 388102
rect 255174 388046 255242 388102
rect 255298 388046 255366 388102
rect 255422 388046 285714 388102
rect 285770 388046 285838 388102
rect 285894 388046 285962 388102
rect 286018 388046 286086 388102
rect 286142 388046 316434 388102
rect 316490 388046 316558 388102
rect 316614 388046 316682 388102
rect 316738 388046 316806 388102
rect 316862 388046 347154 388102
rect 347210 388046 347278 388102
rect 347334 388046 347402 388102
rect 347458 388046 347526 388102
rect 347582 388046 377874 388102
rect 377930 388046 377998 388102
rect 378054 388046 378122 388102
rect 378178 388046 378246 388102
rect 378302 388046 408594 388102
rect 408650 388046 408718 388102
rect 408774 388046 408842 388102
rect 408898 388046 408966 388102
rect 409022 388046 439314 388102
rect 439370 388046 439438 388102
rect 439494 388046 439562 388102
rect 439618 388046 439686 388102
rect 439742 388046 470034 388102
rect 470090 388046 470158 388102
rect 470214 388046 470282 388102
rect 470338 388046 470406 388102
rect 470462 388046 500754 388102
rect 500810 388046 500878 388102
rect 500934 388046 501002 388102
rect 501058 388046 501126 388102
rect 501182 388046 531474 388102
rect 531530 388046 531598 388102
rect 531654 388046 531722 388102
rect 531778 388046 531846 388102
rect 531902 388046 562194 388102
rect 562250 388046 562318 388102
rect 562374 388046 562442 388102
rect 562498 388046 562566 388102
rect 562622 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect -1916 387978 597980 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 9234 387978
rect 9290 387922 9358 387978
rect 9414 387922 9482 387978
rect 9538 387922 9606 387978
rect 9662 387922 39954 387978
rect 40010 387922 40078 387978
rect 40134 387922 40202 387978
rect 40258 387922 40326 387978
rect 40382 387922 70674 387978
rect 70730 387922 70798 387978
rect 70854 387922 70922 387978
rect 70978 387922 71046 387978
rect 71102 387922 101394 387978
rect 101450 387922 101518 387978
rect 101574 387922 101642 387978
rect 101698 387922 101766 387978
rect 101822 387922 132114 387978
rect 132170 387922 132238 387978
rect 132294 387922 132362 387978
rect 132418 387922 132486 387978
rect 132542 387922 162834 387978
rect 162890 387922 162958 387978
rect 163014 387922 163082 387978
rect 163138 387922 163206 387978
rect 163262 387922 193554 387978
rect 193610 387922 193678 387978
rect 193734 387922 193802 387978
rect 193858 387922 193926 387978
rect 193982 387922 224274 387978
rect 224330 387922 224398 387978
rect 224454 387922 224522 387978
rect 224578 387922 224646 387978
rect 224702 387922 254994 387978
rect 255050 387922 255118 387978
rect 255174 387922 255242 387978
rect 255298 387922 255366 387978
rect 255422 387922 285714 387978
rect 285770 387922 285838 387978
rect 285894 387922 285962 387978
rect 286018 387922 286086 387978
rect 286142 387922 316434 387978
rect 316490 387922 316558 387978
rect 316614 387922 316682 387978
rect 316738 387922 316806 387978
rect 316862 387922 347154 387978
rect 347210 387922 347278 387978
rect 347334 387922 347402 387978
rect 347458 387922 347526 387978
rect 347582 387922 377874 387978
rect 377930 387922 377998 387978
rect 378054 387922 378122 387978
rect 378178 387922 378246 387978
rect 378302 387922 408594 387978
rect 408650 387922 408718 387978
rect 408774 387922 408842 387978
rect 408898 387922 408966 387978
rect 409022 387922 439314 387978
rect 439370 387922 439438 387978
rect 439494 387922 439562 387978
rect 439618 387922 439686 387978
rect 439742 387922 470034 387978
rect 470090 387922 470158 387978
rect 470214 387922 470282 387978
rect 470338 387922 470406 387978
rect 470462 387922 500754 387978
rect 500810 387922 500878 387978
rect 500934 387922 501002 387978
rect 501058 387922 501126 387978
rect 501182 387922 531474 387978
rect 531530 387922 531598 387978
rect 531654 387922 531722 387978
rect 531778 387922 531846 387978
rect 531902 387922 562194 387978
rect 562250 387922 562318 387978
rect 562374 387922 562442 387978
rect 562498 387922 562566 387978
rect 562622 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect -1916 387826 597980 387922
rect 237676 385678 286372 385694
rect 237676 385622 237692 385678
rect 237748 385622 286300 385678
rect 286356 385622 286372 385678
rect 237676 385606 286372 385622
rect 303980 385678 373172 385694
rect 303980 385622 303996 385678
rect 304052 385622 373100 385678
rect 373156 385622 373172 385678
rect 303980 385606 373172 385622
rect 7516 385498 267892 385514
rect 7516 385442 7532 385498
rect 7588 385442 267820 385498
rect 267876 385442 267892 385498
rect 7516 385426 267892 385442
rect 273180 385498 583060 385514
rect 273180 385442 273196 385498
rect 273252 385442 582988 385498
rect 583044 385442 583060 385498
rect 273180 385426 583060 385442
rect 27676 385318 269684 385334
rect 27676 385262 27692 385318
rect 27748 385262 269612 385318
rect 269668 385262 269684 385318
rect 27676 385246 269684 385262
rect 271388 385318 579700 385334
rect 271388 385262 271404 385318
rect 271460 385262 579628 385318
rect 579684 385262 579700 385318
rect 271388 385246 579700 385262
rect 287516 384418 464564 384434
rect 287516 384362 287532 384418
rect 287588 384362 464492 384418
rect 464548 384362 464564 384418
rect 287516 384346 464564 384362
rect 288412 384238 476324 384254
rect 288412 384182 288428 384238
rect 288484 384182 476252 384238
rect 476308 384182 476324 384238
rect 288412 384166 476324 384182
rect 290204 384058 479684 384074
rect 290204 384002 290220 384058
rect 290276 384002 479612 384058
rect 479668 384002 479684 384058
rect 290204 383986 479684 384002
rect 289308 383878 481364 383894
rect 289308 383822 289324 383878
rect 289380 383822 481292 383878
rect 481348 383822 481364 383878
rect 289308 383806 481364 383822
rect 235884 382618 520004 382634
rect 235884 382562 235900 382618
rect 235956 382562 519932 382618
rect 519988 382562 520004 382618
rect 235884 382546 520004 382562
rect -1916 382350 597980 382446
rect -1916 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 36234 382350
rect 36290 382294 36358 382350
rect 36414 382294 36482 382350
rect 36538 382294 36606 382350
rect 36662 382294 66954 382350
rect 67010 382294 67078 382350
rect 67134 382294 67202 382350
rect 67258 382294 67326 382350
rect 67382 382294 97674 382350
rect 97730 382294 97798 382350
rect 97854 382294 97922 382350
rect 97978 382294 98046 382350
rect 98102 382294 128394 382350
rect 128450 382294 128518 382350
rect 128574 382294 128642 382350
rect 128698 382294 128766 382350
rect 128822 382294 159114 382350
rect 159170 382294 159238 382350
rect 159294 382294 159362 382350
rect 159418 382294 159486 382350
rect 159542 382294 189834 382350
rect 189890 382294 189958 382350
rect 190014 382294 190082 382350
rect 190138 382294 190206 382350
rect 190262 382294 220554 382350
rect 220610 382294 220678 382350
rect 220734 382294 220802 382350
rect 220858 382294 220926 382350
rect 220982 382294 404874 382350
rect 404930 382294 404998 382350
rect 405054 382294 405122 382350
rect 405178 382294 405246 382350
rect 405302 382294 435594 382350
rect 435650 382294 435718 382350
rect 435774 382294 435842 382350
rect 435898 382294 435966 382350
rect 436022 382294 466314 382350
rect 466370 382294 466438 382350
rect 466494 382294 466562 382350
rect 466618 382294 466686 382350
rect 466742 382294 497034 382350
rect 497090 382294 497158 382350
rect 497214 382294 497282 382350
rect 497338 382294 497406 382350
rect 497462 382294 527754 382350
rect 527810 382294 527878 382350
rect 527934 382294 528002 382350
rect 528058 382294 528126 382350
rect 528182 382294 558474 382350
rect 558530 382294 558598 382350
rect 558654 382294 558722 382350
rect 558778 382294 558846 382350
rect 558902 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597980 382350
rect -1916 382269 597980 382294
rect -1916 382226 240518 382269
rect -1916 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 36234 382226
rect 36290 382170 36358 382226
rect 36414 382170 36482 382226
rect 36538 382170 36606 382226
rect 36662 382170 66954 382226
rect 67010 382170 67078 382226
rect 67134 382170 67202 382226
rect 67258 382170 67326 382226
rect 67382 382170 97674 382226
rect 97730 382170 97798 382226
rect 97854 382170 97922 382226
rect 97978 382170 98046 382226
rect 98102 382170 128394 382226
rect 128450 382170 128518 382226
rect 128574 382170 128642 382226
rect 128698 382170 128766 382226
rect 128822 382170 159114 382226
rect 159170 382170 159238 382226
rect 159294 382170 159362 382226
rect 159418 382170 159486 382226
rect 159542 382170 189834 382226
rect 189890 382170 189958 382226
rect 190014 382170 190082 382226
rect 190138 382170 190206 382226
rect 190262 382170 220554 382226
rect 220610 382170 220678 382226
rect 220734 382170 220802 382226
rect 220858 382170 220926 382226
rect 220982 382213 240518 382226
rect 240574 382213 240642 382269
rect 240698 382213 271238 382269
rect 271294 382213 271362 382269
rect 271418 382213 301958 382269
rect 302014 382213 302082 382269
rect 302138 382213 332678 382269
rect 332734 382213 332802 382269
rect 332858 382213 363398 382269
rect 363454 382213 363522 382269
rect 363578 382226 597980 382269
rect 363578 382213 404874 382226
rect 220982 382170 404874 382213
rect 404930 382170 404998 382226
rect 405054 382170 405122 382226
rect 405178 382170 405246 382226
rect 405302 382170 435594 382226
rect 435650 382170 435718 382226
rect 435774 382170 435842 382226
rect 435898 382170 435966 382226
rect 436022 382170 466314 382226
rect 466370 382170 466438 382226
rect 466494 382170 466562 382226
rect 466618 382170 466686 382226
rect 466742 382170 497034 382226
rect 497090 382170 497158 382226
rect 497214 382170 497282 382226
rect 497338 382170 497406 382226
rect 497462 382170 527754 382226
rect 527810 382170 527878 382226
rect 527934 382170 528002 382226
rect 528058 382170 528126 382226
rect 528182 382170 558474 382226
rect 558530 382170 558598 382226
rect 558654 382170 558722 382226
rect 558778 382170 558846 382226
rect 558902 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597980 382226
rect -1916 382145 597980 382170
rect -1916 382102 240518 382145
rect -1916 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 36234 382102
rect 36290 382046 36358 382102
rect 36414 382046 36482 382102
rect 36538 382046 36606 382102
rect 36662 382046 66954 382102
rect 67010 382046 67078 382102
rect 67134 382046 67202 382102
rect 67258 382046 67326 382102
rect 67382 382046 97674 382102
rect 97730 382046 97798 382102
rect 97854 382046 97922 382102
rect 97978 382046 98046 382102
rect 98102 382046 128394 382102
rect 128450 382046 128518 382102
rect 128574 382046 128642 382102
rect 128698 382046 128766 382102
rect 128822 382046 159114 382102
rect 159170 382046 159238 382102
rect 159294 382046 159362 382102
rect 159418 382046 159486 382102
rect 159542 382046 189834 382102
rect 189890 382046 189958 382102
rect 190014 382046 190082 382102
rect 190138 382046 190206 382102
rect 190262 382046 220554 382102
rect 220610 382046 220678 382102
rect 220734 382046 220802 382102
rect 220858 382046 220926 382102
rect 220982 382089 240518 382102
rect 240574 382089 240642 382145
rect 240698 382089 271238 382145
rect 271294 382089 271362 382145
rect 271418 382089 301958 382145
rect 302014 382089 302082 382145
rect 302138 382089 332678 382145
rect 332734 382089 332802 382145
rect 332858 382089 363398 382145
rect 363454 382089 363522 382145
rect 363578 382102 597980 382145
rect 363578 382089 404874 382102
rect 220982 382046 404874 382089
rect 404930 382046 404998 382102
rect 405054 382046 405122 382102
rect 405178 382046 405246 382102
rect 405302 382046 435594 382102
rect 435650 382046 435718 382102
rect 435774 382046 435842 382102
rect 435898 382046 435966 382102
rect 436022 382046 466314 382102
rect 466370 382046 466438 382102
rect 466494 382046 466562 382102
rect 466618 382046 466686 382102
rect 466742 382046 497034 382102
rect 497090 382046 497158 382102
rect 497214 382046 497282 382102
rect 497338 382046 497406 382102
rect 497462 382046 527754 382102
rect 527810 382046 527878 382102
rect 527934 382046 528002 382102
rect 528058 382046 528126 382102
rect 528182 382046 558474 382102
rect 558530 382046 558598 382102
rect 558654 382046 558722 382102
rect 558778 382046 558846 382102
rect 558902 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597980 382102
rect -1916 382021 597980 382046
rect -1916 381978 240518 382021
rect -1916 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 36234 381978
rect 36290 381922 36358 381978
rect 36414 381922 36482 381978
rect 36538 381922 36606 381978
rect 36662 381922 66954 381978
rect 67010 381922 67078 381978
rect 67134 381922 67202 381978
rect 67258 381922 67326 381978
rect 67382 381922 97674 381978
rect 97730 381922 97798 381978
rect 97854 381922 97922 381978
rect 97978 381922 98046 381978
rect 98102 381922 128394 381978
rect 128450 381922 128518 381978
rect 128574 381922 128642 381978
rect 128698 381922 128766 381978
rect 128822 381922 159114 381978
rect 159170 381922 159238 381978
rect 159294 381922 159362 381978
rect 159418 381922 159486 381978
rect 159542 381922 189834 381978
rect 189890 381922 189958 381978
rect 190014 381922 190082 381978
rect 190138 381922 190206 381978
rect 190262 381922 220554 381978
rect 220610 381922 220678 381978
rect 220734 381922 220802 381978
rect 220858 381922 220926 381978
rect 220982 381965 240518 381978
rect 240574 381965 240642 382021
rect 240698 381965 271238 382021
rect 271294 381965 271362 382021
rect 271418 381965 301958 382021
rect 302014 381965 302082 382021
rect 302138 381965 332678 382021
rect 332734 381965 332802 382021
rect 332858 381965 363398 382021
rect 363454 381965 363522 382021
rect 363578 381978 597980 382021
rect 363578 381965 404874 381978
rect 220982 381922 404874 381965
rect 404930 381922 404998 381978
rect 405054 381922 405122 381978
rect 405178 381922 405246 381978
rect 405302 381922 435594 381978
rect 435650 381922 435718 381978
rect 435774 381922 435842 381978
rect 435898 381922 435966 381978
rect 436022 381922 466314 381978
rect 466370 381922 466438 381978
rect 466494 381922 466562 381978
rect 466618 381922 466686 381978
rect 466742 381922 497034 381978
rect 497090 381922 497158 381978
rect 497214 381922 497282 381978
rect 497338 381922 497406 381978
rect 497462 381922 527754 381978
rect 527810 381922 527878 381978
rect 527934 381922 528002 381978
rect 528058 381922 528126 381978
rect 528182 381922 558474 381978
rect 558530 381922 558598 381978
rect 558654 381922 558722 381978
rect 558778 381922 558846 381978
rect 558902 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597980 381978
rect -1916 381897 597980 381922
rect -1916 381841 240518 381897
rect 240574 381841 240642 381897
rect 240698 381841 271238 381897
rect 271294 381841 271362 381897
rect 271418 381841 301958 381897
rect 302014 381841 302082 381897
rect 302138 381841 332678 381897
rect 332734 381841 332802 381897
rect 332858 381841 363398 381897
rect 363454 381841 363522 381897
rect 363578 381841 597980 381897
rect -1916 381826 597980 381841
rect -1916 370350 597980 370446
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 9234 370350
rect 9290 370294 9358 370350
rect 9414 370294 9482 370350
rect 9538 370294 9606 370350
rect 9662 370294 39954 370350
rect 40010 370294 40078 370350
rect 40134 370294 40202 370350
rect 40258 370294 40326 370350
rect 40382 370294 70674 370350
rect 70730 370294 70798 370350
rect 70854 370294 70922 370350
rect 70978 370294 71046 370350
rect 71102 370294 101394 370350
rect 101450 370294 101518 370350
rect 101574 370294 101642 370350
rect 101698 370294 101766 370350
rect 101822 370294 132114 370350
rect 132170 370294 132238 370350
rect 132294 370294 132362 370350
rect 132418 370294 132486 370350
rect 132542 370294 162834 370350
rect 162890 370294 162958 370350
rect 163014 370294 163082 370350
rect 163138 370294 163206 370350
rect 163262 370294 193554 370350
rect 193610 370294 193678 370350
rect 193734 370294 193802 370350
rect 193858 370294 193926 370350
rect 193982 370294 224274 370350
rect 224330 370294 224398 370350
rect 224454 370294 224522 370350
rect 224578 370294 224646 370350
rect 224702 370294 255878 370350
rect 255934 370294 256002 370350
rect 256058 370294 286598 370350
rect 286654 370294 286722 370350
rect 286778 370294 317318 370350
rect 317374 370294 317442 370350
rect 317498 370294 348038 370350
rect 348094 370294 348162 370350
rect 348218 370294 377874 370350
rect 377930 370294 377998 370350
rect 378054 370294 378122 370350
rect 378178 370294 378246 370350
rect 378302 370294 408594 370350
rect 408650 370294 408718 370350
rect 408774 370294 408842 370350
rect 408898 370294 408966 370350
rect 409022 370294 439314 370350
rect 439370 370294 439438 370350
rect 439494 370294 439562 370350
rect 439618 370294 439686 370350
rect 439742 370294 470034 370350
rect 470090 370294 470158 370350
rect 470214 370294 470282 370350
rect 470338 370294 470406 370350
rect 470462 370294 500754 370350
rect 500810 370294 500878 370350
rect 500934 370294 501002 370350
rect 501058 370294 501126 370350
rect 501182 370294 531474 370350
rect 531530 370294 531598 370350
rect 531654 370294 531722 370350
rect 531778 370294 531846 370350
rect 531902 370294 562194 370350
rect 562250 370294 562318 370350
rect 562374 370294 562442 370350
rect 562498 370294 562566 370350
rect 562622 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect -1916 370226 597980 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 9234 370226
rect 9290 370170 9358 370226
rect 9414 370170 9482 370226
rect 9538 370170 9606 370226
rect 9662 370170 39954 370226
rect 40010 370170 40078 370226
rect 40134 370170 40202 370226
rect 40258 370170 40326 370226
rect 40382 370170 70674 370226
rect 70730 370170 70798 370226
rect 70854 370170 70922 370226
rect 70978 370170 71046 370226
rect 71102 370170 101394 370226
rect 101450 370170 101518 370226
rect 101574 370170 101642 370226
rect 101698 370170 101766 370226
rect 101822 370170 132114 370226
rect 132170 370170 132238 370226
rect 132294 370170 132362 370226
rect 132418 370170 132486 370226
rect 132542 370170 162834 370226
rect 162890 370170 162958 370226
rect 163014 370170 163082 370226
rect 163138 370170 163206 370226
rect 163262 370170 193554 370226
rect 193610 370170 193678 370226
rect 193734 370170 193802 370226
rect 193858 370170 193926 370226
rect 193982 370170 224274 370226
rect 224330 370170 224398 370226
rect 224454 370170 224522 370226
rect 224578 370170 224646 370226
rect 224702 370170 255878 370226
rect 255934 370170 256002 370226
rect 256058 370170 286598 370226
rect 286654 370170 286722 370226
rect 286778 370170 317318 370226
rect 317374 370170 317442 370226
rect 317498 370170 348038 370226
rect 348094 370170 348162 370226
rect 348218 370170 377874 370226
rect 377930 370170 377998 370226
rect 378054 370170 378122 370226
rect 378178 370170 378246 370226
rect 378302 370170 408594 370226
rect 408650 370170 408718 370226
rect 408774 370170 408842 370226
rect 408898 370170 408966 370226
rect 409022 370170 439314 370226
rect 439370 370170 439438 370226
rect 439494 370170 439562 370226
rect 439618 370170 439686 370226
rect 439742 370170 470034 370226
rect 470090 370170 470158 370226
rect 470214 370170 470282 370226
rect 470338 370170 470406 370226
rect 470462 370170 500754 370226
rect 500810 370170 500878 370226
rect 500934 370170 501002 370226
rect 501058 370170 501126 370226
rect 501182 370170 531474 370226
rect 531530 370170 531598 370226
rect 531654 370170 531722 370226
rect 531778 370170 531846 370226
rect 531902 370170 562194 370226
rect 562250 370170 562318 370226
rect 562374 370170 562442 370226
rect 562498 370170 562566 370226
rect 562622 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect -1916 370102 597980 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 9234 370102
rect 9290 370046 9358 370102
rect 9414 370046 9482 370102
rect 9538 370046 9606 370102
rect 9662 370046 39954 370102
rect 40010 370046 40078 370102
rect 40134 370046 40202 370102
rect 40258 370046 40326 370102
rect 40382 370046 70674 370102
rect 70730 370046 70798 370102
rect 70854 370046 70922 370102
rect 70978 370046 71046 370102
rect 71102 370046 101394 370102
rect 101450 370046 101518 370102
rect 101574 370046 101642 370102
rect 101698 370046 101766 370102
rect 101822 370046 132114 370102
rect 132170 370046 132238 370102
rect 132294 370046 132362 370102
rect 132418 370046 132486 370102
rect 132542 370046 162834 370102
rect 162890 370046 162958 370102
rect 163014 370046 163082 370102
rect 163138 370046 163206 370102
rect 163262 370046 193554 370102
rect 193610 370046 193678 370102
rect 193734 370046 193802 370102
rect 193858 370046 193926 370102
rect 193982 370046 224274 370102
rect 224330 370046 224398 370102
rect 224454 370046 224522 370102
rect 224578 370046 224646 370102
rect 224702 370046 255878 370102
rect 255934 370046 256002 370102
rect 256058 370046 286598 370102
rect 286654 370046 286722 370102
rect 286778 370046 317318 370102
rect 317374 370046 317442 370102
rect 317498 370046 348038 370102
rect 348094 370046 348162 370102
rect 348218 370046 377874 370102
rect 377930 370046 377998 370102
rect 378054 370046 378122 370102
rect 378178 370046 378246 370102
rect 378302 370046 408594 370102
rect 408650 370046 408718 370102
rect 408774 370046 408842 370102
rect 408898 370046 408966 370102
rect 409022 370046 439314 370102
rect 439370 370046 439438 370102
rect 439494 370046 439562 370102
rect 439618 370046 439686 370102
rect 439742 370046 470034 370102
rect 470090 370046 470158 370102
rect 470214 370046 470282 370102
rect 470338 370046 470406 370102
rect 470462 370046 500754 370102
rect 500810 370046 500878 370102
rect 500934 370046 501002 370102
rect 501058 370046 501126 370102
rect 501182 370046 531474 370102
rect 531530 370046 531598 370102
rect 531654 370046 531722 370102
rect 531778 370046 531846 370102
rect 531902 370046 562194 370102
rect 562250 370046 562318 370102
rect 562374 370046 562442 370102
rect 562498 370046 562566 370102
rect 562622 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect -1916 369978 597980 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 9234 369978
rect 9290 369922 9358 369978
rect 9414 369922 9482 369978
rect 9538 369922 9606 369978
rect 9662 369922 39954 369978
rect 40010 369922 40078 369978
rect 40134 369922 40202 369978
rect 40258 369922 40326 369978
rect 40382 369922 70674 369978
rect 70730 369922 70798 369978
rect 70854 369922 70922 369978
rect 70978 369922 71046 369978
rect 71102 369922 101394 369978
rect 101450 369922 101518 369978
rect 101574 369922 101642 369978
rect 101698 369922 101766 369978
rect 101822 369922 132114 369978
rect 132170 369922 132238 369978
rect 132294 369922 132362 369978
rect 132418 369922 132486 369978
rect 132542 369922 162834 369978
rect 162890 369922 162958 369978
rect 163014 369922 163082 369978
rect 163138 369922 163206 369978
rect 163262 369922 193554 369978
rect 193610 369922 193678 369978
rect 193734 369922 193802 369978
rect 193858 369922 193926 369978
rect 193982 369922 224274 369978
rect 224330 369922 224398 369978
rect 224454 369922 224522 369978
rect 224578 369922 224646 369978
rect 224702 369922 255878 369978
rect 255934 369922 256002 369978
rect 256058 369922 286598 369978
rect 286654 369922 286722 369978
rect 286778 369922 317318 369978
rect 317374 369922 317442 369978
rect 317498 369922 348038 369978
rect 348094 369922 348162 369978
rect 348218 369922 377874 369978
rect 377930 369922 377998 369978
rect 378054 369922 378122 369978
rect 378178 369922 378246 369978
rect 378302 369922 408594 369978
rect 408650 369922 408718 369978
rect 408774 369922 408842 369978
rect 408898 369922 408966 369978
rect 409022 369922 439314 369978
rect 439370 369922 439438 369978
rect 439494 369922 439562 369978
rect 439618 369922 439686 369978
rect 439742 369922 470034 369978
rect 470090 369922 470158 369978
rect 470214 369922 470282 369978
rect 470338 369922 470406 369978
rect 470462 369922 500754 369978
rect 500810 369922 500878 369978
rect 500934 369922 501002 369978
rect 501058 369922 501126 369978
rect 501182 369922 531474 369978
rect 531530 369922 531598 369978
rect 531654 369922 531722 369978
rect 531778 369922 531846 369978
rect 531902 369922 562194 369978
rect 562250 369922 562318 369978
rect 562374 369922 562442 369978
rect 562498 369922 562566 369978
rect 562622 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect -1916 369826 597980 369922
rect -1916 364350 597980 364446
rect -1916 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 36234 364350
rect 36290 364294 36358 364350
rect 36414 364294 36482 364350
rect 36538 364294 36606 364350
rect 36662 364294 66954 364350
rect 67010 364294 67078 364350
rect 67134 364294 67202 364350
rect 67258 364294 67326 364350
rect 67382 364294 97674 364350
rect 97730 364294 97798 364350
rect 97854 364294 97922 364350
rect 97978 364294 98046 364350
rect 98102 364294 128394 364350
rect 128450 364294 128518 364350
rect 128574 364294 128642 364350
rect 128698 364294 128766 364350
rect 128822 364294 159114 364350
rect 159170 364294 159238 364350
rect 159294 364294 159362 364350
rect 159418 364294 159486 364350
rect 159542 364294 189834 364350
rect 189890 364294 189958 364350
rect 190014 364294 190082 364350
rect 190138 364294 190206 364350
rect 190262 364294 220554 364350
rect 220610 364294 220678 364350
rect 220734 364294 220802 364350
rect 220858 364294 220926 364350
rect 220982 364294 240518 364350
rect 240574 364294 240642 364350
rect 240698 364294 271238 364350
rect 271294 364294 271362 364350
rect 271418 364294 301958 364350
rect 302014 364294 302082 364350
rect 302138 364294 332678 364350
rect 332734 364294 332802 364350
rect 332858 364294 363398 364350
rect 363454 364294 363522 364350
rect 363578 364294 404874 364350
rect 404930 364294 404998 364350
rect 405054 364294 405122 364350
rect 405178 364294 405246 364350
rect 405302 364294 435594 364350
rect 435650 364294 435718 364350
rect 435774 364294 435842 364350
rect 435898 364294 435966 364350
rect 436022 364294 466314 364350
rect 466370 364294 466438 364350
rect 466494 364294 466562 364350
rect 466618 364294 466686 364350
rect 466742 364294 497034 364350
rect 497090 364294 497158 364350
rect 497214 364294 497282 364350
rect 497338 364294 497406 364350
rect 497462 364294 527754 364350
rect 527810 364294 527878 364350
rect 527934 364294 528002 364350
rect 528058 364294 528126 364350
rect 528182 364294 558474 364350
rect 558530 364294 558598 364350
rect 558654 364294 558722 364350
rect 558778 364294 558846 364350
rect 558902 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597980 364350
rect -1916 364226 597980 364294
rect -1916 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 36234 364226
rect 36290 364170 36358 364226
rect 36414 364170 36482 364226
rect 36538 364170 36606 364226
rect 36662 364170 66954 364226
rect 67010 364170 67078 364226
rect 67134 364170 67202 364226
rect 67258 364170 67326 364226
rect 67382 364170 97674 364226
rect 97730 364170 97798 364226
rect 97854 364170 97922 364226
rect 97978 364170 98046 364226
rect 98102 364170 128394 364226
rect 128450 364170 128518 364226
rect 128574 364170 128642 364226
rect 128698 364170 128766 364226
rect 128822 364170 159114 364226
rect 159170 364170 159238 364226
rect 159294 364170 159362 364226
rect 159418 364170 159486 364226
rect 159542 364170 189834 364226
rect 189890 364170 189958 364226
rect 190014 364170 190082 364226
rect 190138 364170 190206 364226
rect 190262 364170 220554 364226
rect 220610 364170 220678 364226
rect 220734 364170 220802 364226
rect 220858 364170 220926 364226
rect 220982 364170 240518 364226
rect 240574 364170 240642 364226
rect 240698 364170 271238 364226
rect 271294 364170 271362 364226
rect 271418 364170 301958 364226
rect 302014 364170 302082 364226
rect 302138 364170 332678 364226
rect 332734 364170 332802 364226
rect 332858 364170 363398 364226
rect 363454 364170 363522 364226
rect 363578 364170 404874 364226
rect 404930 364170 404998 364226
rect 405054 364170 405122 364226
rect 405178 364170 405246 364226
rect 405302 364170 435594 364226
rect 435650 364170 435718 364226
rect 435774 364170 435842 364226
rect 435898 364170 435966 364226
rect 436022 364170 466314 364226
rect 466370 364170 466438 364226
rect 466494 364170 466562 364226
rect 466618 364170 466686 364226
rect 466742 364170 497034 364226
rect 497090 364170 497158 364226
rect 497214 364170 497282 364226
rect 497338 364170 497406 364226
rect 497462 364170 527754 364226
rect 527810 364170 527878 364226
rect 527934 364170 528002 364226
rect 528058 364170 528126 364226
rect 528182 364170 558474 364226
rect 558530 364170 558598 364226
rect 558654 364170 558722 364226
rect 558778 364170 558846 364226
rect 558902 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597980 364226
rect -1916 364102 597980 364170
rect -1916 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 36234 364102
rect 36290 364046 36358 364102
rect 36414 364046 36482 364102
rect 36538 364046 36606 364102
rect 36662 364046 66954 364102
rect 67010 364046 67078 364102
rect 67134 364046 67202 364102
rect 67258 364046 67326 364102
rect 67382 364046 97674 364102
rect 97730 364046 97798 364102
rect 97854 364046 97922 364102
rect 97978 364046 98046 364102
rect 98102 364046 128394 364102
rect 128450 364046 128518 364102
rect 128574 364046 128642 364102
rect 128698 364046 128766 364102
rect 128822 364046 159114 364102
rect 159170 364046 159238 364102
rect 159294 364046 159362 364102
rect 159418 364046 159486 364102
rect 159542 364046 189834 364102
rect 189890 364046 189958 364102
rect 190014 364046 190082 364102
rect 190138 364046 190206 364102
rect 190262 364046 220554 364102
rect 220610 364046 220678 364102
rect 220734 364046 220802 364102
rect 220858 364046 220926 364102
rect 220982 364046 240518 364102
rect 240574 364046 240642 364102
rect 240698 364046 271238 364102
rect 271294 364046 271362 364102
rect 271418 364046 301958 364102
rect 302014 364046 302082 364102
rect 302138 364046 332678 364102
rect 332734 364046 332802 364102
rect 332858 364046 363398 364102
rect 363454 364046 363522 364102
rect 363578 364046 404874 364102
rect 404930 364046 404998 364102
rect 405054 364046 405122 364102
rect 405178 364046 405246 364102
rect 405302 364046 435594 364102
rect 435650 364046 435718 364102
rect 435774 364046 435842 364102
rect 435898 364046 435966 364102
rect 436022 364046 466314 364102
rect 466370 364046 466438 364102
rect 466494 364046 466562 364102
rect 466618 364046 466686 364102
rect 466742 364046 497034 364102
rect 497090 364046 497158 364102
rect 497214 364046 497282 364102
rect 497338 364046 497406 364102
rect 497462 364046 527754 364102
rect 527810 364046 527878 364102
rect 527934 364046 528002 364102
rect 528058 364046 528126 364102
rect 528182 364046 558474 364102
rect 558530 364046 558598 364102
rect 558654 364046 558722 364102
rect 558778 364046 558846 364102
rect 558902 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597980 364102
rect -1916 363978 597980 364046
rect -1916 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 36234 363978
rect 36290 363922 36358 363978
rect 36414 363922 36482 363978
rect 36538 363922 36606 363978
rect 36662 363922 66954 363978
rect 67010 363922 67078 363978
rect 67134 363922 67202 363978
rect 67258 363922 67326 363978
rect 67382 363922 97674 363978
rect 97730 363922 97798 363978
rect 97854 363922 97922 363978
rect 97978 363922 98046 363978
rect 98102 363922 128394 363978
rect 128450 363922 128518 363978
rect 128574 363922 128642 363978
rect 128698 363922 128766 363978
rect 128822 363922 159114 363978
rect 159170 363922 159238 363978
rect 159294 363922 159362 363978
rect 159418 363922 159486 363978
rect 159542 363922 189834 363978
rect 189890 363922 189958 363978
rect 190014 363922 190082 363978
rect 190138 363922 190206 363978
rect 190262 363922 220554 363978
rect 220610 363922 220678 363978
rect 220734 363922 220802 363978
rect 220858 363922 220926 363978
rect 220982 363922 240518 363978
rect 240574 363922 240642 363978
rect 240698 363922 271238 363978
rect 271294 363922 271362 363978
rect 271418 363922 301958 363978
rect 302014 363922 302082 363978
rect 302138 363922 332678 363978
rect 332734 363922 332802 363978
rect 332858 363922 363398 363978
rect 363454 363922 363522 363978
rect 363578 363922 404874 363978
rect 404930 363922 404998 363978
rect 405054 363922 405122 363978
rect 405178 363922 405246 363978
rect 405302 363922 435594 363978
rect 435650 363922 435718 363978
rect 435774 363922 435842 363978
rect 435898 363922 435966 363978
rect 436022 363922 466314 363978
rect 466370 363922 466438 363978
rect 466494 363922 466562 363978
rect 466618 363922 466686 363978
rect 466742 363922 497034 363978
rect 497090 363922 497158 363978
rect 497214 363922 497282 363978
rect 497338 363922 497406 363978
rect 497462 363922 527754 363978
rect 527810 363922 527878 363978
rect 527934 363922 528002 363978
rect 528058 363922 528126 363978
rect 528182 363922 558474 363978
rect 558530 363922 558598 363978
rect 558654 363922 558722 363978
rect 558778 363922 558846 363978
rect 558902 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597980 363978
rect -1916 363826 597980 363922
rect -1916 352350 597980 352446
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 9234 352350
rect 9290 352294 9358 352350
rect 9414 352294 9482 352350
rect 9538 352294 9606 352350
rect 9662 352294 39954 352350
rect 40010 352294 40078 352350
rect 40134 352294 40202 352350
rect 40258 352294 40326 352350
rect 40382 352294 70674 352350
rect 70730 352294 70798 352350
rect 70854 352294 70922 352350
rect 70978 352294 71046 352350
rect 71102 352294 101394 352350
rect 101450 352294 101518 352350
rect 101574 352294 101642 352350
rect 101698 352294 101766 352350
rect 101822 352294 132114 352350
rect 132170 352294 132238 352350
rect 132294 352294 132362 352350
rect 132418 352294 132486 352350
rect 132542 352294 162834 352350
rect 162890 352294 162958 352350
rect 163014 352294 163082 352350
rect 163138 352294 163206 352350
rect 163262 352294 169878 352350
rect 169934 352294 170002 352350
rect 170058 352294 193554 352350
rect 193610 352294 193678 352350
rect 193734 352294 193802 352350
rect 193858 352294 193926 352350
rect 193982 352294 224274 352350
rect 224330 352294 224398 352350
rect 224454 352294 224522 352350
rect 224578 352294 224646 352350
rect 224702 352294 255878 352350
rect 255934 352294 256002 352350
rect 256058 352294 286598 352350
rect 286654 352294 286722 352350
rect 286778 352294 317318 352350
rect 317374 352294 317442 352350
rect 317498 352294 348038 352350
rect 348094 352294 348162 352350
rect 348218 352294 377874 352350
rect 377930 352294 377998 352350
rect 378054 352294 378122 352350
rect 378178 352294 378246 352350
rect 378302 352294 408594 352350
rect 408650 352294 408718 352350
rect 408774 352294 408842 352350
rect 408898 352294 408966 352350
rect 409022 352294 439314 352350
rect 439370 352294 439438 352350
rect 439494 352294 439562 352350
rect 439618 352294 439686 352350
rect 439742 352294 470034 352350
rect 470090 352294 470158 352350
rect 470214 352294 470282 352350
rect 470338 352294 470406 352350
rect 470462 352294 500754 352350
rect 500810 352294 500878 352350
rect 500934 352294 501002 352350
rect 501058 352294 501126 352350
rect 501182 352294 531474 352350
rect 531530 352294 531598 352350
rect 531654 352294 531722 352350
rect 531778 352294 531846 352350
rect 531902 352294 562194 352350
rect 562250 352294 562318 352350
rect 562374 352294 562442 352350
rect 562498 352294 562566 352350
rect 562622 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect -1916 352226 597980 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 9234 352226
rect 9290 352170 9358 352226
rect 9414 352170 9482 352226
rect 9538 352170 9606 352226
rect 9662 352170 39954 352226
rect 40010 352170 40078 352226
rect 40134 352170 40202 352226
rect 40258 352170 40326 352226
rect 40382 352170 70674 352226
rect 70730 352170 70798 352226
rect 70854 352170 70922 352226
rect 70978 352170 71046 352226
rect 71102 352170 101394 352226
rect 101450 352170 101518 352226
rect 101574 352170 101642 352226
rect 101698 352170 101766 352226
rect 101822 352170 132114 352226
rect 132170 352170 132238 352226
rect 132294 352170 132362 352226
rect 132418 352170 132486 352226
rect 132542 352170 162834 352226
rect 162890 352170 162958 352226
rect 163014 352170 163082 352226
rect 163138 352170 163206 352226
rect 163262 352170 169878 352226
rect 169934 352170 170002 352226
rect 170058 352170 193554 352226
rect 193610 352170 193678 352226
rect 193734 352170 193802 352226
rect 193858 352170 193926 352226
rect 193982 352170 224274 352226
rect 224330 352170 224398 352226
rect 224454 352170 224522 352226
rect 224578 352170 224646 352226
rect 224702 352170 255878 352226
rect 255934 352170 256002 352226
rect 256058 352170 286598 352226
rect 286654 352170 286722 352226
rect 286778 352170 317318 352226
rect 317374 352170 317442 352226
rect 317498 352170 348038 352226
rect 348094 352170 348162 352226
rect 348218 352170 377874 352226
rect 377930 352170 377998 352226
rect 378054 352170 378122 352226
rect 378178 352170 378246 352226
rect 378302 352170 408594 352226
rect 408650 352170 408718 352226
rect 408774 352170 408842 352226
rect 408898 352170 408966 352226
rect 409022 352170 439314 352226
rect 439370 352170 439438 352226
rect 439494 352170 439562 352226
rect 439618 352170 439686 352226
rect 439742 352170 470034 352226
rect 470090 352170 470158 352226
rect 470214 352170 470282 352226
rect 470338 352170 470406 352226
rect 470462 352170 500754 352226
rect 500810 352170 500878 352226
rect 500934 352170 501002 352226
rect 501058 352170 501126 352226
rect 501182 352170 531474 352226
rect 531530 352170 531598 352226
rect 531654 352170 531722 352226
rect 531778 352170 531846 352226
rect 531902 352170 562194 352226
rect 562250 352170 562318 352226
rect 562374 352170 562442 352226
rect 562498 352170 562566 352226
rect 562622 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect -1916 352102 597980 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 9234 352102
rect 9290 352046 9358 352102
rect 9414 352046 9482 352102
rect 9538 352046 9606 352102
rect 9662 352046 39954 352102
rect 40010 352046 40078 352102
rect 40134 352046 40202 352102
rect 40258 352046 40326 352102
rect 40382 352046 70674 352102
rect 70730 352046 70798 352102
rect 70854 352046 70922 352102
rect 70978 352046 71046 352102
rect 71102 352046 101394 352102
rect 101450 352046 101518 352102
rect 101574 352046 101642 352102
rect 101698 352046 101766 352102
rect 101822 352046 132114 352102
rect 132170 352046 132238 352102
rect 132294 352046 132362 352102
rect 132418 352046 132486 352102
rect 132542 352046 162834 352102
rect 162890 352046 162958 352102
rect 163014 352046 163082 352102
rect 163138 352046 163206 352102
rect 163262 352046 169878 352102
rect 169934 352046 170002 352102
rect 170058 352046 193554 352102
rect 193610 352046 193678 352102
rect 193734 352046 193802 352102
rect 193858 352046 193926 352102
rect 193982 352046 224274 352102
rect 224330 352046 224398 352102
rect 224454 352046 224522 352102
rect 224578 352046 224646 352102
rect 224702 352046 255878 352102
rect 255934 352046 256002 352102
rect 256058 352046 286598 352102
rect 286654 352046 286722 352102
rect 286778 352046 317318 352102
rect 317374 352046 317442 352102
rect 317498 352046 348038 352102
rect 348094 352046 348162 352102
rect 348218 352046 377874 352102
rect 377930 352046 377998 352102
rect 378054 352046 378122 352102
rect 378178 352046 378246 352102
rect 378302 352046 408594 352102
rect 408650 352046 408718 352102
rect 408774 352046 408842 352102
rect 408898 352046 408966 352102
rect 409022 352046 439314 352102
rect 439370 352046 439438 352102
rect 439494 352046 439562 352102
rect 439618 352046 439686 352102
rect 439742 352046 470034 352102
rect 470090 352046 470158 352102
rect 470214 352046 470282 352102
rect 470338 352046 470406 352102
rect 470462 352046 500754 352102
rect 500810 352046 500878 352102
rect 500934 352046 501002 352102
rect 501058 352046 501126 352102
rect 501182 352046 531474 352102
rect 531530 352046 531598 352102
rect 531654 352046 531722 352102
rect 531778 352046 531846 352102
rect 531902 352046 562194 352102
rect 562250 352046 562318 352102
rect 562374 352046 562442 352102
rect 562498 352046 562566 352102
rect 562622 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect -1916 351978 597980 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 9234 351978
rect 9290 351922 9358 351978
rect 9414 351922 9482 351978
rect 9538 351922 9606 351978
rect 9662 351922 39954 351978
rect 40010 351922 40078 351978
rect 40134 351922 40202 351978
rect 40258 351922 40326 351978
rect 40382 351922 70674 351978
rect 70730 351922 70798 351978
rect 70854 351922 70922 351978
rect 70978 351922 71046 351978
rect 71102 351922 101394 351978
rect 101450 351922 101518 351978
rect 101574 351922 101642 351978
rect 101698 351922 101766 351978
rect 101822 351922 132114 351978
rect 132170 351922 132238 351978
rect 132294 351922 132362 351978
rect 132418 351922 132486 351978
rect 132542 351922 162834 351978
rect 162890 351922 162958 351978
rect 163014 351922 163082 351978
rect 163138 351922 163206 351978
rect 163262 351922 169878 351978
rect 169934 351922 170002 351978
rect 170058 351922 193554 351978
rect 193610 351922 193678 351978
rect 193734 351922 193802 351978
rect 193858 351922 193926 351978
rect 193982 351922 224274 351978
rect 224330 351922 224398 351978
rect 224454 351922 224522 351978
rect 224578 351922 224646 351978
rect 224702 351922 255878 351978
rect 255934 351922 256002 351978
rect 256058 351922 286598 351978
rect 286654 351922 286722 351978
rect 286778 351922 317318 351978
rect 317374 351922 317442 351978
rect 317498 351922 348038 351978
rect 348094 351922 348162 351978
rect 348218 351922 377874 351978
rect 377930 351922 377998 351978
rect 378054 351922 378122 351978
rect 378178 351922 378246 351978
rect 378302 351922 408594 351978
rect 408650 351922 408718 351978
rect 408774 351922 408842 351978
rect 408898 351922 408966 351978
rect 409022 351922 439314 351978
rect 439370 351922 439438 351978
rect 439494 351922 439562 351978
rect 439618 351922 439686 351978
rect 439742 351922 470034 351978
rect 470090 351922 470158 351978
rect 470214 351922 470282 351978
rect 470338 351922 470406 351978
rect 470462 351922 500754 351978
rect 500810 351922 500878 351978
rect 500934 351922 501002 351978
rect 501058 351922 501126 351978
rect 501182 351922 531474 351978
rect 531530 351922 531598 351978
rect 531654 351922 531722 351978
rect 531778 351922 531846 351978
rect 531902 351922 562194 351978
rect 562250 351922 562318 351978
rect 562374 351922 562442 351978
rect 562498 351922 562566 351978
rect 562622 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect -1916 351826 597980 351922
rect -1916 346350 597980 346446
rect -1916 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 36234 346350
rect 36290 346294 36358 346350
rect 36414 346294 36482 346350
rect 36538 346294 36606 346350
rect 36662 346294 66954 346350
rect 67010 346294 67078 346350
rect 67134 346294 67202 346350
rect 67258 346294 67326 346350
rect 67382 346294 97674 346350
rect 97730 346294 97798 346350
rect 97854 346294 97922 346350
rect 97978 346294 98046 346350
rect 98102 346294 128394 346350
rect 128450 346294 128518 346350
rect 128574 346294 128642 346350
rect 128698 346294 128766 346350
rect 128822 346294 154518 346350
rect 154574 346294 154642 346350
rect 154698 346294 159114 346350
rect 159170 346294 159238 346350
rect 159294 346294 159362 346350
rect 159418 346294 159486 346350
rect 159542 346294 185238 346350
rect 185294 346294 185362 346350
rect 185418 346294 189834 346350
rect 189890 346294 189958 346350
rect 190014 346294 190082 346350
rect 190138 346294 190206 346350
rect 190262 346294 220554 346350
rect 220610 346294 220678 346350
rect 220734 346294 220802 346350
rect 220858 346294 220926 346350
rect 220982 346294 240518 346350
rect 240574 346294 240642 346350
rect 240698 346294 271238 346350
rect 271294 346294 271362 346350
rect 271418 346294 301958 346350
rect 302014 346294 302082 346350
rect 302138 346294 332678 346350
rect 332734 346294 332802 346350
rect 332858 346294 363398 346350
rect 363454 346294 363522 346350
rect 363578 346294 404874 346350
rect 404930 346294 404998 346350
rect 405054 346294 405122 346350
rect 405178 346294 405246 346350
rect 405302 346294 435594 346350
rect 435650 346294 435718 346350
rect 435774 346294 435842 346350
rect 435898 346294 435966 346350
rect 436022 346294 466314 346350
rect 466370 346294 466438 346350
rect 466494 346294 466562 346350
rect 466618 346294 466686 346350
rect 466742 346294 497034 346350
rect 497090 346294 497158 346350
rect 497214 346294 497282 346350
rect 497338 346294 497406 346350
rect 497462 346294 527754 346350
rect 527810 346294 527878 346350
rect 527934 346294 528002 346350
rect 528058 346294 528126 346350
rect 528182 346294 558474 346350
rect 558530 346294 558598 346350
rect 558654 346294 558722 346350
rect 558778 346294 558846 346350
rect 558902 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597980 346350
rect -1916 346226 597980 346294
rect -1916 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 36234 346226
rect 36290 346170 36358 346226
rect 36414 346170 36482 346226
rect 36538 346170 36606 346226
rect 36662 346170 66954 346226
rect 67010 346170 67078 346226
rect 67134 346170 67202 346226
rect 67258 346170 67326 346226
rect 67382 346170 97674 346226
rect 97730 346170 97798 346226
rect 97854 346170 97922 346226
rect 97978 346170 98046 346226
rect 98102 346170 128394 346226
rect 128450 346170 128518 346226
rect 128574 346170 128642 346226
rect 128698 346170 128766 346226
rect 128822 346170 154518 346226
rect 154574 346170 154642 346226
rect 154698 346170 159114 346226
rect 159170 346170 159238 346226
rect 159294 346170 159362 346226
rect 159418 346170 159486 346226
rect 159542 346170 185238 346226
rect 185294 346170 185362 346226
rect 185418 346170 189834 346226
rect 189890 346170 189958 346226
rect 190014 346170 190082 346226
rect 190138 346170 190206 346226
rect 190262 346170 220554 346226
rect 220610 346170 220678 346226
rect 220734 346170 220802 346226
rect 220858 346170 220926 346226
rect 220982 346170 240518 346226
rect 240574 346170 240642 346226
rect 240698 346170 271238 346226
rect 271294 346170 271362 346226
rect 271418 346170 301958 346226
rect 302014 346170 302082 346226
rect 302138 346170 332678 346226
rect 332734 346170 332802 346226
rect 332858 346170 363398 346226
rect 363454 346170 363522 346226
rect 363578 346170 404874 346226
rect 404930 346170 404998 346226
rect 405054 346170 405122 346226
rect 405178 346170 405246 346226
rect 405302 346170 435594 346226
rect 435650 346170 435718 346226
rect 435774 346170 435842 346226
rect 435898 346170 435966 346226
rect 436022 346170 466314 346226
rect 466370 346170 466438 346226
rect 466494 346170 466562 346226
rect 466618 346170 466686 346226
rect 466742 346170 497034 346226
rect 497090 346170 497158 346226
rect 497214 346170 497282 346226
rect 497338 346170 497406 346226
rect 497462 346170 527754 346226
rect 527810 346170 527878 346226
rect 527934 346170 528002 346226
rect 528058 346170 528126 346226
rect 528182 346170 558474 346226
rect 558530 346170 558598 346226
rect 558654 346170 558722 346226
rect 558778 346170 558846 346226
rect 558902 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597980 346226
rect -1916 346102 597980 346170
rect -1916 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 36234 346102
rect 36290 346046 36358 346102
rect 36414 346046 36482 346102
rect 36538 346046 36606 346102
rect 36662 346046 66954 346102
rect 67010 346046 67078 346102
rect 67134 346046 67202 346102
rect 67258 346046 67326 346102
rect 67382 346046 97674 346102
rect 97730 346046 97798 346102
rect 97854 346046 97922 346102
rect 97978 346046 98046 346102
rect 98102 346046 128394 346102
rect 128450 346046 128518 346102
rect 128574 346046 128642 346102
rect 128698 346046 128766 346102
rect 128822 346046 154518 346102
rect 154574 346046 154642 346102
rect 154698 346046 159114 346102
rect 159170 346046 159238 346102
rect 159294 346046 159362 346102
rect 159418 346046 159486 346102
rect 159542 346046 185238 346102
rect 185294 346046 185362 346102
rect 185418 346046 189834 346102
rect 189890 346046 189958 346102
rect 190014 346046 190082 346102
rect 190138 346046 190206 346102
rect 190262 346046 220554 346102
rect 220610 346046 220678 346102
rect 220734 346046 220802 346102
rect 220858 346046 220926 346102
rect 220982 346046 240518 346102
rect 240574 346046 240642 346102
rect 240698 346046 271238 346102
rect 271294 346046 271362 346102
rect 271418 346046 301958 346102
rect 302014 346046 302082 346102
rect 302138 346046 332678 346102
rect 332734 346046 332802 346102
rect 332858 346046 363398 346102
rect 363454 346046 363522 346102
rect 363578 346046 404874 346102
rect 404930 346046 404998 346102
rect 405054 346046 405122 346102
rect 405178 346046 405246 346102
rect 405302 346046 435594 346102
rect 435650 346046 435718 346102
rect 435774 346046 435842 346102
rect 435898 346046 435966 346102
rect 436022 346046 466314 346102
rect 466370 346046 466438 346102
rect 466494 346046 466562 346102
rect 466618 346046 466686 346102
rect 466742 346046 497034 346102
rect 497090 346046 497158 346102
rect 497214 346046 497282 346102
rect 497338 346046 497406 346102
rect 497462 346046 527754 346102
rect 527810 346046 527878 346102
rect 527934 346046 528002 346102
rect 528058 346046 528126 346102
rect 528182 346046 558474 346102
rect 558530 346046 558598 346102
rect 558654 346046 558722 346102
rect 558778 346046 558846 346102
rect 558902 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597980 346102
rect -1916 345978 597980 346046
rect -1916 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 36234 345978
rect 36290 345922 36358 345978
rect 36414 345922 36482 345978
rect 36538 345922 36606 345978
rect 36662 345922 66954 345978
rect 67010 345922 67078 345978
rect 67134 345922 67202 345978
rect 67258 345922 67326 345978
rect 67382 345922 97674 345978
rect 97730 345922 97798 345978
rect 97854 345922 97922 345978
rect 97978 345922 98046 345978
rect 98102 345922 128394 345978
rect 128450 345922 128518 345978
rect 128574 345922 128642 345978
rect 128698 345922 128766 345978
rect 128822 345922 154518 345978
rect 154574 345922 154642 345978
rect 154698 345922 159114 345978
rect 159170 345922 159238 345978
rect 159294 345922 159362 345978
rect 159418 345922 159486 345978
rect 159542 345922 185238 345978
rect 185294 345922 185362 345978
rect 185418 345922 189834 345978
rect 189890 345922 189958 345978
rect 190014 345922 190082 345978
rect 190138 345922 190206 345978
rect 190262 345922 220554 345978
rect 220610 345922 220678 345978
rect 220734 345922 220802 345978
rect 220858 345922 220926 345978
rect 220982 345922 240518 345978
rect 240574 345922 240642 345978
rect 240698 345922 271238 345978
rect 271294 345922 271362 345978
rect 271418 345922 301958 345978
rect 302014 345922 302082 345978
rect 302138 345922 332678 345978
rect 332734 345922 332802 345978
rect 332858 345922 363398 345978
rect 363454 345922 363522 345978
rect 363578 345922 404874 345978
rect 404930 345922 404998 345978
rect 405054 345922 405122 345978
rect 405178 345922 405246 345978
rect 405302 345922 435594 345978
rect 435650 345922 435718 345978
rect 435774 345922 435842 345978
rect 435898 345922 435966 345978
rect 436022 345922 466314 345978
rect 466370 345922 466438 345978
rect 466494 345922 466562 345978
rect 466618 345922 466686 345978
rect 466742 345922 497034 345978
rect 497090 345922 497158 345978
rect 497214 345922 497282 345978
rect 497338 345922 497406 345978
rect 497462 345922 527754 345978
rect 527810 345922 527878 345978
rect 527934 345922 528002 345978
rect 528058 345922 528126 345978
rect 528182 345922 558474 345978
rect 558530 345922 558598 345978
rect 558654 345922 558722 345978
rect 558778 345922 558846 345978
rect 558902 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597980 345978
rect -1916 345826 597980 345922
rect -1916 334350 597980 334446
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 9234 334350
rect 9290 334294 9358 334350
rect 9414 334294 9482 334350
rect 9538 334294 9606 334350
rect 9662 334294 39954 334350
rect 40010 334294 40078 334350
rect 40134 334294 40202 334350
rect 40258 334294 40326 334350
rect 40382 334294 70674 334350
rect 70730 334294 70798 334350
rect 70854 334294 70922 334350
rect 70978 334294 71046 334350
rect 71102 334294 101394 334350
rect 101450 334294 101518 334350
rect 101574 334294 101642 334350
rect 101698 334294 101766 334350
rect 101822 334294 132114 334350
rect 132170 334294 132238 334350
rect 132294 334294 132362 334350
rect 132418 334294 132486 334350
rect 132542 334294 162834 334350
rect 162890 334294 162958 334350
rect 163014 334294 163082 334350
rect 163138 334294 163206 334350
rect 163262 334294 169878 334350
rect 169934 334294 170002 334350
rect 170058 334294 193554 334350
rect 193610 334294 193678 334350
rect 193734 334294 193802 334350
rect 193858 334294 193926 334350
rect 193982 334294 224274 334350
rect 224330 334294 224398 334350
rect 224454 334294 224522 334350
rect 224578 334294 224646 334350
rect 224702 334294 255878 334350
rect 255934 334294 256002 334350
rect 256058 334294 286598 334350
rect 286654 334294 286722 334350
rect 286778 334294 317318 334350
rect 317374 334294 317442 334350
rect 317498 334294 348038 334350
rect 348094 334294 348162 334350
rect 348218 334294 377874 334350
rect 377930 334294 377998 334350
rect 378054 334294 378122 334350
rect 378178 334294 378246 334350
rect 378302 334294 408594 334350
rect 408650 334294 408718 334350
rect 408774 334294 408842 334350
rect 408898 334294 408966 334350
rect 409022 334294 439314 334350
rect 439370 334294 439438 334350
rect 439494 334294 439562 334350
rect 439618 334294 439686 334350
rect 439742 334294 470034 334350
rect 470090 334294 470158 334350
rect 470214 334294 470282 334350
rect 470338 334294 470406 334350
rect 470462 334294 500754 334350
rect 500810 334294 500878 334350
rect 500934 334294 501002 334350
rect 501058 334294 501126 334350
rect 501182 334294 531474 334350
rect 531530 334294 531598 334350
rect 531654 334294 531722 334350
rect 531778 334294 531846 334350
rect 531902 334294 562194 334350
rect 562250 334294 562318 334350
rect 562374 334294 562442 334350
rect 562498 334294 562566 334350
rect 562622 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect -1916 334226 597980 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 9234 334226
rect 9290 334170 9358 334226
rect 9414 334170 9482 334226
rect 9538 334170 9606 334226
rect 9662 334170 39954 334226
rect 40010 334170 40078 334226
rect 40134 334170 40202 334226
rect 40258 334170 40326 334226
rect 40382 334170 70674 334226
rect 70730 334170 70798 334226
rect 70854 334170 70922 334226
rect 70978 334170 71046 334226
rect 71102 334170 101394 334226
rect 101450 334170 101518 334226
rect 101574 334170 101642 334226
rect 101698 334170 101766 334226
rect 101822 334170 132114 334226
rect 132170 334170 132238 334226
rect 132294 334170 132362 334226
rect 132418 334170 132486 334226
rect 132542 334170 162834 334226
rect 162890 334170 162958 334226
rect 163014 334170 163082 334226
rect 163138 334170 163206 334226
rect 163262 334170 169878 334226
rect 169934 334170 170002 334226
rect 170058 334170 193554 334226
rect 193610 334170 193678 334226
rect 193734 334170 193802 334226
rect 193858 334170 193926 334226
rect 193982 334170 224274 334226
rect 224330 334170 224398 334226
rect 224454 334170 224522 334226
rect 224578 334170 224646 334226
rect 224702 334170 255878 334226
rect 255934 334170 256002 334226
rect 256058 334170 286598 334226
rect 286654 334170 286722 334226
rect 286778 334170 317318 334226
rect 317374 334170 317442 334226
rect 317498 334170 348038 334226
rect 348094 334170 348162 334226
rect 348218 334170 377874 334226
rect 377930 334170 377998 334226
rect 378054 334170 378122 334226
rect 378178 334170 378246 334226
rect 378302 334170 408594 334226
rect 408650 334170 408718 334226
rect 408774 334170 408842 334226
rect 408898 334170 408966 334226
rect 409022 334170 439314 334226
rect 439370 334170 439438 334226
rect 439494 334170 439562 334226
rect 439618 334170 439686 334226
rect 439742 334170 470034 334226
rect 470090 334170 470158 334226
rect 470214 334170 470282 334226
rect 470338 334170 470406 334226
rect 470462 334170 500754 334226
rect 500810 334170 500878 334226
rect 500934 334170 501002 334226
rect 501058 334170 501126 334226
rect 501182 334170 531474 334226
rect 531530 334170 531598 334226
rect 531654 334170 531722 334226
rect 531778 334170 531846 334226
rect 531902 334170 562194 334226
rect 562250 334170 562318 334226
rect 562374 334170 562442 334226
rect 562498 334170 562566 334226
rect 562622 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect -1916 334102 597980 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 9234 334102
rect 9290 334046 9358 334102
rect 9414 334046 9482 334102
rect 9538 334046 9606 334102
rect 9662 334046 39954 334102
rect 40010 334046 40078 334102
rect 40134 334046 40202 334102
rect 40258 334046 40326 334102
rect 40382 334046 70674 334102
rect 70730 334046 70798 334102
rect 70854 334046 70922 334102
rect 70978 334046 71046 334102
rect 71102 334046 101394 334102
rect 101450 334046 101518 334102
rect 101574 334046 101642 334102
rect 101698 334046 101766 334102
rect 101822 334046 132114 334102
rect 132170 334046 132238 334102
rect 132294 334046 132362 334102
rect 132418 334046 132486 334102
rect 132542 334046 162834 334102
rect 162890 334046 162958 334102
rect 163014 334046 163082 334102
rect 163138 334046 163206 334102
rect 163262 334046 169878 334102
rect 169934 334046 170002 334102
rect 170058 334046 193554 334102
rect 193610 334046 193678 334102
rect 193734 334046 193802 334102
rect 193858 334046 193926 334102
rect 193982 334046 224274 334102
rect 224330 334046 224398 334102
rect 224454 334046 224522 334102
rect 224578 334046 224646 334102
rect 224702 334046 255878 334102
rect 255934 334046 256002 334102
rect 256058 334046 286598 334102
rect 286654 334046 286722 334102
rect 286778 334046 317318 334102
rect 317374 334046 317442 334102
rect 317498 334046 348038 334102
rect 348094 334046 348162 334102
rect 348218 334046 377874 334102
rect 377930 334046 377998 334102
rect 378054 334046 378122 334102
rect 378178 334046 378246 334102
rect 378302 334046 408594 334102
rect 408650 334046 408718 334102
rect 408774 334046 408842 334102
rect 408898 334046 408966 334102
rect 409022 334046 439314 334102
rect 439370 334046 439438 334102
rect 439494 334046 439562 334102
rect 439618 334046 439686 334102
rect 439742 334046 470034 334102
rect 470090 334046 470158 334102
rect 470214 334046 470282 334102
rect 470338 334046 470406 334102
rect 470462 334046 500754 334102
rect 500810 334046 500878 334102
rect 500934 334046 501002 334102
rect 501058 334046 501126 334102
rect 501182 334046 531474 334102
rect 531530 334046 531598 334102
rect 531654 334046 531722 334102
rect 531778 334046 531846 334102
rect 531902 334046 562194 334102
rect 562250 334046 562318 334102
rect 562374 334046 562442 334102
rect 562498 334046 562566 334102
rect 562622 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect -1916 333978 597980 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 9234 333978
rect 9290 333922 9358 333978
rect 9414 333922 9482 333978
rect 9538 333922 9606 333978
rect 9662 333922 39954 333978
rect 40010 333922 40078 333978
rect 40134 333922 40202 333978
rect 40258 333922 40326 333978
rect 40382 333922 70674 333978
rect 70730 333922 70798 333978
rect 70854 333922 70922 333978
rect 70978 333922 71046 333978
rect 71102 333922 101394 333978
rect 101450 333922 101518 333978
rect 101574 333922 101642 333978
rect 101698 333922 101766 333978
rect 101822 333922 132114 333978
rect 132170 333922 132238 333978
rect 132294 333922 132362 333978
rect 132418 333922 132486 333978
rect 132542 333922 162834 333978
rect 162890 333922 162958 333978
rect 163014 333922 163082 333978
rect 163138 333922 163206 333978
rect 163262 333922 169878 333978
rect 169934 333922 170002 333978
rect 170058 333922 193554 333978
rect 193610 333922 193678 333978
rect 193734 333922 193802 333978
rect 193858 333922 193926 333978
rect 193982 333922 224274 333978
rect 224330 333922 224398 333978
rect 224454 333922 224522 333978
rect 224578 333922 224646 333978
rect 224702 333922 255878 333978
rect 255934 333922 256002 333978
rect 256058 333922 286598 333978
rect 286654 333922 286722 333978
rect 286778 333922 317318 333978
rect 317374 333922 317442 333978
rect 317498 333922 348038 333978
rect 348094 333922 348162 333978
rect 348218 333922 377874 333978
rect 377930 333922 377998 333978
rect 378054 333922 378122 333978
rect 378178 333922 378246 333978
rect 378302 333922 408594 333978
rect 408650 333922 408718 333978
rect 408774 333922 408842 333978
rect 408898 333922 408966 333978
rect 409022 333922 439314 333978
rect 439370 333922 439438 333978
rect 439494 333922 439562 333978
rect 439618 333922 439686 333978
rect 439742 333922 470034 333978
rect 470090 333922 470158 333978
rect 470214 333922 470282 333978
rect 470338 333922 470406 333978
rect 470462 333922 500754 333978
rect 500810 333922 500878 333978
rect 500934 333922 501002 333978
rect 501058 333922 501126 333978
rect 501182 333922 531474 333978
rect 531530 333922 531598 333978
rect 531654 333922 531722 333978
rect 531778 333922 531846 333978
rect 531902 333922 562194 333978
rect 562250 333922 562318 333978
rect 562374 333922 562442 333978
rect 562498 333922 562566 333978
rect 562622 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect -1916 333826 597980 333922
rect -1916 328350 597980 328446
rect -1916 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 36234 328350
rect 36290 328294 36358 328350
rect 36414 328294 36482 328350
rect 36538 328294 36606 328350
rect 36662 328294 66954 328350
rect 67010 328294 67078 328350
rect 67134 328294 67202 328350
rect 67258 328294 67326 328350
rect 67382 328294 97674 328350
rect 97730 328294 97798 328350
rect 97854 328294 97922 328350
rect 97978 328294 98046 328350
rect 98102 328294 128394 328350
rect 128450 328294 128518 328350
rect 128574 328294 128642 328350
rect 128698 328294 128766 328350
rect 128822 328294 154518 328350
rect 154574 328294 154642 328350
rect 154698 328294 159114 328350
rect 159170 328294 159238 328350
rect 159294 328294 159362 328350
rect 159418 328294 159486 328350
rect 159542 328294 185238 328350
rect 185294 328294 185362 328350
rect 185418 328294 189834 328350
rect 189890 328294 189958 328350
rect 190014 328294 190082 328350
rect 190138 328294 190206 328350
rect 190262 328294 220554 328350
rect 220610 328294 220678 328350
rect 220734 328294 220802 328350
rect 220858 328294 220926 328350
rect 220982 328294 240518 328350
rect 240574 328294 240642 328350
rect 240698 328294 271238 328350
rect 271294 328294 271362 328350
rect 271418 328294 301958 328350
rect 302014 328294 302082 328350
rect 302138 328294 332678 328350
rect 332734 328294 332802 328350
rect 332858 328294 363398 328350
rect 363454 328294 363522 328350
rect 363578 328294 404874 328350
rect 404930 328294 404998 328350
rect 405054 328294 405122 328350
rect 405178 328294 405246 328350
rect 405302 328294 435594 328350
rect 435650 328294 435718 328350
rect 435774 328294 435842 328350
rect 435898 328294 435966 328350
rect 436022 328294 466314 328350
rect 466370 328294 466438 328350
rect 466494 328294 466562 328350
rect 466618 328294 466686 328350
rect 466742 328294 497034 328350
rect 497090 328294 497158 328350
rect 497214 328294 497282 328350
rect 497338 328294 497406 328350
rect 497462 328294 527754 328350
rect 527810 328294 527878 328350
rect 527934 328294 528002 328350
rect 528058 328294 528126 328350
rect 528182 328294 558474 328350
rect 558530 328294 558598 328350
rect 558654 328294 558722 328350
rect 558778 328294 558846 328350
rect 558902 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597980 328350
rect -1916 328226 597980 328294
rect -1916 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 36234 328226
rect 36290 328170 36358 328226
rect 36414 328170 36482 328226
rect 36538 328170 36606 328226
rect 36662 328170 66954 328226
rect 67010 328170 67078 328226
rect 67134 328170 67202 328226
rect 67258 328170 67326 328226
rect 67382 328170 97674 328226
rect 97730 328170 97798 328226
rect 97854 328170 97922 328226
rect 97978 328170 98046 328226
rect 98102 328170 128394 328226
rect 128450 328170 128518 328226
rect 128574 328170 128642 328226
rect 128698 328170 128766 328226
rect 128822 328170 154518 328226
rect 154574 328170 154642 328226
rect 154698 328170 159114 328226
rect 159170 328170 159238 328226
rect 159294 328170 159362 328226
rect 159418 328170 159486 328226
rect 159542 328170 185238 328226
rect 185294 328170 185362 328226
rect 185418 328170 189834 328226
rect 189890 328170 189958 328226
rect 190014 328170 190082 328226
rect 190138 328170 190206 328226
rect 190262 328170 220554 328226
rect 220610 328170 220678 328226
rect 220734 328170 220802 328226
rect 220858 328170 220926 328226
rect 220982 328170 240518 328226
rect 240574 328170 240642 328226
rect 240698 328170 271238 328226
rect 271294 328170 271362 328226
rect 271418 328170 301958 328226
rect 302014 328170 302082 328226
rect 302138 328170 332678 328226
rect 332734 328170 332802 328226
rect 332858 328170 363398 328226
rect 363454 328170 363522 328226
rect 363578 328170 404874 328226
rect 404930 328170 404998 328226
rect 405054 328170 405122 328226
rect 405178 328170 405246 328226
rect 405302 328170 435594 328226
rect 435650 328170 435718 328226
rect 435774 328170 435842 328226
rect 435898 328170 435966 328226
rect 436022 328170 466314 328226
rect 466370 328170 466438 328226
rect 466494 328170 466562 328226
rect 466618 328170 466686 328226
rect 466742 328170 497034 328226
rect 497090 328170 497158 328226
rect 497214 328170 497282 328226
rect 497338 328170 497406 328226
rect 497462 328170 527754 328226
rect 527810 328170 527878 328226
rect 527934 328170 528002 328226
rect 528058 328170 528126 328226
rect 528182 328170 558474 328226
rect 558530 328170 558598 328226
rect 558654 328170 558722 328226
rect 558778 328170 558846 328226
rect 558902 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597980 328226
rect -1916 328102 597980 328170
rect -1916 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 36234 328102
rect 36290 328046 36358 328102
rect 36414 328046 36482 328102
rect 36538 328046 36606 328102
rect 36662 328046 66954 328102
rect 67010 328046 67078 328102
rect 67134 328046 67202 328102
rect 67258 328046 67326 328102
rect 67382 328046 97674 328102
rect 97730 328046 97798 328102
rect 97854 328046 97922 328102
rect 97978 328046 98046 328102
rect 98102 328046 128394 328102
rect 128450 328046 128518 328102
rect 128574 328046 128642 328102
rect 128698 328046 128766 328102
rect 128822 328046 154518 328102
rect 154574 328046 154642 328102
rect 154698 328046 159114 328102
rect 159170 328046 159238 328102
rect 159294 328046 159362 328102
rect 159418 328046 159486 328102
rect 159542 328046 185238 328102
rect 185294 328046 185362 328102
rect 185418 328046 189834 328102
rect 189890 328046 189958 328102
rect 190014 328046 190082 328102
rect 190138 328046 190206 328102
rect 190262 328046 220554 328102
rect 220610 328046 220678 328102
rect 220734 328046 220802 328102
rect 220858 328046 220926 328102
rect 220982 328046 240518 328102
rect 240574 328046 240642 328102
rect 240698 328046 271238 328102
rect 271294 328046 271362 328102
rect 271418 328046 301958 328102
rect 302014 328046 302082 328102
rect 302138 328046 332678 328102
rect 332734 328046 332802 328102
rect 332858 328046 363398 328102
rect 363454 328046 363522 328102
rect 363578 328046 404874 328102
rect 404930 328046 404998 328102
rect 405054 328046 405122 328102
rect 405178 328046 405246 328102
rect 405302 328046 435594 328102
rect 435650 328046 435718 328102
rect 435774 328046 435842 328102
rect 435898 328046 435966 328102
rect 436022 328046 466314 328102
rect 466370 328046 466438 328102
rect 466494 328046 466562 328102
rect 466618 328046 466686 328102
rect 466742 328046 497034 328102
rect 497090 328046 497158 328102
rect 497214 328046 497282 328102
rect 497338 328046 497406 328102
rect 497462 328046 527754 328102
rect 527810 328046 527878 328102
rect 527934 328046 528002 328102
rect 528058 328046 528126 328102
rect 528182 328046 558474 328102
rect 558530 328046 558598 328102
rect 558654 328046 558722 328102
rect 558778 328046 558846 328102
rect 558902 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597980 328102
rect -1916 327978 597980 328046
rect -1916 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 36234 327978
rect 36290 327922 36358 327978
rect 36414 327922 36482 327978
rect 36538 327922 36606 327978
rect 36662 327922 66954 327978
rect 67010 327922 67078 327978
rect 67134 327922 67202 327978
rect 67258 327922 67326 327978
rect 67382 327922 97674 327978
rect 97730 327922 97798 327978
rect 97854 327922 97922 327978
rect 97978 327922 98046 327978
rect 98102 327922 128394 327978
rect 128450 327922 128518 327978
rect 128574 327922 128642 327978
rect 128698 327922 128766 327978
rect 128822 327922 154518 327978
rect 154574 327922 154642 327978
rect 154698 327922 159114 327978
rect 159170 327922 159238 327978
rect 159294 327922 159362 327978
rect 159418 327922 159486 327978
rect 159542 327922 185238 327978
rect 185294 327922 185362 327978
rect 185418 327922 189834 327978
rect 189890 327922 189958 327978
rect 190014 327922 190082 327978
rect 190138 327922 190206 327978
rect 190262 327922 220554 327978
rect 220610 327922 220678 327978
rect 220734 327922 220802 327978
rect 220858 327922 220926 327978
rect 220982 327922 240518 327978
rect 240574 327922 240642 327978
rect 240698 327922 271238 327978
rect 271294 327922 271362 327978
rect 271418 327922 301958 327978
rect 302014 327922 302082 327978
rect 302138 327922 332678 327978
rect 332734 327922 332802 327978
rect 332858 327922 363398 327978
rect 363454 327922 363522 327978
rect 363578 327922 404874 327978
rect 404930 327922 404998 327978
rect 405054 327922 405122 327978
rect 405178 327922 405246 327978
rect 405302 327922 435594 327978
rect 435650 327922 435718 327978
rect 435774 327922 435842 327978
rect 435898 327922 435966 327978
rect 436022 327922 466314 327978
rect 466370 327922 466438 327978
rect 466494 327922 466562 327978
rect 466618 327922 466686 327978
rect 466742 327922 497034 327978
rect 497090 327922 497158 327978
rect 497214 327922 497282 327978
rect 497338 327922 497406 327978
rect 497462 327922 527754 327978
rect 527810 327922 527878 327978
rect 527934 327922 528002 327978
rect 528058 327922 528126 327978
rect 528182 327922 558474 327978
rect 558530 327922 558598 327978
rect 558654 327922 558722 327978
rect 558778 327922 558846 327978
rect 558902 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597980 327978
rect -1916 327826 597980 327922
rect -1916 316350 597980 316446
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 9234 316350
rect 9290 316294 9358 316350
rect 9414 316294 9482 316350
rect 9538 316294 9606 316350
rect 9662 316294 39954 316350
rect 40010 316294 40078 316350
rect 40134 316294 40202 316350
rect 40258 316294 40326 316350
rect 40382 316294 70674 316350
rect 70730 316294 70798 316350
rect 70854 316294 70922 316350
rect 70978 316294 71046 316350
rect 71102 316294 101394 316350
rect 101450 316294 101518 316350
rect 101574 316294 101642 316350
rect 101698 316294 101766 316350
rect 101822 316294 132114 316350
rect 132170 316294 132238 316350
rect 132294 316294 132362 316350
rect 132418 316294 132486 316350
rect 132542 316294 162834 316350
rect 162890 316294 162958 316350
rect 163014 316294 163082 316350
rect 163138 316294 163206 316350
rect 163262 316294 193554 316350
rect 193610 316294 193678 316350
rect 193734 316294 193802 316350
rect 193858 316294 193926 316350
rect 193982 316294 224274 316350
rect 224330 316294 224398 316350
rect 224454 316294 224522 316350
rect 224578 316294 224646 316350
rect 224702 316294 255878 316350
rect 255934 316294 256002 316350
rect 256058 316294 286598 316350
rect 286654 316294 286722 316350
rect 286778 316294 317318 316350
rect 317374 316294 317442 316350
rect 317498 316294 348038 316350
rect 348094 316294 348162 316350
rect 348218 316294 377874 316350
rect 377930 316294 377998 316350
rect 378054 316294 378122 316350
rect 378178 316294 378246 316350
rect 378302 316294 408594 316350
rect 408650 316294 408718 316350
rect 408774 316294 408842 316350
rect 408898 316294 408966 316350
rect 409022 316294 439314 316350
rect 439370 316294 439438 316350
rect 439494 316294 439562 316350
rect 439618 316294 439686 316350
rect 439742 316294 470034 316350
rect 470090 316294 470158 316350
rect 470214 316294 470282 316350
rect 470338 316294 470406 316350
rect 470462 316294 500754 316350
rect 500810 316294 500878 316350
rect 500934 316294 501002 316350
rect 501058 316294 501126 316350
rect 501182 316294 531474 316350
rect 531530 316294 531598 316350
rect 531654 316294 531722 316350
rect 531778 316294 531846 316350
rect 531902 316294 562194 316350
rect 562250 316294 562318 316350
rect 562374 316294 562442 316350
rect 562498 316294 562566 316350
rect 562622 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect -1916 316226 597980 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 9234 316226
rect 9290 316170 9358 316226
rect 9414 316170 9482 316226
rect 9538 316170 9606 316226
rect 9662 316170 39954 316226
rect 40010 316170 40078 316226
rect 40134 316170 40202 316226
rect 40258 316170 40326 316226
rect 40382 316170 70674 316226
rect 70730 316170 70798 316226
rect 70854 316170 70922 316226
rect 70978 316170 71046 316226
rect 71102 316170 101394 316226
rect 101450 316170 101518 316226
rect 101574 316170 101642 316226
rect 101698 316170 101766 316226
rect 101822 316170 132114 316226
rect 132170 316170 132238 316226
rect 132294 316170 132362 316226
rect 132418 316170 132486 316226
rect 132542 316170 162834 316226
rect 162890 316170 162958 316226
rect 163014 316170 163082 316226
rect 163138 316170 163206 316226
rect 163262 316170 193554 316226
rect 193610 316170 193678 316226
rect 193734 316170 193802 316226
rect 193858 316170 193926 316226
rect 193982 316170 224274 316226
rect 224330 316170 224398 316226
rect 224454 316170 224522 316226
rect 224578 316170 224646 316226
rect 224702 316170 255878 316226
rect 255934 316170 256002 316226
rect 256058 316170 286598 316226
rect 286654 316170 286722 316226
rect 286778 316170 317318 316226
rect 317374 316170 317442 316226
rect 317498 316170 348038 316226
rect 348094 316170 348162 316226
rect 348218 316170 377874 316226
rect 377930 316170 377998 316226
rect 378054 316170 378122 316226
rect 378178 316170 378246 316226
rect 378302 316170 408594 316226
rect 408650 316170 408718 316226
rect 408774 316170 408842 316226
rect 408898 316170 408966 316226
rect 409022 316170 439314 316226
rect 439370 316170 439438 316226
rect 439494 316170 439562 316226
rect 439618 316170 439686 316226
rect 439742 316170 470034 316226
rect 470090 316170 470158 316226
rect 470214 316170 470282 316226
rect 470338 316170 470406 316226
rect 470462 316170 500754 316226
rect 500810 316170 500878 316226
rect 500934 316170 501002 316226
rect 501058 316170 501126 316226
rect 501182 316170 531474 316226
rect 531530 316170 531598 316226
rect 531654 316170 531722 316226
rect 531778 316170 531846 316226
rect 531902 316170 562194 316226
rect 562250 316170 562318 316226
rect 562374 316170 562442 316226
rect 562498 316170 562566 316226
rect 562622 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect -1916 316102 597980 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 9234 316102
rect 9290 316046 9358 316102
rect 9414 316046 9482 316102
rect 9538 316046 9606 316102
rect 9662 316046 39954 316102
rect 40010 316046 40078 316102
rect 40134 316046 40202 316102
rect 40258 316046 40326 316102
rect 40382 316046 70674 316102
rect 70730 316046 70798 316102
rect 70854 316046 70922 316102
rect 70978 316046 71046 316102
rect 71102 316046 101394 316102
rect 101450 316046 101518 316102
rect 101574 316046 101642 316102
rect 101698 316046 101766 316102
rect 101822 316046 132114 316102
rect 132170 316046 132238 316102
rect 132294 316046 132362 316102
rect 132418 316046 132486 316102
rect 132542 316046 162834 316102
rect 162890 316046 162958 316102
rect 163014 316046 163082 316102
rect 163138 316046 163206 316102
rect 163262 316046 193554 316102
rect 193610 316046 193678 316102
rect 193734 316046 193802 316102
rect 193858 316046 193926 316102
rect 193982 316046 224274 316102
rect 224330 316046 224398 316102
rect 224454 316046 224522 316102
rect 224578 316046 224646 316102
rect 224702 316046 255878 316102
rect 255934 316046 256002 316102
rect 256058 316046 286598 316102
rect 286654 316046 286722 316102
rect 286778 316046 317318 316102
rect 317374 316046 317442 316102
rect 317498 316046 348038 316102
rect 348094 316046 348162 316102
rect 348218 316046 377874 316102
rect 377930 316046 377998 316102
rect 378054 316046 378122 316102
rect 378178 316046 378246 316102
rect 378302 316046 408594 316102
rect 408650 316046 408718 316102
rect 408774 316046 408842 316102
rect 408898 316046 408966 316102
rect 409022 316046 439314 316102
rect 439370 316046 439438 316102
rect 439494 316046 439562 316102
rect 439618 316046 439686 316102
rect 439742 316046 470034 316102
rect 470090 316046 470158 316102
rect 470214 316046 470282 316102
rect 470338 316046 470406 316102
rect 470462 316046 500754 316102
rect 500810 316046 500878 316102
rect 500934 316046 501002 316102
rect 501058 316046 501126 316102
rect 501182 316046 531474 316102
rect 531530 316046 531598 316102
rect 531654 316046 531722 316102
rect 531778 316046 531846 316102
rect 531902 316046 562194 316102
rect 562250 316046 562318 316102
rect 562374 316046 562442 316102
rect 562498 316046 562566 316102
rect 562622 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect -1916 315978 597980 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 9234 315978
rect 9290 315922 9358 315978
rect 9414 315922 9482 315978
rect 9538 315922 9606 315978
rect 9662 315922 39954 315978
rect 40010 315922 40078 315978
rect 40134 315922 40202 315978
rect 40258 315922 40326 315978
rect 40382 315922 70674 315978
rect 70730 315922 70798 315978
rect 70854 315922 70922 315978
rect 70978 315922 71046 315978
rect 71102 315922 101394 315978
rect 101450 315922 101518 315978
rect 101574 315922 101642 315978
rect 101698 315922 101766 315978
rect 101822 315922 132114 315978
rect 132170 315922 132238 315978
rect 132294 315922 132362 315978
rect 132418 315922 132486 315978
rect 132542 315922 162834 315978
rect 162890 315922 162958 315978
rect 163014 315922 163082 315978
rect 163138 315922 163206 315978
rect 163262 315922 193554 315978
rect 193610 315922 193678 315978
rect 193734 315922 193802 315978
rect 193858 315922 193926 315978
rect 193982 315922 224274 315978
rect 224330 315922 224398 315978
rect 224454 315922 224522 315978
rect 224578 315922 224646 315978
rect 224702 315922 255878 315978
rect 255934 315922 256002 315978
rect 256058 315922 286598 315978
rect 286654 315922 286722 315978
rect 286778 315922 317318 315978
rect 317374 315922 317442 315978
rect 317498 315922 348038 315978
rect 348094 315922 348162 315978
rect 348218 315922 377874 315978
rect 377930 315922 377998 315978
rect 378054 315922 378122 315978
rect 378178 315922 378246 315978
rect 378302 315922 408594 315978
rect 408650 315922 408718 315978
rect 408774 315922 408842 315978
rect 408898 315922 408966 315978
rect 409022 315922 439314 315978
rect 439370 315922 439438 315978
rect 439494 315922 439562 315978
rect 439618 315922 439686 315978
rect 439742 315922 470034 315978
rect 470090 315922 470158 315978
rect 470214 315922 470282 315978
rect 470338 315922 470406 315978
rect 470462 315922 500754 315978
rect 500810 315922 500878 315978
rect 500934 315922 501002 315978
rect 501058 315922 501126 315978
rect 501182 315922 531474 315978
rect 531530 315922 531598 315978
rect 531654 315922 531722 315978
rect 531778 315922 531846 315978
rect 531902 315922 562194 315978
rect 562250 315922 562318 315978
rect 562374 315922 562442 315978
rect 562498 315922 562566 315978
rect 562622 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect -1916 315826 597980 315922
rect -1916 310350 597980 310446
rect -1916 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 36234 310350
rect 36290 310294 36358 310350
rect 36414 310294 36482 310350
rect 36538 310294 36606 310350
rect 36662 310294 66954 310350
rect 67010 310294 67078 310350
rect 67134 310294 67202 310350
rect 67258 310294 67326 310350
rect 67382 310294 97674 310350
rect 97730 310294 97798 310350
rect 97854 310294 97922 310350
rect 97978 310294 98046 310350
rect 98102 310294 128394 310350
rect 128450 310294 128518 310350
rect 128574 310294 128642 310350
rect 128698 310294 128766 310350
rect 128822 310294 159114 310350
rect 159170 310294 159238 310350
rect 159294 310294 159362 310350
rect 159418 310294 159486 310350
rect 159542 310294 189834 310350
rect 189890 310294 189958 310350
rect 190014 310294 190082 310350
rect 190138 310294 190206 310350
rect 190262 310294 220554 310350
rect 220610 310294 220678 310350
rect 220734 310294 220802 310350
rect 220858 310294 220926 310350
rect 220982 310294 240518 310350
rect 240574 310294 240642 310350
rect 240698 310294 271238 310350
rect 271294 310294 271362 310350
rect 271418 310294 301958 310350
rect 302014 310294 302082 310350
rect 302138 310294 332678 310350
rect 332734 310294 332802 310350
rect 332858 310294 363398 310350
rect 363454 310294 363522 310350
rect 363578 310294 404874 310350
rect 404930 310294 404998 310350
rect 405054 310294 405122 310350
rect 405178 310294 405246 310350
rect 405302 310294 435594 310350
rect 435650 310294 435718 310350
rect 435774 310294 435842 310350
rect 435898 310294 435966 310350
rect 436022 310294 466314 310350
rect 466370 310294 466438 310350
rect 466494 310294 466562 310350
rect 466618 310294 466686 310350
rect 466742 310294 497034 310350
rect 497090 310294 497158 310350
rect 497214 310294 497282 310350
rect 497338 310294 497406 310350
rect 497462 310294 527754 310350
rect 527810 310294 527878 310350
rect 527934 310294 528002 310350
rect 528058 310294 528126 310350
rect 528182 310294 558474 310350
rect 558530 310294 558598 310350
rect 558654 310294 558722 310350
rect 558778 310294 558846 310350
rect 558902 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597980 310350
rect -1916 310226 597980 310294
rect -1916 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 36234 310226
rect 36290 310170 36358 310226
rect 36414 310170 36482 310226
rect 36538 310170 36606 310226
rect 36662 310170 66954 310226
rect 67010 310170 67078 310226
rect 67134 310170 67202 310226
rect 67258 310170 67326 310226
rect 67382 310170 97674 310226
rect 97730 310170 97798 310226
rect 97854 310170 97922 310226
rect 97978 310170 98046 310226
rect 98102 310170 128394 310226
rect 128450 310170 128518 310226
rect 128574 310170 128642 310226
rect 128698 310170 128766 310226
rect 128822 310170 159114 310226
rect 159170 310170 159238 310226
rect 159294 310170 159362 310226
rect 159418 310170 159486 310226
rect 159542 310170 189834 310226
rect 189890 310170 189958 310226
rect 190014 310170 190082 310226
rect 190138 310170 190206 310226
rect 190262 310170 220554 310226
rect 220610 310170 220678 310226
rect 220734 310170 220802 310226
rect 220858 310170 220926 310226
rect 220982 310170 240518 310226
rect 240574 310170 240642 310226
rect 240698 310170 271238 310226
rect 271294 310170 271362 310226
rect 271418 310170 301958 310226
rect 302014 310170 302082 310226
rect 302138 310170 332678 310226
rect 332734 310170 332802 310226
rect 332858 310170 363398 310226
rect 363454 310170 363522 310226
rect 363578 310170 404874 310226
rect 404930 310170 404998 310226
rect 405054 310170 405122 310226
rect 405178 310170 405246 310226
rect 405302 310170 435594 310226
rect 435650 310170 435718 310226
rect 435774 310170 435842 310226
rect 435898 310170 435966 310226
rect 436022 310170 466314 310226
rect 466370 310170 466438 310226
rect 466494 310170 466562 310226
rect 466618 310170 466686 310226
rect 466742 310170 497034 310226
rect 497090 310170 497158 310226
rect 497214 310170 497282 310226
rect 497338 310170 497406 310226
rect 497462 310170 527754 310226
rect 527810 310170 527878 310226
rect 527934 310170 528002 310226
rect 528058 310170 528126 310226
rect 528182 310170 558474 310226
rect 558530 310170 558598 310226
rect 558654 310170 558722 310226
rect 558778 310170 558846 310226
rect 558902 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597980 310226
rect -1916 310102 597980 310170
rect -1916 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 36234 310102
rect 36290 310046 36358 310102
rect 36414 310046 36482 310102
rect 36538 310046 36606 310102
rect 36662 310046 66954 310102
rect 67010 310046 67078 310102
rect 67134 310046 67202 310102
rect 67258 310046 67326 310102
rect 67382 310046 97674 310102
rect 97730 310046 97798 310102
rect 97854 310046 97922 310102
rect 97978 310046 98046 310102
rect 98102 310046 128394 310102
rect 128450 310046 128518 310102
rect 128574 310046 128642 310102
rect 128698 310046 128766 310102
rect 128822 310046 159114 310102
rect 159170 310046 159238 310102
rect 159294 310046 159362 310102
rect 159418 310046 159486 310102
rect 159542 310046 189834 310102
rect 189890 310046 189958 310102
rect 190014 310046 190082 310102
rect 190138 310046 190206 310102
rect 190262 310046 220554 310102
rect 220610 310046 220678 310102
rect 220734 310046 220802 310102
rect 220858 310046 220926 310102
rect 220982 310046 240518 310102
rect 240574 310046 240642 310102
rect 240698 310046 271238 310102
rect 271294 310046 271362 310102
rect 271418 310046 301958 310102
rect 302014 310046 302082 310102
rect 302138 310046 332678 310102
rect 332734 310046 332802 310102
rect 332858 310046 363398 310102
rect 363454 310046 363522 310102
rect 363578 310046 404874 310102
rect 404930 310046 404998 310102
rect 405054 310046 405122 310102
rect 405178 310046 405246 310102
rect 405302 310046 435594 310102
rect 435650 310046 435718 310102
rect 435774 310046 435842 310102
rect 435898 310046 435966 310102
rect 436022 310046 466314 310102
rect 466370 310046 466438 310102
rect 466494 310046 466562 310102
rect 466618 310046 466686 310102
rect 466742 310046 497034 310102
rect 497090 310046 497158 310102
rect 497214 310046 497282 310102
rect 497338 310046 497406 310102
rect 497462 310046 527754 310102
rect 527810 310046 527878 310102
rect 527934 310046 528002 310102
rect 528058 310046 528126 310102
rect 528182 310046 558474 310102
rect 558530 310046 558598 310102
rect 558654 310046 558722 310102
rect 558778 310046 558846 310102
rect 558902 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597980 310102
rect -1916 309978 597980 310046
rect -1916 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 36234 309978
rect 36290 309922 36358 309978
rect 36414 309922 36482 309978
rect 36538 309922 36606 309978
rect 36662 309922 66954 309978
rect 67010 309922 67078 309978
rect 67134 309922 67202 309978
rect 67258 309922 67326 309978
rect 67382 309922 97674 309978
rect 97730 309922 97798 309978
rect 97854 309922 97922 309978
rect 97978 309922 98046 309978
rect 98102 309922 128394 309978
rect 128450 309922 128518 309978
rect 128574 309922 128642 309978
rect 128698 309922 128766 309978
rect 128822 309922 159114 309978
rect 159170 309922 159238 309978
rect 159294 309922 159362 309978
rect 159418 309922 159486 309978
rect 159542 309922 189834 309978
rect 189890 309922 189958 309978
rect 190014 309922 190082 309978
rect 190138 309922 190206 309978
rect 190262 309922 220554 309978
rect 220610 309922 220678 309978
rect 220734 309922 220802 309978
rect 220858 309922 220926 309978
rect 220982 309922 240518 309978
rect 240574 309922 240642 309978
rect 240698 309922 271238 309978
rect 271294 309922 271362 309978
rect 271418 309922 301958 309978
rect 302014 309922 302082 309978
rect 302138 309922 332678 309978
rect 332734 309922 332802 309978
rect 332858 309922 363398 309978
rect 363454 309922 363522 309978
rect 363578 309922 404874 309978
rect 404930 309922 404998 309978
rect 405054 309922 405122 309978
rect 405178 309922 405246 309978
rect 405302 309922 435594 309978
rect 435650 309922 435718 309978
rect 435774 309922 435842 309978
rect 435898 309922 435966 309978
rect 436022 309922 466314 309978
rect 466370 309922 466438 309978
rect 466494 309922 466562 309978
rect 466618 309922 466686 309978
rect 466742 309922 497034 309978
rect 497090 309922 497158 309978
rect 497214 309922 497282 309978
rect 497338 309922 497406 309978
rect 497462 309922 527754 309978
rect 527810 309922 527878 309978
rect 527934 309922 528002 309978
rect 528058 309922 528126 309978
rect 528182 309922 558474 309978
rect 558530 309922 558598 309978
rect 558654 309922 558722 309978
rect 558778 309922 558846 309978
rect 558902 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597980 309978
rect -1916 309826 597980 309922
rect -1916 298422 597980 298446
rect -1916 298366 70674 298422
rect 70730 298366 70798 298422
rect 70854 298366 70922 298422
rect 70978 298366 71046 298422
rect 71102 298366 597980 298422
rect -1916 298350 597980 298366
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 9234 298350
rect 9290 298294 9358 298350
rect 9414 298294 9482 298350
rect 9538 298294 9606 298350
rect 9662 298294 39954 298350
rect 40010 298294 40078 298350
rect 40134 298294 40202 298350
rect 40258 298294 40326 298350
rect 40382 298298 101394 298350
rect 40382 298294 70674 298298
rect -1916 298242 70674 298294
rect 70730 298242 70798 298298
rect 70854 298242 70922 298298
rect 70978 298242 71046 298298
rect 71102 298294 101394 298298
rect 101450 298294 101518 298350
rect 101574 298294 101642 298350
rect 101698 298294 101766 298350
rect 101822 298294 132114 298350
rect 132170 298294 132238 298350
rect 132294 298294 132362 298350
rect 132418 298294 132486 298350
rect 132542 298294 162834 298350
rect 162890 298294 162958 298350
rect 163014 298294 163082 298350
rect 163138 298294 163206 298350
rect 163262 298294 193554 298350
rect 193610 298294 193678 298350
rect 193734 298294 193802 298350
rect 193858 298294 193926 298350
rect 193982 298294 224274 298350
rect 224330 298294 224398 298350
rect 224454 298294 224522 298350
rect 224578 298294 224646 298350
rect 224702 298294 255878 298350
rect 255934 298294 256002 298350
rect 256058 298294 286598 298350
rect 286654 298294 286722 298350
rect 286778 298294 317318 298350
rect 317374 298294 317442 298350
rect 317498 298294 348038 298350
rect 348094 298294 348162 298350
rect 348218 298294 377874 298350
rect 377930 298294 377998 298350
rect 378054 298294 378122 298350
rect 378178 298294 378246 298350
rect 378302 298294 408594 298350
rect 408650 298294 408718 298350
rect 408774 298294 408842 298350
rect 408898 298294 408966 298350
rect 409022 298294 439314 298350
rect 439370 298294 439438 298350
rect 439494 298294 439562 298350
rect 439618 298294 439686 298350
rect 439742 298294 470034 298350
rect 470090 298294 470158 298350
rect 470214 298294 470282 298350
rect 470338 298294 470406 298350
rect 470462 298294 500754 298350
rect 500810 298294 500878 298350
rect 500934 298294 501002 298350
rect 501058 298294 501126 298350
rect 501182 298294 531474 298350
rect 531530 298294 531598 298350
rect 531654 298294 531722 298350
rect 531778 298294 531846 298350
rect 531902 298294 562194 298350
rect 562250 298294 562318 298350
rect 562374 298294 562442 298350
rect 562498 298294 562566 298350
rect 562622 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect 71102 298242 597980 298294
rect -1916 298226 597980 298242
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 9234 298226
rect 9290 298170 9358 298226
rect 9414 298170 9482 298226
rect 9538 298170 9606 298226
rect 9662 298170 39954 298226
rect 40010 298170 40078 298226
rect 40134 298170 40202 298226
rect 40258 298170 40326 298226
rect 40382 298174 101394 298226
rect 40382 298170 70674 298174
rect -1916 298118 70674 298170
rect 70730 298118 70798 298174
rect 70854 298118 70922 298174
rect 70978 298118 71046 298174
rect 71102 298170 101394 298174
rect 101450 298170 101518 298226
rect 101574 298170 101642 298226
rect 101698 298170 101766 298226
rect 101822 298170 132114 298226
rect 132170 298170 132238 298226
rect 132294 298170 132362 298226
rect 132418 298170 132486 298226
rect 132542 298170 162834 298226
rect 162890 298170 162958 298226
rect 163014 298170 163082 298226
rect 163138 298170 163206 298226
rect 163262 298170 193554 298226
rect 193610 298170 193678 298226
rect 193734 298170 193802 298226
rect 193858 298170 193926 298226
rect 193982 298170 224274 298226
rect 224330 298170 224398 298226
rect 224454 298170 224522 298226
rect 224578 298170 224646 298226
rect 224702 298170 255878 298226
rect 255934 298170 256002 298226
rect 256058 298170 286598 298226
rect 286654 298170 286722 298226
rect 286778 298170 317318 298226
rect 317374 298170 317442 298226
rect 317498 298170 348038 298226
rect 348094 298170 348162 298226
rect 348218 298170 377874 298226
rect 377930 298170 377998 298226
rect 378054 298170 378122 298226
rect 378178 298170 378246 298226
rect 378302 298170 408594 298226
rect 408650 298170 408718 298226
rect 408774 298170 408842 298226
rect 408898 298170 408966 298226
rect 409022 298170 439314 298226
rect 439370 298170 439438 298226
rect 439494 298170 439562 298226
rect 439618 298170 439686 298226
rect 439742 298170 470034 298226
rect 470090 298170 470158 298226
rect 470214 298170 470282 298226
rect 470338 298170 470406 298226
rect 470462 298170 500754 298226
rect 500810 298170 500878 298226
rect 500934 298170 501002 298226
rect 501058 298170 501126 298226
rect 501182 298170 531474 298226
rect 531530 298170 531598 298226
rect 531654 298170 531722 298226
rect 531778 298170 531846 298226
rect 531902 298170 562194 298226
rect 562250 298170 562318 298226
rect 562374 298170 562442 298226
rect 562498 298170 562566 298226
rect 562622 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect 71102 298118 597980 298170
rect -1916 298102 597980 298118
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 9234 298102
rect 9290 298046 9358 298102
rect 9414 298046 9482 298102
rect 9538 298046 9606 298102
rect 9662 298046 39954 298102
rect 40010 298046 40078 298102
rect 40134 298046 40202 298102
rect 40258 298046 40326 298102
rect 40382 298046 101394 298102
rect 101450 298046 101518 298102
rect 101574 298046 101642 298102
rect 101698 298046 101766 298102
rect 101822 298046 132114 298102
rect 132170 298046 132238 298102
rect 132294 298046 132362 298102
rect 132418 298046 132486 298102
rect 132542 298046 162834 298102
rect 162890 298046 162958 298102
rect 163014 298046 163082 298102
rect 163138 298046 163206 298102
rect 163262 298046 193554 298102
rect 193610 298046 193678 298102
rect 193734 298046 193802 298102
rect 193858 298046 193926 298102
rect 193982 298046 224274 298102
rect 224330 298046 224398 298102
rect 224454 298046 224522 298102
rect 224578 298046 224646 298102
rect 224702 298046 255878 298102
rect 255934 298046 256002 298102
rect 256058 298046 286598 298102
rect 286654 298046 286722 298102
rect 286778 298046 317318 298102
rect 317374 298046 317442 298102
rect 317498 298046 348038 298102
rect 348094 298046 348162 298102
rect 348218 298046 377874 298102
rect 377930 298046 377998 298102
rect 378054 298046 378122 298102
rect 378178 298046 378246 298102
rect 378302 298046 408594 298102
rect 408650 298046 408718 298102
rect 408774 298046 408842 298102
rect 408898 298046 408966 298102
rect 409022 298046 439314 298102
rect 439370 298046 439438 298102
rect 439494 298046 439562 298102
rect 439618 298046 439686 298102
rect 439742 298046 470034 298102
rect 470090 298046 470158 298102
rect 470214 298046 470282 298102
rect 470338 298046 470406 298102
rect 470462 298046 500754 298102
rect 500810 298046 500878 298102
rect 500934 298046 501002 298102
rect 501058 298046 501126 298102
rect 501182 298046 531474 298102
rect 531530 298046 531598 298102
rect 531654 298046 531722 298102
rect 531778 298046 531846 298102
rect 531902 298046 562194 298102
rect 562250 298046 562318 298102
rect 562374 298046 562442 298102
rect 562498 298046 562566 298102
rect 562622 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect -1916 297978 597980 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 9234 297978
rect 9290 297922 9358 297978
rect 9414 297922 9482 297978
rect 9538 297922 9606 297978
rect 9662 297922 39954 297978
rect 40010 297922 40078 297978
rect 40134 297922 40202 297978
rect 40258 297922 40326 297978
rect 40382 297922 101394 297978
rect 101450 297922 101518 297978
rect 101574 297922 101642 297978
rect 101698 297922 101766 297978
rect 101822 297922 132114 297978
rect 132170 297922 132238 297978
rect 132294 297922 132362 297978
rect 132418 297922 132486 297978
rect 132542 297922 162834 297978
rect 162890 297922 162958 297978
rect 163014 297922 163082 297978
rect 163138 297922 163206 297978
rect 163262 297922 193554 297978
rect 193610 297922 193678 297978
rect 193734 297922 193802 297978
rect 193858 297922 193926 297978
rect 193982 297922 224274 297978
rect 224330 297922 224398 297978
rect 224454 297922 224522 297978
rect 224578 297922 224646 297978
rect 224702 297922 255878 297978
rect 255934 297922 256002 297978
rect 256058 297922 286598 297978
rect 286654 297922 286722 297978
rect 286778 297922 317318 297978
rect 317374 297922 317442 297978
rect 317498 297922 348038 297978
rect 348094 297922 348162 297978
rect 348218 297922 377874 297978
rect 377930 297922 377998 297978
rect 378054 297922 378122 297978
rect 378178 297922 378246 297978
rect 378302 297922 408594 297978
rect 408650 297922 408718 297978
rect 408774 297922 408842 297978
rect 408898 297922 408966 297978
rect 409022 297922 439314 297978
rect 439370 297922 439438 297978
rect 439494 297922 439562 297978
rect 439618 297922 439686 297978
rect 439742 297922 470034 297978
rect 470090 297922 470158 297978
rect 470214 297922 470282 297978
rect 470338 297922 470406 297978
rect 470462 297922 500754 297978
rect 500810 297922 500878 297978
rect 500934 297922 501002 297978
rect 501058 297922 501126 297978
rect 501182 297922 531474 297978
rect 531530 297922 531598 297978
rect 531654 297922 531722 297978
rect 531778 297922 531846 297978
rect 531902 297922 562194 297978
rect 562250 297922 562318 297978
rect 562374 297922 562442 297978
rect 562498 297922 562566 297978
rect 562622 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect -1916 297826 597980 297922
rect -1916 292350 597980 292446
rect -1916 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 36234 292350
rect 36290 292294 36358 292350
rect 36414 292294 36482 292350
rect 36538 292294 36606 292350
rect 36662 292294 44518 292350
rect 44574 292294 44642 292350
rect 44698 292294 75238 292350
rect 75294 292294 75362 292350
rect 75418 292294 97674 292350
rect 97730 292294 97798 292350
rect 97854 292294 97922 292350
rect 97978 292294 98046 292350
rect 98102 292294 128394 292350
rect 128450 292294 128518 292350
rect 128574 292294 128642 292350
rect 128698 292294 128766 292350
rect 128822 292294 159114 292350
rect 159170 292294 159238 292350
rect 159294 292294 159362 292350
rect 159418 292294 159486 292350
rect 159542 292294 189834 292350
rect 189890 292294 189958 292350
rect 190014 292294 190082 292350
rect 190138 292294 190206 292350
rect 190262 292294 220554 292350
rect 220610 292294 220678 292350
rect 220734 292294 220802 292350
rect 220858 292294 220926 292350
rect 220982 292294 240518 292350
rect 240574 292294 240642 292350
rect 240698 292294 271238 292350
rect 271294 292294 271362 292350
rect 271418 292294 301958 292350
rect 302014 292294 302082 292350
rect 302138 292294 332678 292350
rect 332734 292294 332802 292350
rect 332858 292294 363398 292350
rect 363454 292294 363522 292350
rect 363578 292294 404874 292350
rect 404930 292294 404998 292350
rect 405054 292294 405122 292350
rect 405178 292294 405246 292350
rect 405302 292294 435594 292350
rect 435650 292294 435718 292350
rect 435774 292294 435842 292350
rect 435898 292294 435966 292350
rect 436022 292294 466314 292350
rect 466370 292294 466438 292350
rect 466494 292294 466562 292350
rect 466618 292294 466686 292350
rect 466742 292294 497034 292350
rect 497090 292294 497158 292350
rect 497214 292294 497282 292350
rect 497338 292294 497406 292350
rect 497462 292294 527754 292350
rect 527810 292294 527878 292350
rect 527934 292294 528002 292350
rect 528058 292294 528126 292350
rect 528182 292294 558474 292350
rect 558530 292294 558598 292350
rect 558654 292294 558722 292350
rect 558778 292294 558846 292350
rect 558902 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597980 292350
rect -1916 292226 597980 292294
rect -1916 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 36234 292226
rect 36290 292170 36358 292226
rect 36414 292170 36482 292226
rect 36538 292170 36606 292226
rect 36662 292170 44518 292226
rect 44574 292170 44642 292226
rect 44698 292170 75238 292226
rect 75294 292170 75362 292226
rect 75418 292170 97674 292226
rect 97730 292170 97798 292226
rect 97854 292170 97922 292226
rect 97978 292170 98046 292226
rect 98102 292170 128394 292226
rect 128450 292170 128518 292226
rect 128574 292170 128642 292226
rect 128698 292170 128766 292226
rect 128822 292170 159114 292226
rect 159170 292170 159238 292226
rect 159294 292170 159362 292226
rect 159418 292170 159486 292226
rect 159542 292170 189834 292226
rect 189890 292170 189958 292226
rect 190014 292170 190082 292226
rect 190138 292170 190206 292226
rect 190262 292170 220554 292226
rect 220610 292170 220678 292226
rect 220734 292170 220802 292226
rect 220858 292170 220926 292226
rect 220982 292170 240518 292226
rect 240574 292170 240642 292226
rect 240698 292170 271238 292226
rect 271294 292170 271362 292226
rect 271418 292170 301958 292226
rect 302014 292170 302082 292226
rect 302138 292170 332678 292226
rect 332734 292170 332802 292226
rect 332858 292170 363398 292226
rect 363454 292170 363522 292226
rect 363578 292170 404874 292226
rect 404930 292170 404998 292226
rect 405054 292170 405122 292226
rect 405178 292170 405246 292226
rect 405302 292170 435594 292226
rect 435650 292170 435718 292226
rect 435774 292170 435842 292226
rect 435898 292170 435966 292226
rect 436022 292170 466314 292226
rect 466370 292170 466438 292226
rect 466494 292170 466562 292226
rect 466618 292170 466686 292226
rect 466742 292170 497034 292226
rect 497090 292170 497158 292226
rect 497214 292170 497282 292226
rect 497338 292170 497406 292226
rect 497462 292170 527754 292226
rect 527810 292170 527878 292226
rect 527934 292170 528002 292226
rect 528058 292170 528126 292226
rect 528182 292170 558474 292226
rect 558530 292170 558598 292226
rect 558654 292170 558722 292226
rect 558778 292170 558846 292226
rect 558902 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597980 292226
rect -1916 292102 597980 292170
rect -1916 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 36234 292102
rect 36290 292046 36358 292102
rect 36414 292046 36482 292102
rect 36538 292046 36606 292102
rect 36662 292046 44518 292102
rect 44574 292046 44642 292102
rect 44698 292046 75238 292102
rect 75294 292046 75362 292102
rect 75418 292046 97674 292102
rect 97730 292046 97798 292102
rect 97854 292046 97922 292102
rect 97978 292046 98046 292102
rect 98102 292046 128394 292102
rect 128450 292046 128518 292102
rect 128574 292046 128642 292102
rect 128698 292046 128766 292102
rect 128822 292046 159114 292102
rect 159170 292046 159238 292102
rect 159294 292046 159362 292102
rect 159418 292046 159486 292102
rect 159542 292046 189834 292102
rect 189890 292046 189958 292102
rect 190014 292046 190082 292102
rect 190138 292046 190206 292102
rect 190262 292046 220554 292102
rect 220610 292046 220678 292102
rect 220734 292046 220802 292102
rect 220858 292046 220926 292102
rect 220982 292046 240518 292102
rect 240574 292046 240642 292102
rect 240698 292046 271238 292102
rect 271294 292046 271362 292102
rect 271418 292046 301958 292102
rect 302014 292046 302082 292102
rect 302138 292046 332678 292102
rect 332734 292046 332802 292102
rect 332858 292046 363398 292102
rect 363454 292046 363522 292102
rect 363578 292046 404874 292102
rect 404930 292046 404998 292102
rect 405054 292046 405122 292102
rect 405178 292046 405246 292102
rect 405302 292046 435594 292102
rect 435650 292046 435718 292102
rect 435774 292046 435842 292102
rect 435898 292046 435966 292102
rect 436022 292046 466314 292102
rect 466370 292046 466438 292102
rect 466494 292046 466562 292102
rect 466618 292046 466686 292102
rect 466742 292046 497034 292102
rect 497090 292046 497158 292102
rect 497214 292046 497282 292102
rect 497338 292046 497406 292102
rect 497462 292046 527754 292102
rect 527810 292046 527878 292102
rect 527934 292046 528002 292102
rect 528058 292046 528126 292102
rect 528182 292046 558474 292102
rect 558530 292046 558598 292102
rect 558654 292046 558722 292102
rect 558778 292046 558846 292102
rect 558902 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597980 292102
rect -1916 291978 597980 292046
rect -1916 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 36234 291978
rect 36290 291922 36358 291978
rect 36414 291922 36482 291978
rect 36538 291922 36606 291978
rect 36662 291922 44518 291978
rect 44574 291922 44642 291978
rect 44698 291922 75238 291978
rect 75294 291922 75362 291978
rect 75418 291922 97674 291978
rect 97730 291922 97798 291978
rect 97854 291922 97922 291978
rect 97978 291922 98046 291978
rect 98102 291922 128394 291978
rect 128450 291922 128518 291978
rect 128574 291922 128642 291978
rect 128698 291922 128766 291978
rect 128822 291922 159114 291978
rect 159170 291922 159238 291978
rect 159294 291922 159362 291978
rect 159418 291922 159486 291978
rect 159542 291922 189834 291978
rect 189890 291922 189958 291978
rect 190014 291922 190082 291978
rect 190138 291922 190206 291978
rect 190262 291922 220554 291978
rect 220610 291922 220678 291978
rect 220734 291922 220802 291978
rect 220858 291922 220926 291978
rect 220982 291922 240518 291978
rect 240574 291922 240642 291978
rect 240698 291922 271238 291978
rect 271294 291922 271362 291978
rect 271418 291922 301958 291978
rect 302014 291922 302082 291978
rect 302138 291922 332678 291978
rect 332734 291922 332802 291978
rect 332858 291922 363398 291978
rect 363454 291922 363522 291978
rect 363578 291922 404874 291978
rect 404930 291922 404998 291978
rect 405054 291922 405122 291978
rect 405178 291922 405246 291978
rect 405302 291922 435594 291978
rect 435650 291922 435718 291978
rect 435774 291922 435842 291978
rect 435898 291922 435966 291978
rect 436022 291922 466314 291978
rect 466370 291922 466438 291978
rect 466494 291922 466562 291978
rect 466618 291922 466686 291978
rect 466742 291922 497034 291978
rect 497090 291922 497158 291978
rect 497214 291922 497282 291978
rect 497338 291922 497406 291978
rect 497462 291922 527754 291978
rect 527810 291922 527878 291978
rect 527934 291922 528002 291978
rect 528058 291922 528126 291978
rect 528182 291922 558474 291978
rect 558530 291922 558598 291978
rect 558654 291922 558722 291978
rect 558778 291922 558846 291978
rect 558902 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597980 291978
rect -1916 291826 597980 291922
rect 373756 288298 375300 288314
rect 373756 288242 373772 288298
rect 373828 288242 375228 288298
rect 375284 288242 375300 288298
rect 373756 288226 375300 288242
rect 373868 286138 375300 286154
rect 373868 286082 373884 286138
rect 373940 286082 375228 286138
rect 375284 286082 375300 286138
rect 373868 286066 375300 286082
rect -1916 280350 597980 280446
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 9234 280350
rect 9290 280294 9358 280350
rect 9414 280294 9482 280350
rect 9538 280294 9606 280350
rect 9662 280294 39954 280350
rect 40010 280294 40078 280350
rect 40134 280294 40202 280350
rect 40258 280294 40326 280350
rect 40382 280294 59878 280350
rect 59934 280294 60002 280350
rect 60058 280294 90598 280350
rect 90654 280294 90722 280350
rect 90778 280294 101394 280350
rect 101450 280294 101518 280350
rect 101574 280294 101642 280350
rect 101698 280294 101766 280350
rect 101822 280294 132114 280350
rect 132170 280294 132238 280350
rect 132294 280294 132362 280350
rect 132418 280294 132486 280350
rect 132542 280294 162834 280350
rect 162890 280294 162958 280350
rect 163014 280294 163082 280350
rect 163138 280294 163206 280350
rect 163262 280294 167078 280350
rect 167134 280294 167202 280350
rect 167258 280294 172902 280350
rect 172958 280294 173026 280350
rect 173082 280294 178726 280350
rect 178782 280294 178850 280350
rect 178906 280294 184550 280350
rect 184606 280294 184674 280350
rect 184730 280294 193554 280350
rect 193610 280294 193678 280350
rect 193734 280294 193802 280350
rect 193858 280294 193926 280350
rect 193982 280294 224274 280350
rect 224330 280294 224398 280350
rect 224454 280294 224522 280350
rect 224578 280294 224646 280350
rect 224702 280294 255878 280350
rect 255934 280294 256002 280350
rect 256058 280294 286598 280350
rect 286654 280294 286722 280350
rect 286778 280294 317318 280350
rect 317374 280294 317442 280350
rect 317498 280294 348038 280350
rect 348094 280294 348162 280350
rect 348218 280294 377874 280350
rect 377930 280294 377998 280350
rect 378054 280294 378122 280350
rect 378178 280294 378246 280350
rect 378302 280294 408594 280350
rect 408650 280294 408718 280350
rect 408774 280294 408842 280350
rect 408898 280294 408966 280350
rect 409022 280294 439314 280350
rect 439370 280294 439438 280350
rect 439494 280294 439562 280350
rect 439618 280294 439686 280350
rect 439742 280294 470034 280350
rect 470090 280294 470158 280350
rect 470214 280294 470282 280350
rect 470338 280294 470406 280350
rect 470462 280294 500754 280350
rect 500810 280294 500878 280350
rect 500934 280294 501002 280350
rect 501058 280294 501126 280350
rect 501182 280294 531474 280350
rect 531530 280294 531598 280350
rect 531654 280294 531722 280350
rect 531778 280294 531846 280350
rect 531902 280294 562194 280350
rect 562250 280294 562318 280350
rect 562374 280294 562442 280350
rect 562498 280294 562566 280350
rect 562622 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect -1916 280226 597980 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 9234 280226
rect 9290 280170 9358 280226
rect 9414 280170 9482 280226
rect 9538 280170 9606 280226
rect 9662 280170 39954 280226
rect 40010 280170 40078 280226
rect 40134 280170 40202 280226
rect 40258 280170 40326 280226
rect 40382 280170 59878 280226
rect 59934 280170 60002 280226
rect 60058 280170 90598 280226
rect 90654 280170 90722 280226
rect 90778 280170 101394 280226
rect 101450 280170 101518 280226
rect 101574 280170 101642 280226
rect 101698 280170 101766 280226
rect 101822 280170 132114 280226
rect 132170 280170 132238 280226
rect 132294 280170 132362 280226
rect 132418 280170 132486 280226
rect 132542 280170 162834 280226
rect 162890 280170 162958 280226
rect 163014 280170 163082 280226
rect 163138 280170 163206 280226
rect 163262 280170 167078 280226
rect 167134 280170 167202 280226
rect 167258 280170 172902 280226
rect 172958 280170 173026 280226
rect 173082 280170 178726 280226
rect 178782 280170 178850 280226
rect 178906 280170 184550 280226
rect 184606 280170 184674 280226
rect 184730 280170 193554 280226
rect 193610 280170 193678 280226
rect 193734 280170 193802 280226
rect 193858 280170 193926 280226
rect 193982 280170 224274 280226
rect 224330 280170 224398 280226
rect 224454 280170 224522 280226
rect 224578 280170 224646 280226
rect 224702 280170 255878 280226
rect 255934 280170 256002 280226
rect 256058 280170 286598 280226
rect 286654 280170 286722 280226
rect 286778 280170 317318 280226
rect 317374 280170 317442 280226
rect 317498 280170 348038 280226
rect 348094 280170 348162 280226
rect 348218 280170 377874 280226
rect 377930 280170 377998 280226
rect 378054 280170 378122 280226
rect 378178 280170 378246 280226
rect 378302 280170 408594 280226
rect 408650 280170 408718 280226
rect 408774 280170 408842 280226
rect 408898 280170 408966 280226
rect 409022 280170 439314 280226
rect 439370 280170 439438 280226
rect 439494 280170 439562 280226
rect 439618 280170 439686 280226
rect 439742 280170 470034 280226
rect 470090 280170 470158 280226
rect 470214 280170 470282 280226
rect 470338 280170 470406 280226
rect 470462 280170 500754 280226
rect 500810 280170 500878 280226
rect 500934 280170 501002 280226
rect 501058 280170 501126 280226
rect 501182 280170 531474 280226
rect 531530 280170 531598 280226
rect 531654 280170 531722 280226
rect 531778 280170 531846 280226
rect 531902 280170 562194 280226
rect 562250 280170 562318 280226
rect 562374 280170 562442 280226
rect 562498 280170 562566 280226
rect 562622 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect -1916 280102 597980 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 9234 280102
rect 9290 280046 9358 280102
rect 9414 280046 9482 280102
rect 9538 280046 9606 280102
rect 9662 280046 39954 280102
rect 40010 280046 40078 280102
rect 40134 280046 40202 280102
rect 40258 280046 40326 280102
rect 40382 280046 59878 280102
rect 59934 280046 60002 280102
rect 60058 280046 90598 280102
rect 90654 280046 90722 280102
rect 90778 280046 101394 280102
rect 101450 280046 101518 280102
rect 101574 280046 101642 280102
rect 101698 280046 101766 280102
rect 101822 280046 132114 280102
rect 132170 280046 132238 280102
rect 132294 280046 132362 280102
rect 132418 280046 132486 280102
rect 132542 280046 162834 280102
rect 162890 280046 162958 280102
rect 163014 280046 163082 280102
rect 163138 280046 163206 280102
rect 163262 280046 167078 280102
rect 167134 280046 167202 280102
rect 167258 280046 172902 280102
rect 172958 280046 173026 280102
rect 173082 280046 178726 280102
rect 178782 280046 178850 280102
rect 178906 280046 184550 280102
rect 184606 280046 184674 280102
rect 184730 280046 193554 280102
rect 193610 280046 193678 280102
rect 193734 280046 193802 280102
rect 193858 280046 193926 280102
rect 193982 280046 224274 280102
rect 224330 280046 224398 280102
rect 224454 280046 224522 280102
rect 224578 280046 224646 280102
rect 224702 280046 255878 280102
rect 255934 280046 256002 280102
rect 256058 280046 286598 280102
rect 286654 280046 286722 280102
rect 286778 280046 317318 280102
rect 317374 280046 317442 280102
rect 317498 280046 348038 280102
rect 348094 280046 348162 280102
rect 348218 280046 377874 280102
rect 377930 280046 377998 280102
rect 378054 280046 378122 280102
rect 378178 280046 378246 280102
rect 378302 280046 408594 280102
rect 408650 280046 408718 280102
rect 408774 280046 408842 280102
rect 408898 280046 408966 280102
rect 409022 280046 439314 280102
rect 439370 280046 439438 280102
rect 439494 280046 439562 280102
rect 439618 280046 439686 280102
rect 439742 280046 470034 280102
rect 470090 280046 470158 280102
rect 470214 280046 470282 280102
rect 470338 280046 470406 280102
rect 470462 280046 500754 280102
rect 500810 280046 500878 280102
rect 500934 280046 501002 280102
rect 501058 280046 501126 280102
rect 501182 280046 531474 280102
rect 531530 280046 531598 280102
rect 531654 280046 531722 280102
rect 531778 280046 531846 280102
rect 531902 280046 562194 280102
rect 562250 280046 562318 280102
rect 562374 280046 562442 280102
rect 562498 280046 562566 280102
rect 562622 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect -1916 279978 597980 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 9234 279978
rect 9290 279922 9358 279978
rect 9414 279922 9482 279978
rect 9538 279922 9606 279978
rect 9662 279922 39954 279978
rect 40010 279922 40078 279978
rect 40134 279922 40202 279978
rect 40258 279922 40326 279978
rect 40382 279922 59878 279978
rect 59934 279922 60002 279978
rect 60058 279922 90598 279978
rect 90654 279922 90722 279978
rect 90778 279922 101394 279978
rect 101450 279922 101518 279978
rect 101574 279922 101642 279978
rect 101698 279922 101766 279978
rect 101822 279922 132114 279978
rect 132170 279922 132238 279978
rect 132294 279922 132362 279978
rect 132418 279922 132486 279978
rect 132542 279922 162834 279978
rect 162890 279922 162958 279978
rect 163014 279922 163082 279978
rect 163138 279922 163206 279978
rect 163262 279922 167078 279978
rect 167134 279922 167202 279978
rect 167258 279922 172902 279978
rect 172958 279922 173026 279978
rect 173082 279922 178726 279978
rect 178782 279922 178850 279978
rect 178906 279922 184550 279978
rect 184606 279922 184674 279978
rect 184730 279922 193554 279978
rect 193610 279922 193678 279978
rect 193734 279922 193802 279978
rect 193858 279922 193926 279978
rect 193982 279922 224274 279978
rect 224330 279922 224398 279978
rect 224454 279922 224522 279978
rect 224578 279922 224646 279978
rect 224702 279922 255878 279978
rect 255934 279922 256002 279978
rect 256058 279922 286598 279978
rect 286654 279922 286722 279978
rect 286778 279922 317318 279978
rect 317374 279922 317442 279978
rect 317498 279922 348038 279978
rect 348094 279922 348162 279978
rect 348218 279922 377874 279978
rect 377930 279922 377998 279978
rect 378054 279922 378122 279978
rect 378178 279922 378246 279978
rect 378302 279922 408594 279978
rect 408650 279922 408718 279978
rect 408774 279922 408842 279978
rect 408898 279922 408966 279978
rect 409022 279922 439314 279978
rect 439370 279922 439438 279978
rect 439494 279922 439562 279978
rect 439618 279922 439686 279978
rect 439742 279922 470034 279978
rect 470090 279922 470158 279978
rect 470214 279922 470282 279978
rect 470338 279922 470406 279978
rect 470462 279922 500754 279978
rect 500810 279922 500878 279978
rect 500934 279922 501002 279978
rect 501058 279922 501126 279978
rect 501182 279922 531474 279978
rect 531530 279922 531598 279978
rect 531654 279922 531722 279978
rect 531778 279922 531846 279978
rect 531902 279922 562194 279978
rect 562250 279922 562318 279978
rect 562374 279922 562442 279978
rect 562498 279922 562566 279978
rect 562622 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect -1916 279826 597980 279922
rect -1916 274350 597980 274446
rect -1916 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 36234 274350
rect 36290 274294 36358 274350
rect 36414 274294 36482 274350
rect 36538 274294 36606 274350
rect 36662 274294 44518 274350
rect 44574 274294 44642 274350
rect 44698 274294 75238 274350
rect 75294 274294 75362 274350
rect 75418 274294 97674 274350
rect 97730 274294 97798 274350
rect 97854 274294 97922 274350
rect 97978 274294 98046 274350
rect 98102 274294 128394 274350
rect 128450 274294 128518 274350
rect 128574 274294 128642 274350
rect 128698 274294 128766 274350
rect 128822 274294 159114 274350
rect 159170 274294 159238 274350
rect 159294 274294 159362 274350
rect 159418 274294 159486 274350
rect 159542 274294 164166 274350
rect 164222 274294 164290 274350
rect 164346 274294 169990 274350
rect 170046 274294 170114 274350
rect 170170 274294 175814 274350
rect 175870 274294 175938 274350
rect 175994 274294 181638 274350
rect 181694 274294 181762 274350
rect 181818 274294 189834 274350
rect 189890 274294 189958 274350
rect 190014 274294 190082 274350
rect 190138 274294 190206 274350
rect 190262 274294 220554 274350
rect 220610 274294 220678 274350
rect 220734 274294 220802 274350
rect 220858 274294 220926 274350
rect 220982 274294 240518 274350
rect 240574 274294 240642 274350
rect 240698 274294 271238 274350
rect 271294 274294 271362 274350
rect 271418 274294 301958 274350
rect 302014 274294 302082 274350
rect 302138 274294 332678 274350
rect 332734 274294 332802 274350
rect 332858 274294 363398 274350
rect 363454 274294 363522 274350
rect 363578 274294 404874 274350
rect 404930 274294 404998 274350
rect 405054 274294 405122 274350
rect 405178 274294 405246 274350
rect 405302 274294 435594 274350
rect 435650 274294 435718 274350
rect 435774 274294 435842 274350
rect 435898 274294 435966 274350
rect 436022 274294 466314 274350
rect 466370 274294 466438 274350
rect 466494 274294 466562 274350
rect 466618 274294 466686 274350
rect 466742 274294 497034 274350
rect 497090 274294 497158 274350
rect 497214 274294 497282 274350
rect 497338 274294 497406 274350
rect 497462 274294 527754 274350
rect 527810 274294 527878 274350
rect 527934 274294 528002 274350
rect 528058 274294 528126 274350
rect 528182 274294 558474 274350
rect 558530 274294 558598 274350
rect 558654 274294 558722 274350
rect 558778 274294 558846 274350
rect 558902 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597980 274350
rect -1916 274226 597980 274294
rect -1916 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 36234 274226
rect 36290 274170 36358 274226
rect 36414 274170 36482 274226
rect 36538 274170 36606 274226
rect 36662 274170 44518 274226
rect 44574 274170 44642 274226
rect 44698 274170 75238 274226
rect 75294 274170 75362 274226
rect 75418 274170 97674 274226
rect 97730 274170 97798 274226
rect 97854 274170 97922 274226
rect 97978 274170 98046 274226
rect 98102 274170 128394 274226
rect 128450 274170 128518 274226
rect 128574 274170 128642 274226
rect 128698 274170 128766 274226
rect 128822 274170 159114 274226
rect 159170 274170 159238 274226
rect 159294 274170 159362 274226
rect 159418 274170 159486 274226
rect 159542 274170 164166 274226
rect 164222 274170 164290 274226
rect 164346 274170 169990 274226
rect 170046 274170 170114 274226
rect 170170 274170 175814 274226
rect 175870 274170 175938 274226
rect 175994 274170 181638 274226
rect 181694 274170 181762 274226
rect 181818 274170 189834 274226
rect 189890 274170 189958 274226
rect 190014 274170 190082 274226
rect 190138 274170 190206 274226
rect 190262 274170 220554 274226
rect 220610 274170 220678 274226
rect 220734 274170 220802 274226
rect 220858 274170 220926 274226
rect 220982 274170 240518 274226
rect 240574 274170 240642 274226
rect 240698 274170 271238 274226
rect 271294 274170 271362 274226
rect 271418 274170 301958 274226
rect 302014 274170 302082 274226
rect 302138 274170 332678 274226
rect 332734 274170 332802 274226
rect 332858 274170 363398 274226
rect 363454 274170 363522 274226
rect 363578 274170 404874 274226
rect 404930 274170 404998 274226
rect 405054 274170 405122 274226
rect 405178 274170 405246 274226
rect 405302 274170 435594 274226
rect 435650 274170 435718 274226
rect 435774 274170 435842 274226
rect 435898 274170 435966 274226
rect 436022 274170 466314 274226
rect 466370 274170 466438 274226
rect 466494 274170 466562 274226
rect 466618 274170 466686 274226
rect 466742 274170 497034 274226
rect 497090 274170 497158 274226
rect 497214 274170 497282 274226
rect 497338 274170 497406 274226
rect 497462 274170 527754 274226
rect 527810 274170 527878 274226
rect 527934 274170 528002 274226
rect 528058 274170 528126 274226
rect 528182 274170 558474 274226
rect 558530 274170 558598 274226
rect 558654 274170 558722 274226
rect 558778 274170 558846 274226
rect 558902 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597980 274226
rect -1916 274102 597980 274170
rect -1916 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 36234 274102
rect 36290 274046 36358 274102
rect 36414 274046 36482 274102
rect 36538 274046 36606 274102
rect 36662 274046 44518 274102
rect 44574 274046 44642 274102
rect 44698 274046 75238 274102
rect 75294 274046 75362 274102
rect 75418 274046 97674 274102
rect 97730 274046 97798 274102
rect 97854 274046 97922 274102
rect 97978 274046 98046 274102
rect 98102 274046 128394 274102
rect 128450 274046 128518 274102
rect 128574 274046 128642 274102
rect 128698 274046 128766 274102
rect 128822 274046 159114 274102
rect 159170 274046 159238 274102
rect 159294 274046 159362 274102
rect 159418 274046 159486 274102
rect 159542 274046 164166 274102
rect 164222 274046 164290 274102
rect 164346 274046 169990 274102
rect 170046 274046 170114 274102
rect 170170 274046 175814 274102
rect 175870 274046 175938 274102
rect 175994 274046 181638 274102
rect 181694 274046 181762 274102
rect 181818 274046 189834 274102
rect 189890 274046 189958 274102
rect 190014 274046 190082 274102
rect 190138 274046 190206 274102
rect 190262 274046 220554 274102
rect 220610 274046 220678 274102
rect 220734 274046 220802 274102
rect 220858 274046 220926 274102
rect 220982 274046 240518 274102
rect 240574 274046 240642 274102
rect 240698 274046 271238 274102
rect 271294 274046 271362 274102
rect 271418 274046 301958 274102
rect 302014 274046 302082 274102
rect 302138 274046 332678 274102
rect 332734 274046 332802 274102
rect 332858 274046 363398 274102
rect 363454 274046 363522 274102
rect 363578 274046 404874 274102
rect 404930 274046 404998 274102
rect 405054 274046 405122 274102
rect 405178 274046 405246 274102
rect 405302 274046 435594 274102
rect 435650 274046 435718 274102
rect 435774 274046 435842 274102
rect 435898 274046 435966 274102
rect 436022 274046 466314 274102
rect 466370 274046 466438 274102
rect 466494 274046 466562 274102
rect 466618 274046 466686 274102
rect 466742 274046 497034 274102
rect 497090 274046 497158 274102
rect 497214 274046 497282 274102
rect 497338 274046 497406 274102
rect 497462 274046 527754 274102
rect 527810 274046 527878 274102
rect 527934 274046 528002 274102
rect 528058 274046 528126 274102
rect 528182 274046 558474 274102
rect 558530 274046 558598 274102
rect 558654 274046 558722 274102
rect 558778 274046 558846 274102
rect 558902 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597980 274102
rect -1916 273978 597980 274046
rect -1916 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 36234 273978
rect 36290 273922 36358 273978
rect 36414 273922 36482 273978
rect 36538 273922 36606 273978
rect 36662 273922 44518 273978
rect 44574 273922 44642 273978
rect 44698 273922 75238 273978
rect 75294 273922 75362 273978
rect 75418 273922 97674 273978
rect 97730 273922 97798 273978
rect 97854 273922 97922 273978
rect 97978 273922 98046 273978
rect 98102 273922 128394 273978
rect 128450 273922 128518 273978
rect 128574 273922 128642 273978
rect 128698 273922 128766 273978
rect 128822 273922 159114 273978
rect 159170 273922 159238 273978
rect 159294 273922 159362 273978
rect 159418 273922 159486 273978
rect 159542 273922 164166 273978
rect 164222 273922 164290 273978
rect 164346 273922 169990 273978
rect 170046 273922 170114 273978
rect 170170 273922 175814 273978
rect 175870 273922 175938 273978
rect 175994 273922 181638 273978
rect 181694 273922 181762 273978
rect 181818 273922 189834 273978
rect 189890 273922 189958 273978
rect 190014 273922 190082 273978
rect 190138 273922 190206 273978
rect 190262 273922 220554 273978
rect 220610 273922 220678 273978
rect 220734 273922 220802 273978
rect 220858 273922 220926 273978
rect 220982 273922 240518 273978
rect 240574 273922 240642 273978
rect 240698 273922 271238 273978
rect 271294 273922 271362 273978
rect 271418 273922 301958 273978
rect 302014 273922 302082 273978
rect 302138 273922 332678 273978
rect 332734 273922 332802 273978
rect 332858 273922 363398 273978
rect 363454 273922 363522 273978
rect 363578 273922 404874 273978
rect 404930 273922 404998 273978
rect 405054 273922 405122 273978
rect 405178 273922 405246 273978
rect 405302 273922 435594 273978
rect 435650 273922 435718 273978
rect 435774 273922 435842 273978
rect 435898 273922 435966 273978
rect 436022 273922 466314 273978
rect 466370 273922 466438 273978
rect 466494 273922 466562 273978
rect 466618 273922 466686 273978
rect 466742 273922 497034 273978
rect 497090 273922 497158 273978
rect 497214 273922 497282 273978
rect 497338 273922 497406 273978
rect 497462 273922 527754 273978
rect 527810 273922 527878 273978
rect 527934 273922 528002 273978
rect 528058 273922 528126 273978
rect 528182 273922 558474 273978
rect 558530 273922 558598 273978
rect 558654 273922 558722 273978
rect 558778 273922 558846 273978
rect 558902 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597980 273978
rect -1916 273826 597980 273922
rect 189516 268858 237652 268874
rect 189516 268802 189532 268858
rect 189588 268802 237580 268858
rect 237636 268802 237652 268858
rect 189516 268786 237652 268802
rect -1916 262350 597980 262446
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 9234 262350
rect 9290 262294 9358 262350
rect 9414 262294 9482 262350
rect 9538 262294 9606 262350
rect 9662 262294 39954 262350
rect 40010 262294 40078 262350
rect 40134 262294 40202 262350
rect 40258 262294 40326 262350
rect 40382 262294 59878 262350
rect 59934 262294 60002 262350
rect 60058 262294 90598 262350
rect 90654 262294 90722 262350
rect 90778 262294 101394 262350
rect 101450 262294 101518 262350
rect 101574 262294 101642 262350
rect 101698 262294 101766 262350
rect 101822 262294 132114 262350
rect 132170 262294 132238 262350
rect 132294 262294 132362 262350
rect 132418 262294 132486 262350
rect 132542 262294 162834 262350
rect 162890 262294 162958 262350
rect 163014 262294 163082 262350
rect 163138 262294 163206 262350
rect 163262 262294 193554 262350
rect 193610 262294 193678 262350
rect 193734 262294 193802 262350
rect 193858 262294 193926 262350
rect 193982 262294 224274 262350
rect 224330 262294 224398 262350
rect 224454 262294 224522 262350
rect 224578 262294 224646 262350
rect 224702 262294 255878 262350
rect 255934 262294 256002 262350
rect 256058 262294 286598 262350
rect 286654 262294 286722 262350
rect 286778 262294 317318 262350
rect 317374 262294 317442 262350
rect 317498 262294 348038 262350
rect 348094 262294 348162 262350
rect 348218 262294 377874 262350
rect 377930 262294 377998 262350
rect 378054 262294 378122 262350
rect 378178 262294 378246 262350
rect 378302 262294 408594 262350
rect 408650 262294 408718 262350
rect 408774 262294 408842 262350
rect 408898 262294 408966 262350
rect 409022 262294 439314 262350
rect 439370 262294 439438 262350
rect 439494 262294 439562 262350
rect 439618 262294 439686 262350
rect 439742 262294 470034 262350
rect 470090 262294 470158 262350
rect 470214 262294 470282 262350
rect 470338 262294 470406 262350
rect 470462 262294 500754 262350
rect 500810 262294 500878 262350
rect 500934 262294 501002 262350
rect 501058 262294 501126 262350
rect 501182 262294 531474 262350
rect 531530 262294 531598 262350
rect 531654 262294 531722 262350
rect 531778 262294 531846 262350
rect 531902 262294 562194 262350
rect 562250 262294 562318 262350
rect 562374 262294 562442 262350
rect 562498 262294 562566 262350
rect 562622 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect -1916 262226 597980 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 9234 262226
rect 9290 262170 9358 262226
rect 9414 262170 9482 262226
rect 9538 262170 9606 262226
rect 9662 262170 39954 262226
rect 40010 262170 40078 262226
rect 40134 262170 40202 262226
rect 40258 262170 40326 262226
rect 40382 262170 59878 262226
rect 59934 262170 60002 262226
rect 60058 262170 90598 262226
rect 90654 262170 90722 262226
rect 90778 262170 101394 262226
rect 101450 262170 101518 262226
rect 101574 262170 101642 262226
rect 101698 262170 101766 262226
rect 101822 262170 132114 262226
rect 132170 262170 132238 262226
rect 132294 262170 132362 262226
rect 132418 262170 132486 262226
rect 132542 262170 162834 262226
rect 162890 262170 162958 262226
rect 163014 262170 163082 262226
rect 163138 262170 163206 262226
rect 163262 262170 193554 262226
rect 193610 262170 193678 262226
rect 193734 262170 193802 262226
rect 193858 262170 193926 262226
rect 193982 262170 224274 262226
rect 224330 262170 224398 262226
rect 224454 262170 224522 262226
rect 224578 262170 224646 262226
rect 224702 262170 255878 262226
rect 255934 262170 256002 262226
rect 256058 262170 286598 262226
rect 286654 262170 286722 262226
rect 286778 262170 317318 262226
rect 317374 262170 317442 262226
rect 317498 262170 348038 262226
rect 348094 262170 348162 262226
rect 348218 262170 377874 262226
rect 377930 262170 377998 262226
rect 378054 262170 378122 262226
rect 378178 262170 378246 262226
rect 378302 262170 408594 262226
rect 408650 262170 408718 262226
rect 408774 262170 408842 262226
rect 408898 262170 408966 262226
rect 409022 262170 439314 262226
rect 439370 262170 439438 262226
rect 439494 262170 439562 262226
rect 439618 262170 439686 262226
rect 439742 262170 470034 262226
rect 470090 262170 470158 262226
rect 470214 262170 470282 262226
rect 470338 262170 470406 262226
rect 470462 262170 500754 262226
rect 500810 262170 500878 262226
rect 500934 262170 501002 262226
rect 501058 262170 501126 262226
rect 501182 262170 531474 262226
rect 531530 262170 531598 262226
rect 531654 262170 531722 262226
rect 531778 262170 531846 262226
rect 531902 262170 562194 262226
rect 562250 262170 562318 262226
rect 562374 262170 562442 262226
rect 562498 262170 562566 262226
rect 562622 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect -1916 262102 597980 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 9234 262102
rect 9290 262046 9358 262102
rect 9414 262046 9482 262102
rect 9538 262046 9606 262102
rect 9662 262046 39954 262102
rect 40010 262046 40078 262102
rect 40134 262046 40202 262102
rect 40258 262046 40326 262102
rect 40382 262046 59878 262102
rect 59934 262046 60002 262102
rect 60058 262046 90598 262102
rect 90654 262046 90722 262102
rect 90778 262046 101394 262102
rect 101450 262046 101518 262102
rect 101574 262046 101642 262102
rect 101698 262046 101766 262102
rect 101822 262046 132114 262102
rect 132170 262046 132238 262102
rect 132294 262046 132362 262102
rect 132418 262046 132486 262102
rect 132542 262046 162834 262102
rect 162890 262046 162958 262102
rect 163014 262046 163082 262102
rect 163138 262046 163206 262102
rect 163262 262046 193554 262102
rect 193610 262046 193678 262102
rect 193734 262046 193802 262102
rect 193858 262046 193926 262102
rect 193982 262046 224274 262102
rect 224330 262046 224398 262102
rect 224454 262046 224522 262102
rect 224578 262046 224646 262102
rect 224702 262046 255878 262102
rect 255934 262046 256002 262102
rect 256058 262046 286598 262102
rect 286654 262046 286722 262102
rect 286778 262046 317318 262102
rect 317374 262046 317442 262102
rect 317498 262046 348038 262102
rect 348094 262046 348162 262102
rect 348218 262046 377874 262102
rect 377930 262046 377998 262102
rect 378054 262046 378122 262102
rect 378178 262046 378246 262102
rect 378302 262046 408594 262102
rect 408650 262046 408718 262102
rect 408774 262046 408842 262102
rect 408898 262046 408966 262102
rect 409022 262046 439314 262102
rect 439370 262046 439438 262102
rect 439494 262046 439562 262102
rect 439618 262046 439686 262102
rect 439742 262046 470034 262102
rect 470090 262046 470158 262102
rect 470214 262046 470282 262102
rect 470338 262046 470406 262102
rect 470462 262046 500754 262102
rect 500810 262046 500878 262102
rect 500934 262046 501002 262102
rect 501058 262046 501126 262102
rect 501182 262046 531474 262102
rect 531530 262046 531598 262102
rect 531654 262046 531722 262102
rect 531778 262046 531846 262102
rect 531902 262046 562194 262102
rect 562250 262046 562318 262102
rect 562374 262046 562442 262102
rect 562498 262046 562566 262102
rect 562622 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect -1916 261978 597980 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 9234 261978
rect 9290 261922 9358 261978
rect 9414 261922 9482 261978
rect 9538 261922 9606 261978
rect 9662 261922 39954 261978
rect 40010 261922 40078 261978
rect 40134 261922 40202 261978
rect 40258 261922 40326 261978
rect 40382 261922 59878 261978
rect 59934 261922 60002 261978
rect 60058 261922 90598 261978
rect 90654 261922 90722 261978
rect 90778 261922 101394 261978
rect 101450 261922 101518 261978
rect 101574 261922 101642 261978
rect 101698 261922 101766 261978
rect 101822 261922 132114 261978
rect 132170 261922 132238 261978
rect 132294 261922 132362 261978
rect 132418 261922 132486 261978
rect 132542 261922 162834 261978
rect 162890 261922 162958 261978
rect 163014 261922 163082 261978
rect 163138 261922 163206 261978
rect 163262 261922 193554 261978
rect 193610 261922 193678 261978
rect 193734 261922 193802 261978
rect 193858 261922 193926 261978
rect 193982 261922 224274 261978
rect 224330 261922 224398 261978
rect 224454 261922 224522 261978
rect 224578 261922 224646 261978
rect 224702 261922 255878 261978
rect 255934 261922 256002 261978
rect 256058 261922 286598 261978
rect 286654 261922 286722 261978
rect 286778 261922 317318 261978
rect 317374 261922 317442 261978
rect 317498 261922 348038 261978
rect 348094 261922 348162 261978
rect 348218 261922 377874 261978
rect 377930 261922 377998 261978
rect 378054 261922 378122 261978
rect 378178 261922 378246 261978
rect 378302 261922 408594 261978
rect 408650 261922 408718 261978
rect 408774 261922 408842 261978
rect 408898 261922 408966 261978
rect 409022 261922 439314 261978
rect 439370 261922 439438 261978
rect 439494 261922 439562 261978
rect 439618 261922 439686 261978
rect 439742 261922 470034 261978
rect 470090 261922 470158 261978
rect 470214 261922 470282 261978
rect 470338 261922 470406 261978
rect 470462 261922 500754 261978
rect 500810 261922 500878 261978
rect 500934 261922 501002 261978
rect 501058 261922 501126 261978
rect 501182 261922 531474 261978
rect 531530 261922 531598 261978
rect 531654 261922 531722 261978
rect 531778 261922 531846 261978
rect 531902 261922 562194 261978
rect 562250 261922 562318 261978
rect 562374 261922 562442 261978
rect 562498 261922 562566 261978
rect 562622 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect -1916 261826 597980 261922
rect 358636 257878 375300 257894
rect 358636 257822 358652 257878
rect 358708 257822 375228 257878
rect 375284 257822 375300 257878
rect 358636 257806 375300 257822
rect -1916 256350 597980 256446
rect -1916 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 36234 256350
rect 36290 256294 36358 256350
rect 36414 256294 36482 256350
rect 36538 256294 36606 256350
rect 36662 256294 44518 256350
rect 44574 256294 44642 256350
rect 44698 256294 75238 256350
rect 75294 256294 75362 256350
rect 75418 256294 97674 256350
rect 97730 256294 97798 256350
rect 97854 256294 97922 256350
rect 97978 256294 98046 256350
rect 98102 256294 128394 256350
rect 128450 256294 128518 256350
rect 128574 256294 128642 256350
rect 128698 256294 128766 256350
rect 128822 256294 159114 256350
rect 159170 256294 159238 256350
rect 159294 256294 159362 256350
rect 159418 256294 159486 256350
rect 159542 256294 189834 256350
rect 189890 256294 189958 256350
rect 190014 256294 190082 256350
rect 190138 256294 190206 256350
rect 190262 256294 220554 256350
rect 220610 256294 220678 256350
rect 220734 256294 220802 256350
rect 220858 256294 220926 256350
rect 220982 256294 251274 256350
rect 251330 256294 251398 256350
rect 251454 256294 251522 256350
rect 251578 256294 251646 256350
rect 251702 256294 281994 256350
rect 282050 256294 282118 256350
rect 282174 256294 282242 256350
rect 282298 256294 282366 256350
rect 282422 256294 312714 256350
rect 312770 256294 312838 256350
rect 312894 256294 312962 256350
rect 313018 256294 313086 256350
rect 313142 256294 343434 256350
rect 343490 256294 343558 256350
rect 343614 256294 343682 256350
rect 343738 256294 343806 256350
rect 343862 256294 374154 256350
rect 374210 256294 374278 256350
rect 374334 256294 374402 256350
rect 374458 256294 374526 256350
rect 374582 256294 404874 256350
rect 404930 256294 404998 256350
rect 405054 256294 405122 256350
rect 405178 256294 405246 256350
rect 405302 256294 435594 256350
rect 435650 256294 435718 256350
rect 435774 256294 435842 256350
rect 435898 256294 435966 256350
rect 436022 256294 466314 256350
rect 466370 256294 466438 256350
rect 466494 256294 466562 256350
rect 466618 256294 466686 256350
rect 466742 256294 497034 256350
rect 497090 256294 497158 256350
rect 497214 256294 497282 256350
rect 497338 256294 497406 256350
rect 497462 256294 527754 256350
rect 527810 256294 527878 256350
rect 527934 256294 528002 256350
rect 528058 256294 528126 256350
rect 528182 256294 558474 256350
rect 558530 256294 558598 256350
rect 558654 256294 558722 256350
rect 558778 256294 558846 256350
rect 558902 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597980 256350
rect -1916 256226 597980 256294
rect -1916 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 36234 256226
rect 36290 256170 36358 256226
rect 36414 256170 36482 256226
rect 36538 256170 36606 256226
rect 36662 256170 44518 256226
rect 44574 256170 44642 256226
rect 44698 256170 75238 256226
rect 75294 256170 75362 256226
rect 75418 256170 97674 256226
rect 97730 256170 97798 256226
rect 97854 256170 97922 256226
rect 97978 256170 98046 256226
rect 98102 256170 128394 256226
rect 128450 256170 128518 256226
rect 128574 256170 128642 256226
rect 128698 256170 128766 256226
rect 128822 256170 159114 256226
rect 159170 256170 159238 256226
rect 159294 256170 159362 256226
rect 159418 256170 159486 256226
rect 159542 256170 189834 256226
rect 189890 256170 189958 256226
rect 190014 256170 190082 256226
rect 190138 256170 190206 256226
rect 190262 256170 220554 256226
rect 220610 256170 220678 256226
rect 220734 256170 220802 256226
rect 220858 256170 220926 256226
rect 220982 256170 251274 256226
rect 251330 256170 251398 256226
rect 251454 256170 251522 256226
rect 251578 256170 251646 256226
rect 251702 256170 281994 256226
rect 282050 256170 282118 256226
rect 282174 256170 282242 256226
rect 282298 256170 282366 256226
rect 282422 256170 312714 256226
rect 312770 256170 312838 256226
rect 312894 256170 312962 256226
rect 313018 256170 313086 256226
rect 313142 256170 343434 256226
rect 343490 256170 343558 256226
rect 343614 256170 343682 256226
rect 343738 256170 343806 256226
rect 343862 256170 374154 256226
rect 374210 256170 374278 256226
rect 374334 256170 374402 256226
rect 374458 256170 374526 256226
rect 374582 256170 404874 256226
rect 404930 256170 404998 256226
rect 405054 256170 405122 256226
rect 405178 256170 405246 256226
rect 405302 256170 435594 256226
rect 435650 256170 435718 256226
rect 435774 256170 435842 256226
rect 435898 256170 435966 256226
rect 436022 256170 466314 256226
rect 466370 256170 466438 256226
rect 466494 256170 466562 256226
rect 466618 256170 466686 256226
rect 466742 256170 497034 256226
rect 497090 256170 497158 256226
rect 497214 256170 497282 256226
rect 497338 256170 497406 256226
rect 497462 256170 527754 256226
rect 527810 256170 527878 256226
rect 527934 256170 528002 256226
rect 528058 256170 528126 256226
rect 528182 256170 558474 256226
rect 558530 256170 558598 256226
rect 558654 256170 558722 256226
rect 558778 256170 558846 256226
rect 558902 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597980 256226
rect -1916 256102 597980 256170
rect -1916 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 36234 256102
rect 36290 256046 36358 256102
rect 36414 256046 36482 256102
rect 36538 256046 36606 256102
rect 36662 256046 44518 256102
rect 44574 256046 44642 256102
rect 44698 256046 75238 256102
rect 75294 256046 75362 256102
rect 75418 256046 97674 256102
rect 97730 256046 97798 256102
rect 97854 256046 97922 256102
rect 97978 256046 98046 256102
rect 98102 256046 128394 256102
rect 128450 256046 128518 256102
rect 128574 256046 128642 256102
rect 128698 256046 128766 256102
rect 128822 256046 159114 256102
rect 159170 256046 159238 256102
rect 159294 256046 159362 256102
rect 159418 256046 159486 256102
rect 159542 256046 189834 256102
rect 189890 256046 189958 256102
rect 190014 256046 190082 256102
rect 190138 256046 190206 256102
rect 190262 256046 220554 256102
rect 220610 256046 220678 256102
rect 220734 256046 220802 256102
rect 220858 256046 220926 256102
rect 220982 256046 251274 256102
rect 251330 256046 251398 256102
rect 251454 256046 251522 256102
rect 251578 256046 251646 256102
rect 251702 256046 281994 256102
rect 282050 256046 282118 256102
rect 282174 256046 282242 256102
rect 282298 256046 282366 256102
rect 282422 256046 312714 256102
rect 312770 256046 312838 256102
rect 312894 256046 312962 256102
rect 313018 256046 313086 256102
rect 313142 256046 343434 256102
rect 343490 256046 343558 256102
rect 343614 256046 343682 256102
rect 343738 256046 343806 256102
rect 343862 256046 374154 256102
rect 374210 256046 374278 256102
rect 374334 256046 374402 256102
rect 374458 256046 374526 256102
rect 374582 256046 404874 256102
rect 404930 256046 404998 256102
rect 405054 256046 405122 256102
rect 405178 256046 405246 256102
rect 405302 256046 435594 256102
rect 435650 256046 435718 256102
rect 435774 256046 435842 256102
rect 435898 256046 435966 256102
rect 436022 256046 466314 256102
rect 466370 256046 466438 256102
rect 466494 256046 466562 256102
rect 466618 256046 466686 256102
rect 466742 256046 497034 256102
rect 497090 256046 497158 256102
rect 497214 256046 497282 256102
rect 497338 256046 497406 256102
rect 497462 256046 527754 256102
rect 527810 256046 527878 256102
rect 527934 256046 528002 256102
rect 528058 256046 528126 256102
rect 528182 256046 558474 256102
rect 558530 256046 558598 256102
rect 558654 256046 558722 256102
rect 558778 256046 558846 256102
rect 558902 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597980 256102
rect -1916 255978 597980 256046
rect -1916 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 36234 255978
rect 36290 255922 36358 255978
rect 36414 255922 36482 255978
rect 36538 255922 36606 255978
rect 36662 255922 44518 255978
rect 44574 255922 44642 255978
rect 44698 255922 75238 255978
rect 75294 255922 75362 255978
rect 75418 255922 97674 255978
rect 97730 255922 97798 255978
rect 97854 255922 97922 255978
rect 97978 255922 98046 255978
rect 98102 255922 128394 255978
rect 128450 255922 128518 255978
rect 128574 255922 128642 255978
rect 128698 255922 128766 255978
rect 128822 255922 159114 255978
rect 159170 255922 159238 255978
rect 159294 255922 159362 255978
rect 159418 255922 159486 255978
rect 159542 255922 189834 255978
rect 189890 255922 189958 255978
rect 190014 255922 190082 255978
rect 190138 255922 190206 255978
rect 190262 255922 220554 255978
rect 220610 255922 220678 255978
rect 220734 255922 220802 255978
rect 220858 255922 220926 255978
rect 220982 255922 251274 255978
rect 251330 255922 251398 255978
rect 251454 255922 251522 255978
rect 251578 255922 251646 255978
rect 251702 255922 281994 255978
rect 282050 255922 282118 255978
rect 282174 255922 282242 255978
rect 282298 255922 282366 255978
rect 282422 255922 312714 255978
rect 312770 255922 312838 255978
rect 312894 255922 312962 255978
rect 313018 255922 313086 255978
rect 313142 255922 343434 255978
rect 343490 255922 343558 255978
rect 343614 255922 343682 255978
rect 343738 255922 343806 255978
rect 343862 255922 374154 255978
rect 374210 255922 374278 255978
rect 374334 255922 374402 255978
rect 374458 255922 374526 255978
rect 374582 255922 404874 255978
rect 404930 255922 404998 255978
rect 405054 255922 405122 255978
rect 405178 255922 405246 255978
rect 405302 255922 435594 255978
rect 435650 255922 435718 255978
rect 435774 255922 435842 255978
rect 435898 255922 435966 255978
rect 436022 255922 466314 255978
rect 466370 255922 466438 255978
rect 466494 255922 466562 255978
rect 466618 255922 466686 255978
rect 466742 255922 497034 255978
rect 497090 255922 497158 255978
rect 497214 255922 497282 255978
rect 497338 255922 497406 255978
rect 497462 255922 527754 255978
rect 527810 255922 527878 255978
rect 527934 255922 528002 255978
rect 528058 255922 528126 255978
rect 528182 255922 558474 255978
rect 558530 255922 558598 255978
rect 558654 255922 558722 255978
rect 558778 255922 558846 255978
rect 558902 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597980 255978
rect -1916 255826 597980 255922
rect 358748 253198 373956 253214
rect 358748 253142 358764 253198
rect 358820 253142 373884 253198
rect 373940 253142 373956 253198
rect 358748 253126 373956 253142
rect 358972 253018 375748 253034
rect 358972 252962 358988 253018
rect 359044 252962 375676 253018
rect 375732 252962 375748 253018
rect 358972 252946 375748 252962
rect 251900 252838 270580 252854
rect 251900 252782 251916 252838
rect 251972 252782 270508 252838
rect 270564 252782 270580 252838
rect 251900 252766 270580 252782
rect 359196 252838 376532 252854
rect 359196 252782 359212 252838
rect 359268 252782 376460 252838
rect 376516 252782 376532 252838
rect 359196 252766 376532 252782
rect 258844 252658 275620 252674
rect 258844 252602 258860 252658
rect 258916 252602 275548 252658
rect 275604 252602 275620 252658
rect 258844 252586 275620 252602
rect 252572 252478 269684 252494
rect 252572 252422 252588 252478
rect 252644 252422 269612 252478
rect 269668 252422 269684 252478
rect 252572 252406 269684 252422
rect 259740 252298 275732 252314
rect 259740 252242 259756 252298
rect 259812 252242 275660 252298
rect 275716 252242 275732 252298
rect 259740 252226 275732 252242
rect 260636 252118 269572 252134
rect 260636 252062 260652 252118
rect 260708 252062 269500 252118
rect 269556 252062 269572 252118
rect 260636 252046 269572 252062
rect 230956 249418 274724 249434
rect 230956 249362 230972 249418
rect 231028 249362 274652 249418
rect 274708 249362 274724 249418
rect 230956 249346 274724 249362
rect 4044 247078 46244 247094
rect 4044 247022 4060 247078
rect 4116 247022 46172 247078
rect 46228 247022 46244 247078
rect 4044 247006 46244 247022
rect 231852 246178 268788 246194
rect 231852 246122 231868 246178
rect 231924 246122 268716 246178
rect 268772 246122 268788 246178
rect 231852 246106 268788 246122
rect -1916 244350 597980 244446
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 9234 244350
rect 9290 244294 9358 244350
rect 9414 244294 9482 244350
rect 9538 244294 9606 244350
rect 9662 244294 39954 244350
rect 40010 244294 40078 244350
rect 40134 244294 40202 244350
rect 40258 244294 40326 244350
rect 40382 244294 59878 244350
rect 59934 244294 60002 244350
rect 60058 244294 70674 244350
rect 70730 244294 70798 244350
rect 70854 244294 70922 244350
rect 70978 244294 71046 244350
rect 71102 244294 90598 244350
rect 90654 244294 90722 244350
rect 90778 244294 101394 244350
rect 101450 244294 101518 244350
rect 101574 244294 101642 244350
rect 101698 244294 101766 244350
rect 101822 244294 132114 244350
rect 132170 244294 132238 244350
rect 132294 244294 132362 244350
rect 132418 244294 132486 244350
rect 132542 244294 162834 244350
rect 162890 244294 162958 244350
rect 163014 244294 163082 244350
rect 163138 244294 163206 244350
rect 163262 244294 193554 244350
rect 193610 244294 193678 244350
rect 193734 244294 193802 244350
rect 193858 244294 193926 244350
rect 193982 244294 224274 244350
rect 224330 244294 224398 244350
rect 224454 244294 224522 244350
rect 224578 244294 224646 244350
rect 224702 244294 254994 244350
rect 255050 244294 255118 244350
rect 255174 244294 255242 244350
rect 255298 244294 255366 244350
rect 255422 244294 285714 244350
rect 285770 244294 285838 244350
rect 285894 244294 285962 244350
rect 286018 244294 286086 244350
rect 286142 244294 316434 244350
rect 316490 244294 316558 244350
rect 316614 244294 316682 244350
rect 316738 244294 316806 244350
rect 316862 244294 347154 244350
rect 347210 244294 347278 244350
rect 347334 244294 347402 244350
rect 347458 244294 347526 244350
rect 347582 244294 377874 244350
rect 377930 244294 377998 244350
rect 378054 244294 378122 244350
rect 378178 244294 378246 244350
rect 378302 244294 408594 244350
rect 408650 244294 408718 244350
rect 408774 244294 408842 244350
rect 408898 244294 408966 244350
rect 409022 244294 439314 244350
rect 439370 244294 439438 244350
rect 439494 244294 439562 244350
rect 439618 244294 439686 244350
rect 439742 244294 470034 244350
rect 470090 244294 470158 244350
rect 470214 244294 470282 244350
rect 470338 244294 470406 244350
rect 470462 244294 500754 244350
rect 500810 244294 500878 244350
rect 500934 244294 501002 244350
rect 501058 244294 501126 244350
rect 501182 244294 531474 244350
rect 531530 244294 531598 244350
rect 531654 244294 531722 244350
rect 531778 244294 531846 244350
rect 531902 244294 562194 244350
rect 562250 244294 562318 244350
rect 562374 244294 562442 244350
rect 562498 244294 562566 244350
rect 562622 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect -1916 244226 597980 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 9234 244226
rect 9290 244170 9358 244226
rect 9414 244170 9482 244226
rect 9538 244170 9606 244226
rect 9662 244170 39954 244226
rect 40010 244170 40078 244226
rect 40134 244170 40202 244226
rect 40258 244170 40326 244226
rect 40382 244170 59878 244226
rect 59934 244170 60002 244226
rect 60058 244170 70674 244226
rect 70730 244170 70798 244226
rect 70854 244170 70922 244226
rect 70978 244170 71046 244226
rect 71102 244170 90598 244226
rect 90654 244170 90722 244226
rect 90778 244170 101394 244226
rect 101450 244170 101518 244226
rect 101574 244170 101642 244226
rect 101698 244170 101766 244226
rect 101822 244170 132114 244226
rect 132170 244170 132238 244226
rect 132294 244170 132362 244226
rect 132418 244170 132486 244226
rect 132542 244170 162834 244226
rect 162890 244170 162958 244226
rect 163014 244170 163082 244226
rect 163138 244170 163206 244226
rect 163262 244170 193554 244226
rect 193610 244170 193678 244226
rect 193734 244170 193802 244226
rect 193858 244170 193926 244226
rect 193982 244170 224274 244226
rect 224330 244170 224398 244226
rect 224454 244170 224522 244226
rect 224578 244170 224646 244226
rect 224702 244170 254994 244226
rect 255050 244170 255118 244226
rect 255174 244170 255242 244226
rect 255298 244170 255366 244226
rect 255422 244170 285714 244226
rect 285770 244170 285838 244226
rect 285894 244170 285962 244226
rect 286018 244170 286086 244226
rect 286142 244170 316434 244226
rect 316490 244170 316558 244226
rect 316614 244170 316682 244226
rect 316738 244170 316806 244226
rect 316862 244170 347154 244226
rect 347210 244170 347278 244226
rect 347334 244170 347402 244226
rect 347458 244170 347526 244226
rect 347582 244170 377874 244226
rect 377930 244170 377998 244226
rect 378054 244170 378122 244226
rect 378178 244170 378246 244226
rect 378302 244170 408594 244226
rect 408650 244170 408718 244226
rect 408774 244170 408842 244226
rect 408898 244170 408966 244226
rect 409022 244170 439314 244226
rect 439370 244170 439438 244226
rect 439494 244170 439562 244226
rect 439618 244170 439686 244226
rect 439742 244170 470034 244226
rect 470090 244170 470158 244226
rect 470214 244170 470282 244226
rect 470338 244170 470406 244226
rect 470462 244170 500754 244226
rect 500810 244170 500878 244226
rect 500934 244170 501002 244226
rect 501058 244170 501126 244226
rect 501182 244170 531474 244226
rect 531530 244170 531598 244226
rect 531654 244170 531722 244226
rect 531778 244170 531846 244226
rect 531902 244170 562194 244226
rect 562250 244170 562318 244226
rect 562374 244170 562442 244226
rect 562498 244170 562566 244226
rect 562622 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect -1916 244102 597980 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 9234 244102
rect 9290 244046 9358 244102
rect 9414 244046 9482 244102
rect 9538 244046 9606 244102
rect 9662 244046 39954 244102
rect 40010 244046 40078 244102
rect 40134 244046 40202 244102
rect 40258 244046 40326 244102
rect 40382 244046 59878 244102
rect 59934 244046 60002 244102
rect 60058 244046 70674 244102
rect 70730 244046 70798 244102
rect 70854 244046 70922 244102
rect 70978 244046 71046 244102
rect 71102 244046 90598 244102
rect 90654 244046 90722 244102
rect 90778 244046 101394 244102
rect 101450 244046 101518 244102
rect 101574 244046 101642 244102
rect 101698 244046 101766 244102
rect 101822 244046 132114 244102
rect 132170 244046 132238 244102
rect 132294 244046 132362 244102
rect 132418 244046 132486 244102
rect 132542 244046 162834 244102
rect 162890 244046 162958 244102
rect 163014 244046 163082 244102
rect 163138 244046 163206 244102
rect 163262 244046 193554 244102
rect 193610 244046 193678 244102
rect 193734 244046 193802 244102
rect 193858 244046 193926 244102
rect 193982 244046 224274 244102
rect 224330 244046 224398 244102
rect 224454 244046 224522 244102
rect 224578 244046 224646 244102
rect 224702 244046 254994 244102
rect 255050 244046 255118 244102
rect 255174 244046 255242 244102
rect 255298 244046 255366 244102
rect 255422 244046 285714 244102
rect 285770 244046 285838 244102
rect 285894 244046 285962 244102
rect 286018 244046 286086 244102
rect 286142 244046 316434 244102
rect 316490 244046 316558 244102
rect 316614 244046 316682 244102
rect 316738 244046 316806 244102
rect 316862 244046 347154 244102
rect 347210 244046 347278 244102
rect 347334 244046 347402 244102
rect 347458 244046 347526 244102
rect 347582 244046 377874 244102
rect 377930 244046 377998 244102
rect 378054 244046 378122 244102
rect 378178 244046 378246 244102
rect 378302 244046 408594 244102
rect 408650 244046 408718 244102
rect 408774 244046 408842 244102
rect 408898 244046 408966 244102
rect 409022 244046 439314 244102
rect 439370 244046 439438 244102
rect 439494 244046 439562 244102
rect 439618 244046 439686 244102
rect 439742 244046 470034 244102
rect 470090 244046 470158 244102
rect 470214 244046 470282 244102
rect 470338 244046 470406 244102
rect 470462 244046 500754 244102
rect 500810 244046 500878 244102
rect 500934 244046 501002 244102
rect 501058 244046 501126 244102
rect 501182 244046 531474 244102
rect 531530 244046 531598 244102
rect 531654 244046 531722 244102
rect 531778 244046 531846 244102
rect 531902 244046 562194 244102
rect 562250 244046 562318 244102
rect 562374 244046 562442 244102
rect 562498 244046 562566 244102
rect 562622 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect -1916 243978 597980 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 9234 243978
rect 9290 243922 9358 243978
rect 9414 243922 9482 243978
rect 9538 243922 9606 243978
rect 9662 243922 39954 243978
rect 40010 243922 40078 243978
rect 40134 243922 40202 243978
rect 40258 243922 40326 243978
rect 40382 243922 59878 243978
rect 59934 243922 60002 243978
rect 60058 243922 70674 243978
rect 70730 243922 70798 243978
rect 70854 243922 70922 243978
rect 70978 243922 71046 243978
rect 71102 243922 90598 243978
rect 90654 243922 90722 243978
rect 90778 243922 101394 243978
rect 101450 243922 101518 243978
rect 101574 243922 101642 243978
rect 101698 243922 101766 243978
rect 101822 243922 132114 243978
rect 132170 243922 132238 243978
rect 132294 243922 132362 243978
rect 132418 243922 132486 243978
rect 132542 243922 162834 243978
rect 162890 243922 162958 243978
rect 163014 243922 163082 243978
rect 163138 243922 163206 243978
rect 163262 243922 193554 243978
rect 193610 243922 193678 243978
rect 193734 243922 193802 243978
rect 193858 243922 193926 243978
rect 193982 243922 224274 243978
rect 224330 243922 224398 243978
rect 224454 243922 224522 243978
rect 224578 243922 224646 243978
rect 224702 243922 254994 243978
rect 255050 243922 255118 243978
rect 255174 243922 255242 243978
rect 255298 243922 255366 243978
rect 255422 243922 285714 243978
rect 285770 243922 285838 243978
rect 285894 243922 285962 243978
rect 286018 243922 286086 243978
rect 286142 243922 316434 243978
rect 316490 243922 316558 243978
rect 316614 243922 316682 243978
rect 316738 243922 316806 243978
rect 316862 243922 347154 243978
rect 347210 243922 347278 243978
rect 347334 243922 347402 243978
rect 347458 243922 347526 243978
rect 347582 243922 377874 243978
rect 377930 243922 377998 243978
rect 378054 243922 378122 243978
rect 378178 243922 378246 243978
rect 378302 243922 408594 243978
rect 408650 243922 408718 243978
rect 408774 243922 408842 243978
rect 408898 243922 408966 243978
rect 409022 243922 439314 243978
rect 439370 243922 439438 243978
rect 439494 243922 439562 243978
rect 439618 243922 439686 243978
rect 439742 243922 470034 243978
rect 470090 243922 470158 243978
rect 470214 243922 470282 243978
rect 470338 243922 470406 243978
rect 470462 243922 500754 243978
rect 500810 243922 500878 243978
rect 500934 243922 501002 243978
rect 501058 243922 501126 243978
rect 501182 243922 531474 243978
rect 531530 243922 531598 243978
rect 531654 243922 531722 243978
rect 531778 243922 531846 243978
rect 531902 243922 562194 243978
rect 562250 243922 562318 243978
rect 562374 243922 562442 243978
rect 562498 243922 562566 243978
rect 562622 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect -1916 243826 597980 243922
rect -1916 238350 597980 238446
rect -1916 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 36234 238350
rect 36290 238294 36358 238350
rect 36414 238294 36482 238350
rect 36538 238294 36606 238350
rect 36662 238294 66954 238350
rect 67010 238294 67078 238350
rect 67134 238294 67202 238350
rect 67258 238294 67326 238350
rect 67382 238294 97674 238350
rect 97730 238294 97798 238350
rect 97854 238294 97922 238350
rect 97978 238294 98046 238350
rect 98102 238294 128394 238350
rect 128450 238294 128518 238350
rect 128574 238294 128642 238350
rect 128698 238294 128766 238350
rect 128822 238294 159114 238350
rect 159170 238294 159238 238350
rect 159294 238294 159362 238350
rect 159418 238294 159486 238350
rect 159542 238294 189834 238350
rect 189890 238294 189958 238350
rect 190014 238294 190082 238350
rect 190138 238294 190206 238350
rect 190262 238294 220554 238350
rect 220610 238294 220678 238350
rect 220734 238294 220802 238350
rect 220858 238294 220926 238350
rect 220982 238294 251274 238350
rect 251330 238294 251398 238350
rect 251454 238294 251522 238350
rect 251578 238294 251646 238350
rect 251702 238294 281994 238350
rect 282050 238294 282118 238350
rect 282174 238294 282242 238350
rect 282298 238294 282366 238350
rect 282422 238294 312714 238350
rect 312770 238294 312838 238350
rect 312894 238294 312962 238350
rect 313018 238294 313086 238350
rect 313142 238294 343434 238350
rect 343490 238294 343558 238350
rect 343614 238294 343682 238350
rect 343738 238294 343806 238350
rect 343862 238294 374154 238350
rect 374210 238294 374278 238350
rect 374334 238294 374402 238350
rect 374458 238294 374526 238350
rect 374582 238294 404874 238350
rect 404930 238294 404998 238350
rect 405054 238294 405122 238350
rect 405178 238294 405246 238350
rect 405302 238294 435594 238350
rect 435650 238294 435718 238350
rect 435774 238294 435842 238350
rect 435898 238294 435966 238350
rect 436022 238294 466314 238350
rect 466370 238294 466438 238350
rect 466494 238294 466562 238350
rect 466618 238294 466686 238350
rect 466742 238294 497034 238350
rect 497090 238294 497158 238350
rect 497214 238294 497282 238350
rect 497338 238294 497406 238350
rect 497462 238294 527754 238350
rect 527810 238294 527878 238350
rect 527934 238294 528002 238350
rect 528058 238294 528126 238350
rect 528182 238294 558474 238350
rect 558530 238294 558598 238350
rect 558654 238294 558722 238350
rect 558778 238294 558846 238350
rect 558902 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597980 238350
rect -1916 238226 597980 238294
rect -1916 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 36234 238226
rect 36290 238170 36358 238226
rect 36414 238170 36482 238226
rect 36538 238170 36606 238226
rect 36662 238170 66954 238226
rect 67010 238170 67078 238226
rect 67134 238170 67202 238226
rect 67258 238170 67326 238226
rect 67382 238170 97674 238226
rect 97730 238170 97798 238226
rect 97854 238170 97922 238226
rect 97978 238170 98046 238226
rect 98102 238170 128394 238226
rect 128450 238170 128518 238226
rect 128574 238170 128642 238226
rect 128698 238170 128766 238226
rect 128822 238170 159114 238226
rect 159170 238170 159238 238226
rect 159294 238170 159362 238226
rect 159418 238170 159486 238226
rect 159542 238170 189834 238226
rect 189890 238170 189958 238226
rect 190014 238170 190082 238226
rect 190138 238170 190206 238226
rect 190262 238170 220554 238226
rect 220610 238170 220678 238226
rect 220734 238170 220802 238226
rect 220858 238170 220926 238226
rect 220982 238170 251274 238226
rect 251330 238170 251398 238226
rect 251454 238170 251522 238226
rect 251578 238170 251646 238226
rect 251702 238170 281994 238226
rect 282050 238170 282118 238226
rect 282174 238170 282242 238226
rect 282298 238170 282366 238226
rect 282422 238170 312714 238226
rect 312770 238170 312838 238226
rect 312894 238170 312962 238226
rect 313018 238170 313086 238226
rect 313142 238170 343434 238226
rect 343490 238170 343558 238226
rect 343614 238170 343682 238226
rect 343738 238170 343806 238226
rect 343862 238170 374154 238226
rect 374210 238170 374278 238226
rect 374334 238170 374402 238226
rect 374458 238170 374526 238226
rect 374582 238170 404874 238226
rect 404930 238170 404998 238226
rect 405054 238170 405122 238226
rect 405178 238170 405246 238226
rect 405302 238170 435594 238226
rect 435650 238170 435718 238226
rect 435774 238170 435842 238226
rect 435898 238170 435966 238226
rect 436022 238170 466314 238226
rect 466370 238170 466438 238226
rect 466494 238170 466562 238226
rect 466618 238170 466686 238226
rect 466742 238170 497034 238226
rect 497090 238170 497158 238226
rect 497214 238170 497282 238226
rect 497338 238170 497406 238226
rect 497462 238170 527754 238226
rect 527810 238170 527878 238226
rect 527934 238170 528002 238226
rect 528058 238170 528126 238226
rect 528182 238170 558474 238226
rect 558530 238170 558598 238226
rect 558654 238170 558722 238226
rect 558778 238170 558846 238226
rect 558902 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597980 238226
rect -1916 238102 597980 238170
rect -1916 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 36234 238102
rect 36290 238046 36358 238102
rect 36414 238046 36482 238102
rect 36538 238046 36606 238102
rect 36662 238046 66954 238102
rect 67010 238046 67078 238102
rect 67134 238046 67202 238102
rect 67258 238046 67326 238102
rect 67382 238046 97674 238102
rect 97730 238046 97798 238102
rect 97854 238046 97922 238102
rect 97978 238046 98046 238102
rect 98102 238046 128394 238102
rect 128450 238046 128518 238102
rect 128574 238046 128642 238102
rect 128698 238046 128766 238102
rect 128822 238046 159114 238102
rect 159170 238046 159238 238102
rect 159294 238046 159362 238102
rect 159418 238046 159486 238102
rect 159542 238046 189834 238102
rect 189890 238046 189958 238102
rect 190014 238046 190082 238102
rect 190138 238046 190206 238102
rect 190262 238046 220554 238102
rect 220610 238046 220678 238102
rect 220734 238046 220802 238102
rect 220858 238046 220926 238102
rect 220982 238046 251274 238102
rect 251330 238046 251398 238102
rect 251454 238046 251522 238102
rect 251578 238046 251646 238102
rect 251702 238046 281994 238102
rect 282050 238046 282118 238102
rect 282174 238046 282242 238102
rect 282298 238046 282366 238102
rect 282422 238046 312714 238102
rect 312770 238046 312838 238102
rect 312894 238046 312962 238102
rect 313018 238046 313086 238102
rect 313142 238046 343434 238102
rect 343490 238046 343558 238102
rect 343614 238046 343682 238102
rect 343738 238046 343806 238102
rect 343862 238046 374154 238102
rect 374210 238046 374278 238102
rect 374334 238046 374402 238102
rect 374458 238046 374526 238102
rect 374582 238046 404874 238102
rect 404930 238046 404998 238102
rect 405054 238046 405122 238102
rect 405178 238046 405246 238102
rect 405302 238046 435594 238102
rect 435650 238046 435718 238102
rect 435774 238046 435842 238102
rect 435898 238046 435966 238102
rect 436022 238046 466314 238102
rect 466370 238046 466438 238102
rect 466494 238046 466562 238102
rect 466618 238046 466686 238102
rect 466742 238046 497034 238102
rect 497090 238046 497158 238102
rect 497214 238046 497282 238102
rect 497338 238046 497406 238102
rect 497462 238046 527754 238102
rect 527810 238046 527878 238102
rect 527934 238046 528002 238102
rect 528058 238046 528126 238102
rect 528182 238046 558474 238102
rect 558530 238046 558598 238102
rect 558654 238046 558722 238102
rect 558778 238046 558846 238102
rect 558902 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597980 238102
rect -1916 237978 597980 238046
rect -1916 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 36234 237978
rect 36290 237922 36358 237978
rect 36414 237922 36482 237978
rect 36538 237922 36606 237978
rect 36662 237922 66954 237978
rect 67010 237922 67078 237978
rect 67134 237922 67202 237978
rect 67258 237922 67326 237978
rect 67382 237922 97674 237978
rect 97730 237922 97798 237978
rect 97854 237922 97922 237978
rect 97978 237922 98046 237978
rect 98102 237922 128394 237978
rect 128450 237922 128518 237978
rect 128574 237922 128642 237978
rect 128698 237922 128766 237978
rect 128822 237922 159114 237978
rect 159170 237922 159238 237978
rect 159294 237922 159362 237978
rect 159418 237922 159486 237978
rect 159542 237922 189834 237978
rect 189890 237922 189958 237978
rect 190014 237922 190082 237978
rect 190138 237922 190206 237978
rect 190262 237922 220554 237978
rect 220610 237922 220678 237978
rect 220734 237922 220802 237978
rect 220858 237922 220926 237978
rect 220982 237922 251274 237978
rect 251330 237922 251398 237978
rect 251454 237922 251522 237978
rect 251578 237922 251646 237978
rect 251702 237922 281994 237978
rect 282050 237922 282118 237978
rect 282174 237922 282242 237978
rect 282298 237922 282366 237978
rect 282422 237922 312714 237978
rect 312770 237922 312838 237978
rect 312894 237922 312962 237978
rect 313018 237922 313086 237978
rect 313142 237922 343434 237978
rect 343490 237922 343558 237978
rect 343614 237922 343682 237978
rect 343738 237922 343806 237978
rect 343862 237922 374154 237978
rect 374210 237922 374278 237978
rect 374334 237922 374402 237978
rect 374458 237922 374526 237978
rect 374582 237922 404874 237978
rect 404930 237922 404998 237978
rect 405054 237922 405122 237978
rect 405178 237922 405246 237978
rect 405302 237922 435594 237978
rect 435650 237922 435718 237978
rect 435774 237922 435842 237978
rect 435898 237922 435966 237978
rect 436022 237922 466314 237978
rect 466370 237922 466438 237978
rect 466494 237922 466562 237978
rect 466618 237922 466686 237978
rect 466742 237922 497034 237978
rect 497090 237922 497158 237978
rect 497214 237922 497282 237978
rect 497338 237922 497406 237978
rect 497462 237922 527754 237978
rect 527810 237922 527878 237978
rect 527934 237922 528002 237978
rect 528058 237922 528126 237978
rect 528182 237922 558474 237978
rect 558530 237922 558598 237978
rect 558654 237922 558722 237978
rect 558778 237922 558846 237978
rect 558902 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597980 237978
rect -1916 237826 597980 237922
rect 76956 237718 103364 237734
rect 76956 237662 76972 237718
rect 77028 237662 103292 237718
rect 103348 237662 103364 237718
rect 76956 237646 103364 237662
rect 74940 237538 100004 237554
rect 74940 237482 74956 237538
rect 75012 237482 99932 237538
rect 99988 237482 100004 237538
rect 74940 237466 100004 237482
rect -1916 226350 597980 226446
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 9234 226350
rect 9290 226294 9358 226350
rect 9414 226294 9482 226350
rect 9538 226294 9606 226350
rect 9662 226294 39954 226350
rect 40010 226294 40078 226350
rect 40134 226294 40202 226350
rect 40258 226294 40326 226350
rect 40382 226294 70674 226350
rect 70730 226294 70798 226350
rect 70854 226294 70922 226350
rect 70978 226294 71046 226350
rect 71102 226294 101394 226350
rect 101450 226294 101518 226350
rect 101574 226294 101642 226350
rect 101698 226294 101766 226350
rect 101822 226294 132114 226350
rect 132170 226294 132238 226350
rect 132294 226294 132362 226350
rect 132418 226294 132486 226350
rect 132542 226294 162834 226350
rect 162890 226294 162958 226350
rect 163014 226294 163082 226350
rect 163138 226294 163206 226350
rect 163262 226294 193554 226350
rect 193610 226294 193678 226350
rect 193734 226294 193802 226350
rect 193858 226294 193926 226350
rect 193982 226294 224274 226350
rect 224330 226294 224398 226350
rect 224454 226294 224522 226350
rect 224578 226294 224646 226350
rect 224702 226294 254994 226350
rect 255050 226294 255118 226350
rect 255174 226294 255242 226350
rect 255298 226294 255366 226350
rect 255422 226294 285714 226350
rect 285770 226294 285838 226350
rect 285894 226294 285962 226350
rect 286018 226294 286086 226350
rect 286142 226294 316434 226350
rect 316490 226294 316558 226350
rect 316614 226294 316682 226350
rect 316738 226294 316806 226350
rect 316862 226294 347154 226350
rect 347210 226294 347278 226350
rect 347334 226294 347402 226350
rect 347458 226294 347526 226350
rect 347582 226294 377874 226350
rect 377930 226294 377998 226350
rect 378054 226294 378122 226350
rect 378178 226294 378246 226350
rect 378302 226294 408594 226350
rect 408650 226294 408718 226350
rect 408774 226294 408842 226350
rect 408898 226294 408966 226350
rect 409022 226294 439314 226350
rect 439370 226294 439438 226350
rect 439494 226294 439562 226350
rect 439618 226294 439686 226350
rect 439742 226294 470034 226350
rect 470090 226294 470158 226350
rect 470214 226294 470282 226350
rect 470338 226294 470406 226350
rect 470462 226294 489822 226350
rect 489878 226294 489946 226350
rect 490002 226294 498390 226350
rect 498446 226294 498514 226350
rect 498570 226294 506958 226350
rect 507014 226294 507082 226350
rect 507138 226294 515526 226350
rect 515582 226294 515650 226350
rect 515706 226294 531474 226350
rect 531530 226294 531598 226350
rect 531654 226294 531722 226350
rect 531778 226294 531846 226350
rect 531902 226294 562194 226350
rect 562250 226294 562318 226350
rect 562374 226294 562442 226350
rect 562498 226294 562566 226350
rect 562622 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect -1916 226226 597980 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 9234 226226
rect 9290 226170 9358 226226
rect 9414 226170 9482 226226
rect 9538 226170 9606 226226
rect 9662 226170 39954 226226
rect 40010 226170 40078 226226
rect 40134 226170 40202 226226
rect 40258 226170 40326 226226
rect 40382 226170 70674 226226
rect 70730 226170 70798 226226
rect 70854 226170 70922 226226
rect 70978 226170 71046 226226
rect 71102 226170 101394 226226
rect 101450 226170 101518 226226
rect 101574 226170 101642 226226
rect 101698 226170 101766 226226
rect 101822 226170 132114 226226
rect 132170 226170 132238 226226
rect 132294 226170 132362 226226
rect 132418 226170 132486 226226
rect 132542 226170 162834 226226
rect 162890 226170 162958 226226
rect 163014 226170 163082 226226
rect 163138 226170 163206 226226
rect 163262 226170 193554 226226
rect 193610 226170 193678 226226
rect 193734 226170 193802 226226
rect 193858 226170 193926 226226
rect 193982 226170 224274 226226
rect 224330 226170 224398 226226
rect 224454 226170 224522 226226
rect 224578 226170 224646 226226
rect 224702 226170 254994 226226
rect 255050 226170 255118 226226
rect 255174 226170 255242 226226
rect 255298 226170 255366 226226
rect 255422 226170 285714 226226
rect 285770 226170 285838 226226
rect 285894 226170 285962 226226
rect 286018 226170 286086 226226
rect 286142 226170 316434 226226
rect 316490 226170 316558 226226
rect 316614 226170 316682 226226
rect 316738 226170 316806 226226
rect 316862 226170 347154 226226
rect 347210 226170 347278 226226
rect 347334 226170 347402 226226
rect 347458 226170 347526 226226
rect 347582 226170 377874 226226
rect 377930 226170 377998 226226
rect 378054 226170 378122 226226
rect 378178 226170 378246 226226
rect 378302 226170 408594 226226
rect 408650 226170 408718 226226
rect 408774 226170 408842 226226
rect 408898 226170 408966 226226
rect 409022 226170 439314 226226
rect 439370 226170 439438 226226
rect 439494 226170 439562 226226
rect 439618 226170 439686 226226
rect 439742 226170 470034 226226
rect 470090 226170 470158 226226
rect 470214 226170 470282 226226
rect 470338 226170 470406 226226
rect 470462 226170 489822 226226
rect 489878 226170 489946 226226
rect 490002 226170 498390 226226
rect 498446 226170 498514 226226
rect 498570 226170 506958 226226
rect 507014 226170 507082 226226
rect 507138 226170 515526 226226
rect 515582 226170 515650 226226
rect 515706 226170 531474 226226
rect 531530 226170 531598 226226
rect 531654 226170 531722 226226
rect 531778 226170 531846 226226
rect 531902 226170 562194 226226
rect 562250 226170 562318 226226
rect 562374 226170 562442 226226
rect 562498 226170 562566 226226
rect 562622 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect -1916 226102 597980 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 9234 226102
rect 9290 226046 9358 226102
rect 9414 226046 9482 226102
rect 9538 226046 9606 226102
rect 9662 226046 39954 226102
rect 40010 226046 40078 226102
rect 40134 226046 40202 226102
rect 40258 226046 40326 226102
rect 40382 226046 70674 226102
rect 70730 226046 70798 226102
rect 70854 226046 70922 226102
rect 70978 226046 71046 226102
rect 71102 226046 101394 226102
rect 101450 226046 101518 226102
rect 101574 226046 101642 226102
rect 101698 226046 101766 226102
rect 101822 226046 132114 226102
rect 132170 226046 132238 226102
rect 132294 226046 132362 226102
rect 132418 226046 132486 226102
rect 132542 226046 162834 226102
rect 162890 226046 162958 226102
rect 163014 226046 163082 226102
rect 163138 226046 163206 226102
rect 163262 226046 193554 226102
rect 193610 226046 193678 226102
rect 193734 226046 193802 226102
rect 193858 226046 193926 226102
rect 193982 226046 224274 226102
rect 224330 226046 224398 226102
rect 224454 226046 224522 226102
rect 224578 226046 224646 226102
rect 224702 226046 254994 226102
rect 255050 226046 255118 226102
rect 255174 226046 255242 226102
rect 255298 226046 255366 226102
rect 255422 226046 285714 226102
rect 285770 226046 285838 226102
rect 285894 226046 285962 226102
rect 286018 226046 286086 226102
rect 286142 226046 316434 226102
rect 316490 226046 316558 226102
rect 316614 226046 316682 226102
rect 316738 226046 316806 226102
rect 316862 226046 347154 226102
rect 347210 226046 347278 226102
rect 347334 226046 347402 226102
rect 347458 226046 347526 226102
rect 347582 226046 377874 226102
rect 377930 226046 377998 226102
rect 378054 226046 378122 226102
rect 378178 226046 378246 226102
rect 378302 226046 408594 226102
rect 408650 226046 408718 226102
rect 408774 226046 408842 226102
rect 408898 226046 408966 226102
rect 409022 226046 439314 226102
rect 439370 226046 439438 226102
rect 439494 226046 439562 226102
rect 439618 226046 439686 226102
rect 439742 226046 470034 226102
rect 470090 226046 470158 226102
rect 470214 226046 470282 226102
rect 470338 226046 470406 226102
rect 470462 226046 489822 226102
rect 489878 226046 489946 226102
rect 490002 226046 498390 226102
rect 498446 226046 498514 226102
rect 498570 226046 506958 226102
rect 507014 226046 507082 226102
rect 507138 226046 515526 226102
rect 515582 226046 515650 226102
rect 515706 226046 531474 226102
rect 531530 226046 531598 226102
rect 531654 226046 531722 226102
rect 531778 226046 531846 226102
rect 531902 226046 562194 226102
rect 562250 226046 562318 226102
rect 562374 226046 562442 226102
rect 562498 226046 562566 226102
rect 562622 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect -1916 225978 597980 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 9234 225978
rect 9290 225922 9358 225978
rect 9414 225922 9482 225978
rect 9538 225922 9606 225978
rect 9662 225922 39954 225978
rect 40010 225922 40078 225978
rect 40134 225922 40202 225978
rect 40258 225922 40326 225978
rect 40382 225922 70674 225978
rect 70730 225922 70798 225978
rect 70854 225922 70922 225978
rect 70978 225922 71046 225978
rect 71102 225922 101394 225978
rect 101450 225922 101518 225978
rect 101574 225922 101642 225978
rect 101698 225922 101766 225978
rect 101822 225922 132114 225978
rect 132170 225922 132238 225978
rect 132294 225922 132362 225978
rect 132418 225922 132486 225978
rect 132542 225922 162834 225978
rect 162890 225922 162958 225978
rect 163014 225922 163082 225978
rect 163138 225922 163206 225978
rect 163262 225922 193554 225978
rect 193610 225922 193678 225978
rect 193734 225922 193802 225978
rect 193858 225922 193926 225978
rect 193982 225922 224274 225978
rect 224330 225922 224398 225978
rect 224454 225922 224522 225978
rect 224578 225922 224646 225978
rect 224702 225922 254994 225978
rect 255050 225922 255118 225978
rect 255174 225922 255242 225978
rect 255298 225922 255366 225978
rect 255422 225922 285714 225978
rect 285770 225922 285838 225978
rect 285894 225922 285962 225978
rect 286018 225922 286086 225978
rect 286142 225922 316434 225978
rect 316490 225922 316558 225978
rect 316614 225922 316682 225978
rect 316738 225922 316806 225978
rect 316862 225922 347154 225978
rect 347210 225922 347278 225978
rect 347334 225922 347402 225978
rect 347458 225922 347526 225978
rect 347582 225922 377874 225978
rect 377930 225922 377998 225978
rect 378054 225922 378122 225978
rect 378178 225922 378246 225978
rect 378302 225922 408594 225978
rect 408650 225922 408718 225978
rect 408774 225922 408842 225978
rect 408898 225922 408966 225978
rect 409022 225922 439314 225978
rect 439370 225922 439438 225978
rect 439494 225922 439562 225978
rect 439618 225922 439686 225978
rect 439742 225922 470034 225978
rect 470090 225922 470158 225978
rect 470214 225922 470282 225978
rect 470338 225922 470406 225978
rect 470462 225922 489822 225978
rect 489878 225922 489946 225978
rect 490002 225922 498390 225978
rect 498446 225922 498514 225978
rect 498570 225922 506958 225978
rect 507014 225922 507082 225978
rect 507138 225922 515526 225978
rect 515582 225922 515650 225978
rect 515706 225922 531474 225978
rect 531530 225922 531598 225978
rect 531654 225922 531722 225978
rect 531778 225922 531846 225978
rect 531902 225922 562194 225978
rect 562250 225922 562318 225978
rect 562374 225922 562442 225978
rect 562498 225922 562566 225978
rect 562622 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect -1916 225826 597980 225922
rect -1916 220350 597980 220446
rect -1916 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 36234 220350
rect 36290 220294 36358 220350
rect 36414 220294 36482 220350
rect 36538 220294 36606 220350
rect 36662 220294 66954 220350
rect 67010 220294 67078 220350
rect 67134 220294 67202 220350
rect 67258 220294 67326 220350
rect 67382 220294 97674 220350
rect 97730 220294 97798 220350
rect 97854 220294 97922 220350
rect 97978 220294 98046 220350
rect 98102 220294 128394 220350
rect 128450 220294 128518 220350
rect 128574 220294 128642 220350
rect 128698 220294 128766 220350
rect 128822 220294 159114 220350
rect 159170 220294 159238 220350
rect 159294 220294 159362 220350
rect 159418 220294 159486 220350
rect 159542 220294 189834 220350
rect 189890 220294 189958 220350
rect 190014 220294 190082 220350
rect 190138 220294 190206 220350
rect 190262 220294 220554 220350
rect 220610 220294 220678 220350
rect 220734 220294 220802 220350
rect 220858 220294 220926 220350
rect 220982 220294 251274 220350
rect 251330 220294 251398 220350
rect 251454 220294 251522 220350
rect 251578 220294 251646 220350
rect 251702 220294 281994 220350
rect 282050 220294 282118 220350
rect 282174 220294 282242 220350
rect 282298 220294 282366 220350
rect 282422 220294 312714 220350
rect 312770 220294 312838 220350
rect 312894 220294 312962 220350
rect 313018 220294 313086 220350
rect 313142 220294 343434 220350
rect 343490 220294 343558 220350
rect 343614 220294 343682 220350
rect 343738 220294 343806 220350
rect 343862 220294 374154 220350
rect 374210 220294 374278 220350
rect 374334 220294 374402 220350
rect 374458 220294 374526 220350
rect 374582 220294 404874 220350
rect 404930 220294 404998 220350
rect 405054 220294 405122 220350
rect 405178 220294 405246 220350
rect 405302 220294 435594 220350
rect 435650 220294 435718 220350
rect 435774 220294 435842 220350
rect 435898 220294 435966 220350
rect 436022 220294 466314 220350
rect 466370 220294 466438 220350
rect 466494 220294 466562 220350
rect 466618 220294 466686 220350
rect 466742 220294 485538 220350
rect 485594 220294 485662 220350
rect 485718 220294 494106 220350
rect 494162 220294 494230 220350
rect 494286 220294 502674 220350
rect 502730 220294 502798 220350
rect 502854 220294 511242 220350
rect 511298 220294 511366 220350
rect 511422 220294 527754 220350
rect 527810 220294 527878 220350
rect 527934 220294 528002 220350
rect 528058 220294 528126 220350
rect 528182 220294 558474 220350
rect 558530 220294 558598 220350
rect 558654 220294 558722 220350
rect 558778 220294 558846 220350
rect 558902 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597980 220350
rect -1916 220226 597980 220294
rect -1916 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 36234 220226
rect 36290 220170 36358 220226
rect 36414 220170 36482 220226
rect 36538 220170 36606 220226
rect 36662 220170 66954 220226
rect 67010 220170 67078 220226
rect 67134 220170 67202 220226
rect 67258 220170 67326 220226
rect 67382 220170 97674 220226
rect 97730 220170 97798 220226
rect 97854 220170 97922 220226
rect 97978 220170 98046 220226
rect 98102 220170 128394 220226
rect 128450 220170 128518 220226
rect 128574 220170 128642 220226
rect 128698 220170 128766 220226
rect 128822 220170 159114 220226
rect 159170 220170 159238 220226
rect 159294 220170 159362 220226
rect 159418 220170 159486 220226
rect 159542 220170 189834 220226
rect 189890 220170 189958 220226
rect 190014 220170 190082 220226
rect 190138 220170 190206 220226
rect 190262 220170 220554 220226
rect 220610 220170 220678 220226
rect 220734 220170 220802 220226
rect 220858 220170 220926 220226
rect 220982 220170 251274 220226
rect 251330 220170 251398 220226
rect 251454 220170 251522 220226
rect 251578 220170 251646 220226
rect 251702 220170 281994 220226
rect 282050 220170 282118 220226
rect 282174 220170 282242 220226
rect 282298 220170 282366 220226
rect 282422 220170 312714 220226
rect 312770 220170 312838 220226
rect 312894 220170 312962 220226
rect 313018 220170 313086 220226
rect 313142 220170 343434 220226
rect 343490 220170 343558 220226
rect 343614 220170 343682 220226
rect 343738 220170 343806 220226
rect 343862 220170 374154 220226
rect 374210 220170 374278 220226
rect 374334 220170 374402 220226
rect 374458 220170 374526 220226
rect 374582 220170 404874 220226
rect 404930 220170 404998 220226
rect 405054 220170 405122 220226
rect 405178 220170 405246 220226
rect 405302 220170 435594 220226
rect 435650 220170 435718 220226
rect 435774 220170 435842 220226
rect 435898 220170 435966 220226
rect 436022 220170 466314 220226
rect 466370 220170 466438 220226
rect 466494 220170 466562 220226
rect 466618 220170 466686 220226
rect 466742 220170 485538 220226
rect 485594 220170 485662 220226
rect 485718 220170 494106 220226
rect 494162 220170 494230 220226
rect 494286 220170 502674 220226
rect 502730 220170 502798 220226
rect 502854 220170 511242 220226
rect 511298 220170 511366 220226
rect 511422 220170 527754 220226
rect 527810 220170 527878 220226
rect 527934 220170 528002 220226
rect 528058 220170 528126 220226
rect 528182 220170 558474 220226
rect 558530 220170 558598 220226
rect 558654 220170 558722 220226
rect 558778 220170 558846 220226
rect 558902 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597980 220226
rect -1916 220102 597980 220170
rect -1916 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 36234 220102
rect 36290 220046 36358 220102
rect 36414 220046 36482 220102
rect 36538 220046 36606 220102
rect 36662 220046 66954 220102
rect 67010 220046 67078 220102
rect 67134 220046 67202 220102
rect 67258 220046 67326 220102
rect 67382 220046 97674 220102
rect 97730 220046 97798 220102
rect 97854 220046 97922 220102
rect 97978 220046 98046 220102
rect 98102 220046 128394 220102
rect 128450 220046 128518 220102
rect 128574 220046 128642 220102
rect 128698 220046 128766 220102
rect 128822 220046 159114 220102
rect 159170 220046 159238 220102
rect 159294 220046 159362 220102
rect 159418 220046 159486 220102
rect 159542 220046 189834 220102
rect 189890 220046 189958 220102
rect 190014 220046 190082 220102
rect 190138 220046 190206 220102
rect 190262 220046 220554 220102
rect 220610 220046 220678 220102
rect 220734 220046 220802 220102
rect 220858 220046 220926 220102
rect 220982 220046 251274 220102
rect 251330 220046 251398 220102
rect 251454 220046 251522 220102
rect 251578 220046 251646 220102
rect 251702 220046 281994 220102
rect 282050 220046 282118 220102
rect 282174 220046 282242 220102
rect 282298 220046 282366 220102
rect 282422 220046 312714 220102
rect 312770 220046 312838 220102
rect 312894 220046 312962 220102
rect 313018 220046 313086 220102
rect 313142 220046 343434 220102
rect 343490 220046 343558 220102
rect 343614 220046 343682 220102
rect 343738 220046 343806 220102
rect 343862 220046 374154 220102
rect 374210 220046 374278 220102
rect 374334 220046 374402 220102
rect 374458 220046 374526 220102
rect 374582 220046 404874 220102
rect 404930 220046 404998 220102
rect 405054 220046 405122 220102
rect 405178 220046 405246 220102
rect 405302 220046 435594 220102
rect 435650 220046 435718 220102
rect 435774 220046 435842 220102
rect 435898 220046 435966 220102
rect 436022 220046 466314 220102
rect 466370 220046 466438 220102
rect 466494 220046 466562 220102
rect 466618 220046 466686 220102
rect 466742 220046 485538 220102
rect 485594 220046 485662 220102
rect 485718 220046 494106 220102
rect 494162 220046 494230 220102
rect 494286 220046 502674 220102
rect 502730 220046 502798 220102
rect 502854 220046 511242 220102
rect 511298 220046 511366 220102
rect 511422 220046 527754 220102
rect 527810 220046 527878 220102
rect 527934 220046 528002 220102
rect 528058 220046 528126 220102
rect 528182 220046 558474 220102
rect 558530 220046 558598 220102
rect 558654 220046 558722 220102
rect 558778 220046 558846 220102
rect 558902 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597980 220102
rect -1916 219978 597980 220046
rect -1916 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 36234 219978
rect 36290 219922 36358 219978
rect 36414 219922 36482 219978
rect 36538 219922 36606 219978
rect 36662 219922 66954 219978
rect 67010 219922 67078 219978
rect 67134 219922 67202 219978
rect 67258 219922 67326 219978
rect 67382 219922 97674 219978
rect 97730 219922 97798 219978
rect 97854 219922 97922 219978
rect 97978 219922 98046 219978
rect 98102 219922 128394 219978
rect 128450 219922 128518 219978
rect 128574 219922 128642 219978
rect 128698 219922 128766 219978
rect 128822 219922 159114 219978
rect 159170 219922 159238 219978
rect 159294 219922 159362 219978
rect 159418 219922 159486 219978
rect 159542 219922 189834 219978
rect 189890 219922 189958 219978
rect 190014 219922 190082 219978
rect 190138 219922 190206 219978
rect 190262 219922 220554 219978
rect 220610 219922 220678 219978
rect 220734 219922 220802 219978
rect 220858 219922 220926 219978
rect 220982 219922 251274 219978
rect 251330 219922 251398 219978
rect 251454 219922 251522 219978
rect 251578 219922 251646 219978
rect 251702 219922 281994 219978
rect 282050 219922 282118 219978
rect 282174 219922 282242 219978
rect 282298 219922 282366 219978
rect 282422 219922 312714 219978
rect 312770 219922 312838 219978
rect 312894 219922 312962 219978
rect 313018 219922 313086 219978
rect 313142 219922 343434 219978
rect 343490 219922 343558 219978
rect 343614 219922 343682 219978
rect 343738 219922 343806 219978
rect 343862 219922 374154 219978
rect 374210 219922 374278 219978
rect 374334 219922 374402 219978
rect 374458 219922 374526 219978
rect 374582 219922 404874 219978
rect 404930 219922 404998 219978
rect 405054 219922 405122 219978
rect 405178 219922 405246 219978
rect 405302 219922 435594 219978
rect 435650 219922 435718 219978
rect 435774 219922 435842 219978
rect 435898 219922 435966 219978
rect 436022 219922 466314 219978
rect 466370 219922 466438 219978
rect 466494 219922 466562 219978
rect 466618 219922 466686 219978
rect 466742 219922 485538 219978
rect 485594 219922 485662 219978
rect 485718 219922 494106 219978
rect 494162 219922 494230 219978
rect 494286 219922 502674 219978
rect 502730 219922 502798 219978
rect 502854 219922 511242 219978
rect 511298 219922 511366 219978
rect 511422 219922 527754 219978
rect 527810 219922 527878 219978
rect 527934 219922 528002 219978
rect 528058 219922 528126 219978
rect 528182 219922 558474 219978
rect 558530 219922 558598 219978
rect 558654 219922 558722 219978
rect 558778 219922 558846 219978
rect 558902 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597980 219978
rect -1916 219826 597980 219922
rect 236220 211078 291636 211094
rect 236220 211022 236236 211078
rect 236292 211022 291564 211078
rect 291620 211022 291636 211078
rect 236220 211006 291636 211022
rect 237900 210898 296564 210914
rect 237900 210842 237916 210898
rect 237972 210842 296492 210898
rect 296548 210842 296564 210898
rect 237900 210826 296564 210842
rect -1916 208350 597980 208446
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 9234 208350
rect 9290 208294 9358 208350
rect 9414 208294 9482 208350
rect 9538 208294 9606 208350
rect 9662 208294 39954 208350
rect 40010 208294 40078 208350
rect 40134 208294 40202 208350
rect 40258 208294 40326 208350
rect 40382 208294 285714 208350
rect 285770 208294 285838 208350
rect 285894 208294 285962 208350
rect 286018 208294 286086 208350
rect 286142 208294 316434 208350
rect 316490 208294 316558 208350
rect 316614 208294 316682 208350
rect 316738 208294 316806 208350
rect 316862 208294 347154 208350
rect 347210 208294 347278 208350
rect 347334 208294 347402 208350
rect 347458 208294 347526 208350
rect 347582 208294 377874 208350
rect 377930 208294 377998 208350
rect 378054 208294 378122 208350
rect 378178 208294 378246 208350
rect 378302 208294 408594 208350
rect 408650 208294 408718 208350
rect 408774 208294 408842 208350
rect 408898 208294 408966 208350
rect 409022 208294 439314 208350
rect 439370 208294 439438 208350
rect 439494 208294 439562 208350
rect 439618 208294 439686 208350
rect 439742 208294 470034 208350
rect 470090 208294 470158 208350
rect 470214 208294 470282 208350
rect 470338 208294 470406 208350
rect 470462 208294 489822 208350
rect 489878 208294 489946 208350
rect 490002 208294 498390 208350
rect 498446 208294 498514 208350
rect 498570 208294 506958 208350
rect 507014 208294 507082 208350
rect 507138 208294 515526 208350
rect 515582 208294 515650 208350
rect 515706 208294 531474 208350
rect 531530 208294 531598 208350
rect 531654 208294 531722 208350
rect 531778 208294 531846 208350
rect 531902 208294 562194 208350
rect 562250 208294 562318 208350
rect 562374 208294 562442 208350
rect 562498 208294 562566 208350
rect 562622 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect -1916 208226 597980 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 9234 208226
rect 9290 208170 9358 208226
rect 9414 208170 9482 208226
rect 9538 208170 9606 208226
rect 9662 208170 39954 208226
rect 40010 208170 40078 208226
rect 40134 208170 40202 208226
rect 40258 208170 40326 208226
rect 40382 208170 285714 208226
rect 285770 208170 285838 208226
rect 285894 208170 285962 208226
rect 286018 208170 286086 208226
rect 286142 208170 316434 208226
rect 316490 208170 316558 208226
rect 316614 208170 316682 208226
rect 316738 208170 316806 208226
rect 316862 208170 347154 208226
rect 347210 208170 347278 208226
rect 347334 208170 347402 208226
rect 347458 208170 347526 208226
rect 347582 208170 377874 208226
rect 377930 208170 377998 208226
rect 378054 208170 378122 208226
rect 378178 208170 378246 208226
rect 378302 208170 408594 208226
rect 408650 208170 408718 208226
rect 408774 208170 408842 208226
rect 408898 208170 408966 208226
rect 409022 208170 439314 208226
rect 439370 208170 439438 208226
rect 439494 208170 439562 208226
rect 439618 208170 439686 208226
rect 439742 208170 470034 208226
rect 470090 208170 470158 208226
rect 470214 208170 470282 208226
rect 470338 208170 470406 208226
rect 470462 208170 489822 208226
rect 489878 208170 489946 208226
rect 490002 208170 498390 208226
rect 498446 208170 498514 208226
rect 498570 208170 506958 208226
rect 507014 208170 507082 208226
rect 507138 208170 515526 208226
rect 515582 208170 515650 208226
rect 515706 208170 531474 208226
rect 531530 208170 531598 208226
rect 531654 208170 531722 208226
rect 531778 208170 531846 208226
rect 531902 208170 562194 208226
rect 562250 208170 562318 208226
rect 562374 208170 562442 208226
rect 562498 208170 562566 208226
rect 562622 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect -1916 208102 597980 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 9234 208102
rect 9290 208046 9358 208102
rect 9414 208046 9482 208102
rect 9538 208046 9606 208102
rect 9662 208046 39954 208102
rect 40010 208046 40078 208102
rect 40134 208046 40202 208102
rect 40258 208046 40326 208102
rect 40382 208046 285714 208102
rect 285770 208046 285838 208102
rect 285894 208046 285962 208102
rect 286018 208046 286086 208102
rect 286142 208046 316434 208102
rect 316490 208046 316558 208102
rect 316614 208046 316682 208102
rect 316738 208046 316806 208102
rect 316862 208046 347154 208102
rect 347210 208046 347278 208102
rect 347334 208046 347402 208102
rect 347458 208046 347526 208102
rect 347582 208046 377874 208102
rect 377930 208046 377998 208102
rect 378054 208046 378122 208102
rect 378178 208046 378246 208102
rect 378302 208046 408594 208102
rect 408650 208046 408718 208102
rect 408774 208046 408842 208102
rect 408898 208046 408966 208102
rect 409022 208046 439314 208102
rect 439370 208046 439438 208102
rect 439494 208046 439562 208102
rect 439618 208046 439686 208102
rect 439742 208046 470034 208102
rect 470090 208046 470158 208102
rect 470214 208046 470282 208102
rect 470338 208046 470406 208102
rect 470462 208046 489822 208102
rect 489878 208046 489946 208102
rect 490002 208046 498390 208102
rect 498446 208046 498514 208102
rect 498570 208046 506958 208102
rect 507014 208046 507082 208102
rect 507138 208046 515526 208102
rect 515582 208046 515650 208102
rect 515706 208046 531474 208102
rect 531530 208046 531598 208102
rect 531654 208046 531722 208102
rect 531778 208046 531846 208102
rect 531902 208046 562194 208102
rect 562250 208046 562318 208102
rect 562374 208046 562442 208102
rect 562498 208046 562566 208102
rect 562622 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect -1916 207978 597980 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 9234 207978
rect 9290 207922 9358 207978
rect 9414 207922 9482 207978
rect 9538 207922 9606 207978
rect 9662 207922 39954 207978
rect 40010 207922 40078 207978
rect 40134 207922 40202 207978
rect 40258 207922 40326 207978
rect 40382 207922 285714 207978
rect 285770 207922 285838 207978
rect 285894 207922 285962 207978
rect 286018 207922 286086 207978
rect 286142 207922 316434 207978
rect 316490 207922 316558 207978
rect 316614 207922 316682 207978
rect 316738 207922 316806 207978
rect 316862 207922 347154 207978
rect 347210 207922 347278 207978
rect 347334 207922 347402 207978
rect 347458 207922 347526 207978
rect 347582 207922 377874 207978
rect 377930 207922 377998 207978
rect 378054 207922 378122 207978
rect 378178 207922 378246 207978
rect 378302 207922 408594 207978
rect 408650 207922 408718 207978
rect 408774 207922 408842 207978
rect 408898 207922 408966 207978
rect 409022 207922 439314 207978
rect 439370 207922 439438 207978
rect 439494 207922 439562 207978
rect 439618 207922 439686 207978
rect 439742 207922 470034 207978
rect 470090 207922 470158 207978
rect 470214 207922 470282 207978
rect 470338 207922 470406 207978
rect 470462 207922 489822 207978
rect 489878 207922 489946 207978
rect 490002 207922 498390 207978
rect 498446 207922 498514 207978
rect 498570 207922 506958 207978
rect 507014 207922 507082 207978
rect 507138 207922 515526 207978
rect 515582 207922 515650 207978
rect 515706 207922 531474 207978
rect 531530 207922 531598 207978
rect 531654 207922 531722 207978
rect 531778 207922 531846 207978
rect 531902 207922 562194 207978
rect 562250 207922 562318 207978
rect 562374 207922 562442 207978
rect 562498 207922 562566 207978
rect 562622 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect -1916 207826 597980 207922
rect 4156 206578 50388 206594
rect 4156 206522 4172 206578
rect 4228 206522 50316 206578
rect 50372 206522 50388 206578
rect 4156 206506 50388 206522
rect -1916 202350 597980 202446
rect -1916 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 36234 202350
rect 36290 202294 36358 202350
rect 36414 202294 36482 202350
rect 36538 202294 36606 202350
rect 36662 202294 44518 202350
rect 44574 202294 44642 202350
rect 44698 202294 75238 202350
rect 75294 202294 75362 202350
rect 75418 202294 105958 202350
rect 106014 202294 106082 202350
rect 106138 202294 136678 202350
rect 136734 202294 136802 202350
rect 136858 202294 167398 202350
rect 167454 202294 167522 202350
rect 167578 202294 198118 202350
rect 198174 202294 198242 202350
rect 198298 202294 228838 202350
rect 228894 202294 228962 202350
rect 229018 202294 259558 202350
rect 259614 202294 259682 202350
rect 259738 202294 281994 202350
rect 282050 202294 282118 202350
rect 282174 202294 282242 202350
rect 282298 202294 282366 202350
rect 282422 202294 312714 202350
rect 312770 202294 312838 202350
rect 312894 202294 312962 202350
rect 313018 202294 313086 202350
rect 313142 202294 343434 202350
rect 343490 202294 343558 202350
rect 343614 202294 343682 202350
rect 343738 202294 343806 202350
rect 343862 202294 374154 202350
rect 374210 202294 374278 202350
rect 374334 202294 374402 202350
rect 374458 202294 374526 202350
rect 374582 202294 404874 202350
rect 404930 202294 404998 202350
rect 405054 202294 405122 202350
rect 405178 202294 405246 202350
rect 405302 202294 435594 202350
rect 435650 202294 435718 202350
rect 435774 202294 435842 202350
rect 435898 202294 435966 202350
rect 436022 202294 466314 202350
rect 466370 202294 466438 202350
rect 466494 202294 466562 202350
rect 466618 202294 466686 202350
rect 466742 202294 497034 202350
rect 497090 202294 497158 202350
rect 497214 202294 497282 202350
rect 497338 202294 497406 202350
rect 497462 202294 527754 202350
rect 527810 202294 527878 202350
rect 527934 202294 528002 202350
rect 528058 202294 528126 202350
rect 528182 202294 558474 202350
rect 558530 202294 558598 202350
rect 558654 202294 558722 202350
rect 558778 202294 558846 202350
rect 558902 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597980 202350
rect -1916 202226 597980 202294
rect -1916 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 36234 202226
rect 36290 202170 36358 202226
rect 36414 202170 36482 202226
rect 36538 202170 36606 202226
rect 36662 202170 44518 202226
rect 44574 202170 44642 202226
rect 44698 202170 75238 202226
rect 75294 202170 75362 202226
rect 75418 202170 105958 202226
rect 106014 202170 106082 202226
rect 106138 202170 136678 202226
rect 136734 202170 136802 202226
rect 136858 202170 167398 202226
rect 167454 202170 167522 202226
rect 167578 202170 198118 202226
rect 198174 202170 198242 202226
rect 198298 202170 228838 202226
rect 228894 202170 228962 202226
rect 229018 202170 259558 202226
rect 259614 202170 259682 202226
rect 259738 202170 281994 202226
rect 282050 202170 282118 202226
rect 282174 202170 282242 202226
rect 282298 202170 282366 202226
rect 282422 202170 312714 202226
rect 312770 202170 312838 202226
rect 312894 202170 312962 202226
rect 313018 202170 313086 202226
rect 313142 202170 343434 202226
rect 343490 202170 343558 202226
rect 343614 202170 343682 202226
rect 343738 202170 343806 202226
rect 343862 202170 374154 202226
rect 374210 202170 374278 202226
rect 374334 202170 374402 202226
rect 374458 202170 374526 202226
rect 374582 202170 404874 202226
rect 404930 202170 404998 202226
rect 405054 202170 405122 202226
rect 405178 202170 405246 202226
rect 405302 202170 435594 202226
rect 435650 202170 435718 202226
rect 435774 202170 435842 202226
rect 435898 202170 435966 202226
rect 436022 202170 466314 202226
rect 466370 202170 466438 202226
rect 466494 202170 466562 202226
rect 466618 202170 466686 202226
rect 466742 202170 497034 202226
rect 497090 202170 497158 202226
rect 497214 202170 497282 202226
rect 497338 202170 497406 202226
rect 497462 202170 527754 202226
rect 527810 202170 527878 202226
rect 527934 202170 528002 202226
rect 528058 202170 528126 202226
rect 528182 202170 558474 202226
rect 558530 202170 558598 202226
rect 558654 202170 558722 202226
rect 558778 202170 558846 202226
rect 558902 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597980 202226
rect -1916 202102 597980 202170
rect -1916 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 36234 202102
rect 36290 202046 36358 202102
rect 36414 202046 36482 202102
rect 36538 202046 36606 202102
rect 36662 202046 44518 202102
rect 44574 202046 44642 202102
rect 44698 202046 75238 202102
rect 75294 202046 75362 202102
rect 75418 202046 105958 202102
rect 106014 202046 106082 202102
rect 106138 202046 136678 202102
rect 136734 202046 136802 202102
rect 136858 202046 167398 202102
rect 167454 202046 167522 202102
rect 167578 202046 198118 202102
rect 198174 202046 198242 202102
rect 198298 202046 228838 202102
rect 228894 202046 228962 202102
rect 229018 202046 259558 202102
rect 259614 202046 259682 202102
rect 259738 202046 281994 202102
rect 282050 202046 282118 202102
rect 282174 202046 282242 202102
rect 282298 202046 282366 202102
rect 282422 202046 312714 202102
rect 312770 202046 312838 202102
rect 312894 202046 312962 202102
rect 313018 202046 313086 202102
rect 313142 202046 343434 202102
rect 343490 202046 343558 202102
rect 343614 202046 343682 202102
rect 343738 202046 343806 202102
rect 343862 202046 374154 202102
rect 374210 202046 374278 202102
rect 374334 202046 374402 202102
rect 374458 202046 374526 202102
rect 374582 202046 404874 202102
rect 404930 202046 404998 202102
rect 405054 202046 405122 202102
rect 405178 202046 405246 202102
rect 405302 202046 435594 202102
rect 435650 202046 435718 202102
rect 435774 202046 435842 202102
rect 435898 202046 435966 202102
rect 436022 202046 466314 202102
rect 466370 202046 466438 202102
rect 466494 202046 466562 202102
rect 466618 202046 466686 202102
rect 466742 202046 497034 202102
rect 497090 202046 497158 202102
rect 497214 202046 497282 202102
rect 497338 202046 497406 202102
rect 497462 202046 527754 202102
rect 527810 202046 527878 202102
rect 527934 202046 528002 202102
rect 528058 202046 528126 202102
rect 528182 202046 558474 202102
rect 558530 202046 558598 202102
rect 558654 202046 558722 202102
rect 558778 202046 558846 202102
rect 558902 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597980 202102
rect -1916 201978 597980 202046
rect -1916 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 36234 201978
rect 36290 201922 36358 201978
rect 36414 201922 36482 201978
rect 36538 201922 36606 201978
rect 36662 201922 44518 201978
rect 44574 201922 44642 201978
rect 44698 201922 75238 201978
rect 75294 201922 75362 201978
rect 75418 201922 105958 201978
rect 106014 201922 106082 201978
rect 106138 201922 136678 201978
rect 136734 201922 136802 201978
rect 136858 201922 167398 201978
rect 167454 201922 167522 201978
rect 167578 201922 198118 201978
rect 198174 201922 198242 201978
rect 198298 201922 228838 201978
rect 228894 201922 228962 201978
rect 229018 201922 259558 201978
rect 259614 201922 259682 201978
rect 259738 201922 281994 201978
rect 282050 201922 282118 201978
rect 282174 201922 282242 201978
rect 282298 201922 282366 201978
rect 282422 201922 312714 201978
rect 312770 201922 312838 201978
rect 312894 201922 312962 201978
rect 313018 201922 313086 201978
rect 313142 201922 343434 201978
rect 343490 201922 343558 201978
rect 343614 201922 343682 201978
rect 343738 201922 343806 201978
rect 343862 201922 374154 201978
rect 374210 201922 374278 201978
rect 374334 201922 374402 201978
rect 374458 201922 374526 201978
rect 374582 201922 404874 201978
rect 404930 201922 404998 201978
rect 405054 201922 405122 201978
rect 405178 201922 405246 201978
rect 405302 201922 435594 201978
rect 435650 201922 435718 201978
rect 435774 201922 435842 201978
rect 435898 201922 435966 201978
rect 436022 201922 466314 201978
rect 466370 201922 466438 201978
rect 466494 201922 466562 201978
rect 466618 201922 466686 201978
rect 466742 201922 497034 201978
rect 497090 201922 497158 201978
rect 497214 201922 497282 201978
rect 497338 201922 497406 201978
rect 497462 201922 527754 201978
rect 527810 201922 527878 201978
rect 527934 201922 528002 201978
rect 528058 201922 528126 201978
rect 528182 201922 558474 201978
rect 558530 201922 558598 201978
rect 558654 201922 558722 201978
rect 558778 201922 558846 201978
rect 558902 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597980 201978
rect -1916 201826 597980 201922
rect 464476 198118 497716 198134
rect 464476 198062 464492 198118
rect 464548 198062 497644 198118
rect 497700 198062 497716 198118
rect 464476 198046 497716 198062
rect 476236 197938 499172 197954
rect 476236 197882 476252 197938
rect 476308 197882 499100 197938
rect 499156 197882 499172 197938
rect 476236 197866 499172 197882
rect 479596 197758 502308 197774
rect 479596 197702 479612 197758
rect 479668 197702 502236 197758
rect 502292 197702 502308 197758
rect 479596 197686 502308 197702
rect -1916 190350 597980 190446
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 9234 190350
rect 9290 190294 9358 190350
rect 9414 190294 9482 190350
rect 9538 190294 9606 190350
rect 9662 190294 39954 190350
rect 40010 190294 40078 190350
rect 40134 190294 40202 190350
rect 40258 190294 40326 190350
rect 40382 190294 59878 190350
rect 59934 190294 60002 190350
rect 60058 190294 90598 190350
rect 90654 190294 90722 190350
rect 90778 190294 121318 190350
rect 121374 190294 121442 190350
rect 121498 190294 152038 190350
rect 152094 190294 152162 190350
rect 152218 190294 182758 190350
rect 182814 190294 182882 190350
rect 182938 190294 213478 190350
rect 213534 190294 213602 190350
rect 213658 190294 244198 190350
rect 244254 190294 244322 190350
rect 244378 190294 285714 190350
rect 285770 190294 285838 190350
rect 285894 190294 285962 190350
rect 286018 190294 286086 190350
rect 286142 190294 316434 190350
rect 316490 190294 316558 190350
rect 316614 190294 316682 190350
rect 316738 190294 316806 190350
rect 316862 190294 347154 190350
rect 347210 190294 347278 190350
rect 347334 190294 347402 190350
rect 347458 190294 347526 190350
rect 347582 190294 377874 190350
rect 377930 190294 377998 190350
rect 378054 190294 378122 190350
rect 378178 190294 378246 190350
rect 378302 190294 408594 190350
rect 408650 190294 408718 190350
rect 408774 190294 408842 190350
rect 408898 190294 408966 190350
rect 409022 190294 439314 190350
rect 439370 190294 439438 190350
rect 439494 190294 439562 190350
rect 439618 190294 439686 190350
rect 439742 190294 470034 190350
rect 470090 190294 470158 190350
rect 470214 190294 470282 190350
rect 470338 190294 470406 190350
rect 470462 190294 500754 190350
rect 500810 190294 500878 190350
rect 500934 190294 501002 190350
rect 501058 190294 501126 190350
rect 501182 190294 531474 190350
rect 531530 190294 531598 190350
rect 531654 190294 531722 190350
rect 531778 190294 531846 190350
rect 531902 190294 562194 190350
rect 562250 190294 562318 190350
rect 562374 190294 562442 190350
rect 562498 190294 562566 190350
rect 562622 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect -1916 190226 597980 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 9234 190226
rect 9290 190170 9358 190226
rect 9414 190170 9482 190226
rect 9538 190170 9606 190226
rect 9662 190170 39954 190226
rect 40010 190170 40078 190226
rect 40134 190170 40202 190226
rect 40258 190170 40326 190226
rect 40382 190170 59878 190226
rect 59934 190170 60002 190226
rect 60058 190170 90598 190226
rect 90654 190170 90722 190226
rect 90778 190170 121318 190226
rect 121374 190170 121442 190226
rect 121498 190170 152038 190226
rect 152094 190170 152162 190226
rect 152218 190170 182758 190226
rect 182814 190170 182882 190226
rect 182938 190170 213478 190226
rect 213534 190170 213602 190226
rect 213658 190170 244198 190226
rect 244254 190170 244322 190226
rect 244378 190170 285714 190226
rect 285770 190170 285838 190226
rect 285894 190170 285962 190226
rect 286018 190170 286086 190226
rect 286142 190170 316434 190226
rect 316490 190170 316558 190226
rect 316614 190170 316682 190226
rect 316738 190170 316806 190226
rect 316862 190170 347154 190226
rect 347210 190170 347278 190226
rect 347334 190170 347402 190226
rect 347458 190170 347526 190226
rect 347582 190170 377874 190226
rect 377930 190170 377998 190226
rect 378054 190170 378122 190226
rect 378178 190170 378246 190226
rect 378302 190170 408594 190226
rect 408650 190170 408718 190226
rect 408774 190170 408842 190226
rect 408898 190170 408966 190226
rect 409022 190170 439314 190226
rect 439370 190170 439438 190226
rect 439494 190170 439562 190226
rect 439618 190170 439686 190226
rect 439742 190170 470034 190226
rect 470090 190170 470158 190226
rect 470214 190170 470282 190226
rect 470338 190170 470406 190226
rect 470462 190170 500754 190226
rect 500810 190170 500878 190226
rect 500934 190170 501002 190226
rect 501058 190170 501126 190226
rect 501182 190170 531474 190226
rect 531530 190170 531598 190226
rect 531654 190170 531722 190226
rect 531778 190170 531846 190226
rect 531902 190170 562194 190226
rect 562250 190170 562318 190226
rect 562374 190170 562442 190226
rect 562498 190170 562566 190226
rect 562622 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect -1916 190102 597980 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 9234 190102
rect 9290 190046 9358 190102
rect 9414 190046 9482 190102
rect 9538 190046 9606 190102
rect 9662 190046 39954 190102
rect 40010 190046 40078 190102
rect 40134 190046 40202 190102
rect 40258 190046 40326 190102
rect 40382 190046 59878 190102
rect 59934 190046 60002 190102
rect 60058 190046 90598 190102
rect 90654 190046 90722 190102
rect 90778 190046 121318 190102
rect 121374 190046 121442 190102
rect 121498 190046 152038 190102
rect 152094 190046 152162 190102
rect 152218 190046 182758 190102
rect 182814 190046 182882 190102
rect 182938 190046 213478 190102
rect 213534 190046 213602 190102
rect 213658 190046 244198 190102
rect 244254 190046 244322 190102
rect 244378 190046 285714 190102
rect 285770 190046 285838 190102
rect 285894 190046 285962 190102
rect 286018 190046 286086 190102
rect 286142 190046 316434 190102
rect 316490 190046 316558 190102
rect 316614 190046 316682 190102
rect 316738 190046 316806 190102
rect 316862 190046 347154 190102
rect 347210 190046 347278 190102
rect 347334 190046 347402 190102
rect 347458 190046 347526 190102
rect 347582 190046 377874 190102
rect 377930 190046 377998 190102
rect 378054 190046 378122 190102
rect 378178 190046 378246 190102
rect 378302 190046 408594 190102
rect 408650 190046 408718 190102
rect 408774 190046 408842 190102
rect 408898 190046 408966 190102
rect 409022 190046 439314 190102
rect 439370 190046 439438 190102
rect 439494 190046 439562 190102
rect 439618 190046 439686 190102
rect 439742 190046 470034 190102
rect 470090 190046 470158 190102
rect 470214 190046 470282 190102
rect 470338 190046 470406 190102
rect 470462 190046 500754 190102
rect 500810 190046 500878 190102
rect 500934 190046 501002 190102
rect 501058 190046 501126 190102
rect 501182 190046 531474 190102
rect 531530 190046 531598 190102
rect 531654 190046 531722 190102
rect 531778 190046 531846 190102
rect 531902 190046 562194 190102
rect 562250 190046 562318 190102
rect 562374 190046 562442 190102
rect 562498 190046 562566 190102
rect 562622 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect -1916 189978 597980 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 9234 189978
rect 9290 189922 9358 189978
rect 9414 189922 9482 189978
rect 9538 189922 9606 189978
rect 9662 189922 39954 189978
rect 40010 189922 40078 189978
rect 40134 189922 40202 189978
rect 40258 189922 40326 189978
rect 40382 189922 59878 189978
rect 59934 189922 60002 189978
rect 60058 189922 90598 189978
rect 90654 189922 90722 189978
rect 90778 189922 121318 189978
rect 121374 189922 121442 189978
rect 121498 189922 152038 189978
rect 152094 189922 152162 189978
rect 152218 189922 182758 189978
rect 182814 189922 182882 189978
rect 182938 189922 213478 189978
rect 213534 189922 213602 189978
rect 213658 189922 244198 189978
rect 244254 189922 244322 189978
rect 244378 189922 285714 189978
rect 285770 189922 285838 189978
rect 285894 189922 285962 189978
rect 286018 189922 286086 189978
rect 286142 189922 316434 189978
rect 316490 189922 316558 189978
rect 316614 189922 316682 189978
rect 316738 189922 316806 189978
rect 316862 189922 347154 189978
rect 347210 189922 347278 189978
rect 347334 189922 347402 189978
rect 347458 189922 347526 189978
rect 347582 189922 377874 189978
rect 377930 189922 377998 189978
rect 378054 189922 378122 189978
rect 378178 189922 378246 189978
rect 378302 189922 408594 189978
rect 408650 189922 408718 189978
rect 408774 189922 408842 189978
rect 408898 189922 408966 189978
rect 409022 189922 439314 189978
rect 439370 189922 439438 189978
rect 439494 189922 439562 189978
rect 439618 189922 439686 189978
rect 439742 189922 470034 189978
rect 470090 189922 470158 189978
rect 470214 189922 470282 189978
rect 470338 189922 470406 189978
rect 470462 189922 500754 189978
rect 500810 189922 500878 189978
rect 500934 189922 501002 189978
rect 501058 189922 501126 189978
rect 501182 189922 531474 189978
rect 531530 189922 531598 189978
rect 531654 189922 531722 189978
rect 531778 189922 531846 189978
rect 531902 189922 562194 189978
rect 562250 189922 562318 189978
rect 562374 189922 562442 189978
rect 562498 189922 562566 189978
rect 562622 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect -1916 189826 597980 189922
rect -1916 184350 597980 184446
rect -1916 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 36234 184350
rect 36290 184294 36358 184350
rect 36414 184294 36482 184350
rect 36538 184294 36606 184350
rect 36662 184294 44518 184350
rect 44574 184294 44642 184350
rect 44698 184294 75238 184350
rect 75294 184294 75362 184350
rect 75418 184294 105958 184350
rect 106014 184294 106082 184350
rect 106138 184294 136678 184350
rect 136734 184294 136802 184350
rect 136858 184294 167398 184350
rect 167454 184294 167522 184350
rect 167578 184294 198118 184350
rect 198174 184294 198242 184350
rect 198298 184294 228838 184350
rect 228894 184294 228962 184350
rect 229018 184294 259558 184350
rect 259614 184294 259682 184350
rect 259738 184294 281994 184350
rect 282050 184294 282118 184350
rect 282174 184294 282242 184350
rect 282298 184294 282366 184350
rect 282422 184294 312714 184350
rect 312770 184294 312838 184350
rect 312894 184294 312962 184350
rect 313018 184294 313086 184350
rect 313142 184294 343434 184350
rect 343490 184294 343558 184350
rect 343614 184294 343682 184350
rect 343738 184294 343806 184350
rect 343862 184294 374154 184350
rect 374210 184294 374278 184350
rect 374334 184294 374402 184350
rect 374458 184294 374526 184350
rect 374582 184294 404874 184350
rect 404930 184294 404998 184350
rect 405054 184294 405122 184350
rect 405178 184294 405246 184350
rect 405302 184294 435594 184350
rect 435650 184294 435718 184350
rect 435774 184294 435842 184350
rect 435898 184294 435966 184350
rect 436022 184294 466314 184350
rect 466370 184294 466438 184350
rect 466494 184294 466562 184350
rect 466618 184294 466686 184350
rect 466742 184294 497034 184350
rect 497090 184294 497158 184350
rect 497214 184294 497282 184350
rect 497338 184294 497406 184350
rect 497462 184294 527754 184350
rect 527810 184294 527878 184350
rect 527934 184294 528002 184350
rect 528058 184294 528126 184350
rect 528182 184294 558474 184350
rect 558530 184294 558598 184350
rect 558654 184294 558722 184350
rect 558778 184294 558846 184350
rect 558902 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597980 184350
rect -1916 184226 597980 184294
rect -1916 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 36234 184226
rect 36290 184170 36358 184226
rect 36414 184170 36482 184226
rect 36538 184170 36606 184226
rect 36662 184170 44518 184226
rect 44574 184170 44642 184226
rect 44698 184170 75238 184226
rect 75294 184170 75362 184226
rect 75418 184170 105958 184226
rect 106014 184170 106082 184226
rect 106138 184170 136678 184226
rect 136734 184170 136802 184226
rect 136858 184170 167398 184226
rect 167454 184170 167522 184226
rect 167578 184170 198118 184226
rect 198174 184170 198242 184226
rect 198298 184170 228838 184226
rect 228894 184170 228962 184226
rect 229018 184170 259558 184226
rect 259614 184170 259682 184226
rect 259738 184170 281994 184226
rect 282050 184170 282118 184226
rect 282174 184170 282242 184226
rect 282298 184170 282366 184226
rect 282422 184170 312714 184226
rect 312770 184170 312838 184226
rect 312894 184170 312962 184226
rect 313018 184170 313086 184226
rect 313142 184170 343434 184226
rect 343490 184170 343558 184226
rect 343614 184170 343682 184226
rect 343738 184170 343806 184226
rect 343862 184170 374154 184226
rect 374210 184170 374278 184226
rect 374334 184170 374402 184226
rect 374458 184170 374526 184226
rect 374582 184170 404874 184226
rect 404930 184170 404998 184226
rect 405054 184170 405122 184226
rect 405178 184170 405246 184226
rect 405302 184170 435594 184226
rect 435650 184170 435718 184226
rect 435774 184170 435842 184226
rect 435898 184170 435966 184226
rect 436022 184170 466314 184226
rect 466370 184170 466438 184226
rect 466494 184170 466562 184226
rect 466618 184170 466686 184226
rect 466742 184170 497034 184226
rect 497090 184170 497158 184226
rect 497214 184170 497282 184226
rect 497338 184170 497406 184226
rect 497462 184170 527754 184226
rect 527810 184170 527878 184226
rect 527934 184170 528002 184226
rect 528058 184170 528126 184226
rect 528182 184170 558474 184226
rect 558530 184170 558598 184226
rect 558654 184170 558722 184226
rect 558778 184170 558846 184226
rect 558902 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597980 184226
rect -1916 184102 597980 184170
rect -1916 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 36234 184102
rect 36290 184046 36358 184102
rect 36414 184046 36482 184102
rect 36538 184046 36606 184102
rect 36662 184046 44518 184102
rect 44574 184046 44642 184102
rect 44698 184046 75238 184102
rect 75294 184046 75362 184102
rect 75418 184046 105958 184102
rect 106014 184046 106082 184102
rect 106138 184046 136678 184102
rect 136734 184046 136802 184102
rect 136858 184046 167398 184102
rect 167454 184046 167522 184102
rect 167578 184046 198118 184102
rect 198174 184046 198242 184102
rect 198298 184046 228838 184102
rect 228894 184046 228962 184102
rect 229018 184046 259558 184102
rect 259614 184046 259682 184102
rect 259738 184046 281994 184102
rect 282050 184046 282118 184102
rect 282174 184046 282242 184102
rect 282298 184046 282366 184102
rect 282422 184046 312714 184102
rect 312770 184046 312838 184102
rect 312894 184046 312962 184102
rect 313018 184046 313086 184102
rect 313142 184046 343434 184102
rect 343490 184046 343558 184102
rect 343614 184046 343682 184102
rect 343738 184046 343806 184102
rect 343862 184046 374154 184102
rect 374210 184046 374278 184102
rect 374334 184046 374402 184102
rect 374458 184046 374526 184102
rect 374582 184046 404874 184102
rect 404930 184046 404998 184102
rect 405054 184046 405122 184102
rect 405178 184046 405246 184102
rect 405302 184046 435594 184102
rect 435650 184046 435718 184102
rect 435774 184046 435842 184102
rect 435898 184046 435966 184102
rect 436022 184046 466314 184102
rect 466370 184046 466438 184102
rect 466494 184046 466562 184102
rect 466618 184046 466686 184102
rect 466742 184046 497034 184102
rect 497090 184046 497158 184102
rect 497214 184046 497282 184102
rect 497338 184046 497406 184102
rect 497462 184046 527754 184102
rect 527810 184046 527878 184102
rect 527934 184046 528002 184102
rect 528058 184046 528126 184102
rect 528182 184046 558474 184102
rect 558530 184046 558598 184102
rect 558654 184046 558722 184102
rect 558778 184046 558846 184102
rect 558902 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597980 184102
rect -1916 183978 597980 184046
rect -1916 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 36234 183978
rect 36290 183922 36358 183978
rect 36414 183922 36482 183978
rect 36538 183922 36606 183978
rect 36662 183922 44518 183978
rect 44574 183922 44642 183978
rect 44698 183922 75238 183978
rect 75294 183922 75362 183978
rect 75418 183922 105958 183978
rect 106014 183922 106082 183978
rect 106138 183922 136678 183978
rect 136734 183922 136802 183978
rect 136858 183922 167398 183978
rect 167454 183922 167522 183978
rect 167578 183922 198118 183978
rect 198174 183922 198242 183978
rect 198298 183922 228838 183978
rect 228894 183922 228962 183978
rect 229018 183922 259558 183978
rect 259614 183922 259682 183978
rect 259738 183922 281994 183978
rect 282050 183922 282118 183978
rect 282174 183922 282242 183978
rect 282298 183922 282366 183978
rect 282422 183922 312714 183978
rect 312770 183922 312838 183978
rect 312894 183922 312962 183978
rect 313018 183922 313086 183978
rect 313142 183922 343434 183978
rect 343490 183922 343558 183978
rect 343614 183922 343682 183978
rect 343738 183922 343806 183978
rect 343862 183922 374154 183978
rect 374210 183922 374278 183978
rect 374334 183922 374402 183978
rect 374458 183922 374526 183978
rect 374582 183922 404874 183978
rect 404930 183922 404998 183978
rect 405054 183922 405122 183978
rect 405178 183922 405246 183978
rect 405302 183922 435594 183978
rect 435650 183922 435718 183978
rect 435774 183922 435842 183978
rect 435898 183922 435966 183978
rect 436022 183922 466314 183978
rect 466370 183922 466438 183978
rect 466494 183922 466562 183978
rect 466618 183922 466686 183978
rect 466742 183922 497034 183978
rect 497090 183922 497158 183978
rect 497214 183922 497282 183978
rect 497338 183922 497406 183978
rect 497462 183922 527754 183978
rect 527810 183922 527878 183978
rect 527934 183922 528002 183978
rect 528058 183922 528126 183978
rect 528182 183922 558474 183978
rect 558530 183922 558598 183978
rect 558654 183922 558722 183978
rect 558778 183922 558846 183978
rect 558902 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597980 183978
rect -1916 183826 597980 183922
rect -1916 172350 597980 172446
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 9234 172350
rect 9290 172294 9358 172350
rect 9414 172294 9482 172350
rect 9538 172294 9606 172350
rect 9662 172294 39954 172350
rect 40010 172294 40078 172350
rect 40134 172294 40202 172350
rect 40258 172294 40326 172350
rect 40382 172294 59878 172350
rect 59934 172294 60002 172350
rect 60058 172294 90598 172350
rect 90654 172294 90722 172350
rect 90778 172294 121318 172350
rect 121374 172294 121442 172350
rect 121498 172294 152038 172350
rect 152094 172294 152162 172350
rect 152218 172294 182758 172350
rect 182814 172294 182882 172350
rect 182938 172294 213478 172350
rect 213534 172294 213602 172350
rect 213658 172294 244198 172350
rect 244254 172294 244322 172350
rect 244378 172294 285714 172350
rect 285770 172294 285838 172350
rect 285894 172294 285962 172350
rect 286018 172294 286086 172350
rect 286142 172294 316434 172350
rect 316490 172294 316558 172350
rect 316614 172294 316682 172350
rect 316738 172294 316806 172350
rect 316862 172294 347154 172350
rect 347210 172294 347278 172350
rect 347334 172294 347402 172350
rect 347458 172294 347526 172350
rect 347582 172294 377874 172350
rect 377930 172294 377998 172350
rect 378054 172294 378122 172350
rect 378178 172294 378246 172350
rect 378302 172294 408594 172350
rect 408650 172294 408718 172350
rect 408774 172294 408842 172350
rect 408898 172294 408966 172350
rect 409022 172294 439314 172350
rect 439370 172294 439438 172350
rect 439494 172294 439562 172350
rect 439618 172294 439686 172350
rect 439742 172294 470034 172350
rect 470090 172294 470158 172350
rect 470214 172294 470282 172350
rect 470338 172294 470406 172350
rect 470462 172294 500754 172350
rect 500810 172294 500878 172350
rect 500934 172294 501002 172350
rect 501058 172294 501126 172350
rect 501182 172294 531474 172350
rect 531530 172294 531598 172350
rect 531654 172294 531722 172350
rect 531778 172294 531846 172350
rect 531902 172294 562194 172350
rect 562250 172294 562318 172350
rect 562374 172294 562442 172350
rect 562498 172294 562566 172350
rect 562622 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect -1916 172226 597980 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 9234 172226
rect 9290 172170 9358 172226
rect 9414 172170 9482 172226
rect 9538 172170 9606 172226
rect 9662 172170 39954 172226
rect 40010 172170 40078 172226
rect 40134 172170 40202 172226
rect 40258 172170 40326 172226
rect 40382 172170 59878 172226
rect 59934 172170 60002 172226
rect 60058 172170 90598 172226
rect 90654 172170 90722 172226
rect 90778 172170 121318 172226
rect 121374 172170 121442 172226
rect 121498 172170 152038 172226
rect 152094 172170 152162 172226
rect 152218 172170 182758 172226
rect 182814 172170 182882 172226
rect 182938 172170 213478 172226
rect 213534 172170 213602 172226
rect 213658 172170 244198 172226
rect 244254 172170 244322 172226
rect 244378 172170 285714 172226
rect 285770 172170 285838 172226
rect 285894 172170 285962 172226
rect 286018 172170 286086 172226
rect 286142 172170 316434 172226
rect 316490 172170 316558 172226
rect 316614 172170 316682 172226
rect 316738 172170 316806 172226
rect 316862 172170 347154 172226
rect 347210 172170 347278 172226
rect 347334 172170 347402 172226
rect 347458 172170 347526 172226
rect 347582 172170 377874 172226
rect 377930 172170 377998 172226
rect 378054 172170 378122 172226
rect 378178 172170 378246 172226
rect 378302 172170 408594 172226
rect 408650 172170 408718 172226
rect 408774 172170 408842 172226
rect 408898 172170 408966 172226
rect 409022 172170 439314 172226
rect 439370 172170 439438 172226
rect 439494 172170 439562 172226
rect 439618 172170 439686 172226
rect 439742 172170 470034 172226
rect 470090 172170 470158 172226
rect 470214 172170 470282 172226
rect 470338 172170 470406 172226
rect 470462 172170 500754 172226
rect 500810 172170 500878 172226
rect 500934 172170 501002 172226
rect 501058 172170 501126 172226
rect 501182 172170 531474 172226
rect 531530 172170 531598 172226
rect 531654 172170 531722 172226
rect 531778 172170 531846 172226
rect 531902 172170 562194 172226
rect 562250 172170 562318 172226
rect 562374 172170 562442 172226
rect 562498 172170 562566 172226
rect 562622 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect -1916 172102 597980 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 9234 172102
rect 9290 172046 9358 172102
rect 9414 172046 9482 172102
rect 9538 172046 9606 172102
rect 9662 172046 39954 172102
rect 40010 172046 40078 172102
rect 40134 172046 40202 172102
rect 40258 172046 40326 172102
rect 40382 172046 59878 172102
rect 59934 172046 60002 172102
rect 60058 172046 90598 172102
rect 90654 172046 90722 172102
rect 90778 172046 121318 172102
rect 121374 172046 121442 172102
rect 121498 172046 152038 172102
rect 152094 172046 152162 172102
rect 152218 172046 182758 172102
rect 182814 172046 182882 172102
rect 182938 172046 213478 172102
rect 213534 172046 213602 172102
rect 213658 172046 244198 172102
rect 244254 172046 244322 172102
rect 244378 172046 285714 172102
rect 285770 172046 285838 172102
rect 285894 172046 285962 172102
rect 286018 172046 286086 172102
rect 286142 172046 316434 172102
rect 316490 172046 316558 172102
rect 316614 172046 316682 172102
rect 316738 172046 316806 172102
rect 316862 172046 347154 172102
rect 347210 172046 347278 172102
rect 347334 172046 347402 172102
rect 347458 172046 347526 172102
rect 347582 172046 377874 172102
rect 377930 172046 377998 172102
rect 378054 172046 378122 172102
rect 378178 172046 378246 172102
rect 378302 172046 408594 172102
rect 408650 172046 408718 172102
rect 408774 172046 408842 172102
rect 408898 172046 408966 172102
rect 409022 172046 439314 172102
rect 439370 172046 439438 172102
rect 439494 172046 439562 172102
rect 439618 172046 439686 172102
rect 439742 172046 470034 172102
rect 470090 172046 470158 172102
rect 470214 172046 470282 172102
rect 470338 172046 470406 172102
rect 470462 172046 500754 172102
rect 500810 172046 500878 172102
rect 500934 172046 501002 172102
rect 501058 172046 501126 172102
rect 501182 172046 531474 172102
rect 531530 172046 531598 172102
rect 531654 172046 531722 172102
rect 531778 172046 531846 172102
rect 531902 172046 562194 172102
rect 562250 172046 562318 172102
rect 562374 172046 562442 172102
rect 562498 172046 562566 172102
rect 562622 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect -1916 171978 597980 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 9234 171978
rect 9290 171922 9358 171978
rect 9414 171922 9482 171978
rect 9538 171922 9606 171978
rect 9662 171922 39954 171978
rect 40010 171922 40078 171978
rect 40134 171922 40202 171978
rect 40258 171922 40326 171978
rect 40382 171922 59878 171978
rect 59934 171922 60002 171978
rect 60058 171922 90598 171978
rect 90654 171922 90722 171978
rect 90778 171922 121318 171978
rect 121374 171922 121442 171978
rect 121498 171922 152038 171978
rect 152094 171922 152162 171978
rect 152218 171922 182758 171978
rect 182814 171922 182882 171978
rect 182938 171922 213478 171978
rect 213534 171922 213602 171978
rect 213658 171922 244198 171978
rect 244254 171922 244322 171978
rect 244378 171922 285714 171978
rect 285770 171922 285838 171978
rect 285894 171922 285962 171978
rect 286018 171922 286086 171978
rect 286142 171922 316434 171978
rect 316490 171922 316558 171978
rect 316614 171922 316682 171978
rect 316738 171922 316806 171978
rect 316862 171922 347154 171978
rect 347210 171922 347278 171978
rect 347334 171922 347402 171978
rect 347458 171922 347526 171978
rect 347582 171922 377874 171978
rect 377930 171922 377998 171978
rect 378054 171922 378122 171978
rect 378178 171922 378246 171978
rect 378302 171922 408594 171978
rect 408650 171922 408718 171978
rect 408774 171922 408842 171978
rect 408898 171922 408966 171978
rect 409022 171922 439314 171978
rect 439370 171922 439438 171978
rect 439494 171922 439562 171978
rect 439618 171922 439686 171978
rect 439742 171922 470034 171978
rect 470090 171922 470158 171978
rect 470214 171922 470282 171978
rect 470338 171922 470406 171978
rect 470462 171922 500754 171978
rect 500810 171922 500878 171978
rect 500934 171922 501002 171978
rect 501058 171922 501126 171978
rect 501182 171922 531474 171978
rect 531530 171922 531598 171978
rect 531654 171922 531722 171978
rect 531778 171922 531846 171978
rect 531902 171922 562194 171978
rect 562250 171922 562318 171978
rect 562374 171922 562442 171978
rect 562498 171922 562566 171978
rect 562622 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect -1916 171826 597980 171922
rect -1916 166350 597980 166446
rect -1916 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 36234 166350
rect 36290 166294 36358 166350
rect 36414 166294 36482 166350
rect 36538 166294 36606 166350
rect 36662 166294 44518 166350
rect 44574 166294 44642 166350
rect 44698 166294 75238 166350
rect 75294 166294 75362 166350
rect 75418 166294 105958 166350
rect 106014 166294 106082 166350
rect 106138 166294 136678 166350
rect 136734 166294 136802 166350
rect 136858 166294 167398 166350
rect 167454 166294 167522 166350
rect 167578 166294 198118 166350
rect 198174 166294 198242 166350
rect 198298 166294 228838 166350
rect 228894 166294 228962 166350
rect 229018 166294 259558 166350
rect 259614 166294 259682 166350
rect 259738 166294 281994 166350
rect 282050 166294 282118 166350
rect 282174 166294 282242 166350
rect 282298 166294 282366 166350
rect 282422 166294 312714 166350
rect 312770 166294 312838 166350
rect 312894 166294 312962 166350
rect 313018 166294 313086 166350
rect 313142 166294 343434 166350
rect 343490 166294 343558 166350
rect 343614 166294 343682 166350
rect 343738 166294 343806 166350
rect 343862 166294 374154 166350
rect 374210 166294 374278 166350
rect 374334 166294 374402 166350
rect 374458 166294 374526 166350
rect 374582 166294 404874 166350
rect 404930 166294 404998 166350
rect 405054 166294 405122 166350
rect 405178 166294 405246 166350
rect 405302 166294 435594 166350
rect 435650 166294 435718 166350
rect 435774 166294 435842 166350
rect 435898 166294 435966 166350
rect 436022 166294 466314 166350
rect 466370 166294 466438 166350
rect 466494 166294 466562 166350
rect 466618 166294 466686 166350
rect 466742 166294 497034 166350
rect 497090 166294 497158 166350
rect 497214 166294 497282 166350
rect 497338 166294 497406 166350
rect 497462 166294 527754 166350
rect 527810 166294 527878 166350
rect 527934 166294 528002 166350
rect 528058 166294 528126 166350
rect 528182 166294 558474 166350
rect 558530 166294 558598 166350
rect 558654 166294 558722 166350
rect 558778 166294 558846 166350
rect 558902 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597980 166350
rect -1916 166226 597980 166294
rect -1916 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 36234 166226
rect 36290 166170 36358 166226
rect 36414 166170 36482 166226
rect 36538 166170 36606 166226
rect 36662 166170 44518 166226
rect 44574 166170 44642 166226
rect 44698 166170 75238 166226
rect 75294 166170 75362 166226
rect 75418 166170 105958 166226
rect 106014 166170 106082 166226
rect 106138 166170 136678 166226
rect 136734 166170 136802 166226
rect 136858 166170 167398 166226
rect 167454 166170 167522 166226
rect 167578 166170 198118 166226
rect 198174 166170 198242 166226
rect 198298 166170 228838 166226
rect 228894 166170 228962 166226
rect 229018 166170 259558 166226
rect 259614 166170 259682 166226
rect 259738 166170 281994 166226
rect 282050 166170 282118 166226
rect 282174 166170 282242 166226
rect 282298 166170 282366 166226
rect 282422 166170 312714 166226
rect 312770 166170 312838 166226
rect 312894 166170 312962 166226
rect 313018 166170 313086 166226
rect 313142 166170 343434 166226
rect 343490 166170 343558 166226
rect 343614 166170 343682 166226
rect 343738 166170 343806 166226
rect 343862 166170 374154 166226
rect 374210 166170 374278 166226
rect 374334 166170 374402 166226
rect 374458 166170 374526 166226
rect 374582 166170 404874 166226
rect 404930 166170 404998 166226
rect 405054 166170 405122 166226
rect 405178 166170 405246 166226
rect 405302 166170 435594 166226
rect 435650 166170 435718 166226
rect 435774 166170 435842 166226
rect 435898 166170 435966 166226
rect 436022 166170 466314 166226
rect 466370 166170 466438 166226
rect 466494 166170 466562 166226
rect 466618 166170 466686 166226
rect 466742 166170 497034 166226
rect 497090 166170 497158 166226
rect 497214 166170 497282 166226
rect 497338 166170 497406 166226
rect 497462 166170 527754 166226
rect 527810 166170 527878 166226
rect 527934 166170 528002 166226
rect 528058 166170 528126 166226
rect 528182 166170 558474 166226
rect 558530 166170 558598 166226
rect 558654 166170 558722 166226
rect 558778 166170 558846 166226
rect 558902 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597980 166226
rect -1916 166102 597980 166170
rect -1916 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 36234 166102
rect 36290 166046 36358 166102
rect 36414 166046 36482 166102
rect 36538 166046 36606 166102
rect 36662 166046 44518 166102
rect 44574 166046 44642 166102
rect 44698 166046 75238 166102
rect 75294 166046 75362 166102
rect 75418 166046 105958 166102
rect 106014 166046 106082 166102
rect 106138 166046 136678 166102
rect 136734 166046 136802 166102
rect 136858 166046 167398 166102
rect 167454 166046 167522 166102
rect 167578 166046 198118 166102
rect 198174 166046 198242 166102
rect 198298 166046 228838 166102
rect 228894 166046 228962 166102
rect 229018 166046 259558 166102
rect 259614 166046 259682 166102
rect 259738 166046 281994 166102
rect 282050 166046 282118 166102
rect 282174 166046 282242 166102
rect 282298 166046 282366 166102
rect 282422 166046 312714 166102
rect 312770 166046 312838 166102
rect 312894 166046 312962 166102
rect 313018 166046 313086 166102
rect 313142 166046 343434 166102
rect 343490 166046 343558 166102
rect 343614 166046 343682 166102
rect 343738 166046 343806 166102
rect 343862 166046 374154 166102
rect 374210 166046 374278 166102
rect 374334 166046 374402 166102
rect 374458 166046 374526 166102
rect 374582 166046 404874 166102
rect 404930 166046 404998 166102
rect 405054 166046 405122 166102
rect 405178 166046 405246 166102
rect 405302 166046 435594 166102
rect 435650 166046 435718 166102
rect 435774 166046 435842 166102
rect 435898 166046 435966 166102
rect 436022 166046 466314 166102
rect 466370 166046 466438 166102
rect 466494 166046 466562 166102
rect 466618 166046 466686 166102
rect 466742 166046 497034 166102
rect 497090 166046 497158 166102
rect 497214 166046 497282 166102
rect 497338 166046 497406 166102
rect 497462 166046 527754 166102
rect 527810 166046 527878 166102
rect 527934 166046 528002 166102
rect 528058 166046 528126 166102
rect 528182 166046 558474 166102
rect 558530 166046 558598 166102
rect 558654 166046 558722 166102
rect 558778 166046 558846 166102
rect 558902 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597980 166102
rect -1916 165978 597980 166046
rect -1916 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 36234 165978
rect 36290 165922 36358 165978
rect 36414 165922 36482 165978
rect 36538 165922 36606 165978
rect 36662 165922 44518 165978
rect 44574 165922 44642 165978
rect 44698 165922 75238 165978
rect 75294 165922 75362 165978
rect 75418 165922 105958 165978
rect 106014 165922 106082 165978
rect 106138 165922 136678 165978
rect 136734 165922 136802 165978
rect 136858 165922 167398 165978
rect 167454 165922 167522 165978
rect 167578 165922 198118 165978
rect 198174 165922 198242 165978
rect 198298 165922 228838 165978
rect 228894 165922 228962 165978
rect 229018 165922 259558 165978
rect 259614 165922 259682 165978
rect 259738 165922 281994 165978
rect 282050 165922 282118 165978
rect 282174 165922 282242 165978
rect 282298 165922 282366 165978
rect 282422 165922 312714 165978
rect 312770 165922 312838 165978
rect 312894 165922 312962 165978
rect 313018 165922 313086 165978
rect 313142 165922 343434 165978
rect 343490 165922 343558 165978
rect 343614 165922 343682 165978
rect 343738 165922 343806 165978
rect 343862 165922 374154 165978
rect 374210 165922 374278 165978
rect 374334 165922 374402 165978
rect 374458 165922 374526 165978
rect 374582 165922 404874 165978
rect 404930 165922 404998 165978
rect 405054 165922 405122 165978
rect 405178 165922 405246 165978
rect 405302 165922 435594 165978
rect 435650 165922 435718 165978
rect 435774 165922 435842 165978
rect 435898 165922 435966 165978
rect 436022 165922 466314 165978
rect 466370 165922 466438 165978
rect 466494 165922 466562 165978
rect 466618 165922 466686 165978
rect 466742 165922 497034 165978
rect 497090 165922 497158 165978
rect 497214 165922 497282 165978
rect 497338 165922 497406 165978
rect 497462 165922 527754 165978
rect 527810 165922 527878 165978
rect 527934 165922 528002 165978
rect 528058 165922 528126 165978
rect 528182 165922 558474 165978
rect 558530 165922 558598 165978
rect 558654 165922 558722 165978
rect 558778 165922 558846 165978
rect 558902 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597980 165978
rect -1916 165826 597980 165922
rect 4156 164638 49604 164654
rect 4156 164582 4172 164638
rect 4228 164582 49532 164638
rect 49588 164582 49604 164638
rect 4156 164566 49604 164582
rect -1916 154350 597980 154446
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 9234 154350
rect 9290 154294 9358 154350
rect 9414 154294 9482 154350
rect 9538 154294 9606 154350
rect 9662 154294 39954 154350
rect 40010 154294 40078 154350
rect 40134 154294 40202 154350
rect 40258 154294 40326 154350
rect 40382 154294 59878 154350
rect 59934 154294 60002 154350
rect 60058 154294 90598 154350
rect 90654 154294 90722 154350
rect 90778 154294 121318 154350
rect 121374 154294 121442 154350
rect 121498 154294 152038 154350
rect 152094 154294 152162 154350
rect 152218 154294 182758 154350
rect 182814 154294 182882 154350
rect 182938 154294 213478 154350
rect 213534 154294 213602 154350
rect 213658 154294 244198 154350
rect 244254 154294 244322 154350
rect 244378 154294 285714 154350
rect 285770 154294 285838 154350
rect 285894 154294 285962 154350
rect 286018 154294 286086 154350
rect 286142 154294 316434 154350
rect 316490 154294 316558 154350
rect 316614 154294 316682 154350
rect 316738 154294 316806 154350
rect 316862 154294 347154 154350
rect 347210 154294 347278 154350
rect 347334 154294 347402 154350
rect 347458 154294 347526 154350
rect 347582 154294 377874 154350
rect 377930 154294 377998 154350
rect 378054 154294 378122 154350
rect 378178 154294 378246 154350
rect 378302 154294 408594 154350
rect 408650 154294 408718 154350
rect 408774 154294 408842 154350
rect 408898 154294 408966 154350
rect 409022 154294 439314 154350
rect 439370 154294 439438 154350
rect 439494 154294 439562 154350
rect 439618 154294 439686 154350
rect 439742 154294 470034 154350
rect 470090 154294 470158 154350
rect 470214 154294 470282 154350
rect 470338 154294 470406 154350
rect 470462 154294 500754 154350
rect 500810 154294 500878 154350
rect 500934 154294 501002 154350
rect 501058 154294 501126 154350
rect 501182 154294 531474 154350
rect 531530 154294 531598 154350
rect 531654 154294 531722 154350
rect 531778 154294 531846 154350
rect 531902 154294 562194 154350
rect 562250 154294 562318 154350
rect 562374 154294 562442 154350
rect 562498 154294 562566 154350
rect 562622 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect -1916 154226 597980 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 9234 154226
rect 9290 154170 9358 154226
rect 9414 154170 9482 154226
rect 9538 154170 9606 154226
rect 9662 154170 39954 154226
rect 40010 154170 40078 154226
rect 40134 154170 40202 154226
rect 40258 154170 40326 154226
rect 40382 154170 59878 154226
rect 59934 154170 60002 154226
rect 60058 154170 90598 154226
rect 90654 154170 90722 154226
rect 90778 154170 121318 154226
rect 121374 154170 121442 154226
rect 121498 154170 152038 154226
rect 152094 154170 152162 154226
rect 152218 154170 182758 154226
rect 182814 154170 182882 154226
rect 182938 154170 213478 154226
rect 213534 154170 213602 154226
rect 213658 154170 244198 154226
rect 244254 154170 244322 154226
rect 244378 154170 285714 154226
rect 285770 154170 285838 154226
rect 285894 154170 285962 154226
rect 286018 154170 286086 154226
rect 286142 154170 316434 154226
rect 316490 154170 316558 154226
rect 316614 154170 316682 154226
rect 316738 154170 316806 154226
rect 316862 154170 347154 154226
rect 347210 154170 347278 154226
rect 347334 154170 347402 154226
rect 347458 154170 347526 154226
rect 347582 154170 377874 154226
rect 377930 154170 377998 154226
rect 378054 154170 378122 154226
rect 378178 154170 378246 154226
rect 378302 154170 408594 154226
rect 408650 154170 408718 154226
rect 408774 154170 408842 154226
rect 408898 154170 408966 154226
rect 409022 154170 439314 154226
rect 439370 154170 439438 154226
rect 439494 154170 439562 154226
rect 439618 154170 439686 154226
rect 439742 154170 470034 154226
rect 470090 154170 470158 154226
rect 470214 154170 470282 154226
rect 470338 154170 470406 154226
rect 470462 154170 500754 154226
rect 500810 154170 500878 154226
rect 500934 154170 501002 154226
rect 501058 154170 501126 154226
rect 501182 154170 531474 154226
rect 531530 154170 531598 154226
rect 531654 154170 531722 154226
rect 531778 154170 531846 154226
rect 531902 154170 562194 154226
rect 562250 154170 562318 154226
rect 562374 154170 562442 154226
rect 562498 154170 562566 154226
rect 562622 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect -1916 154102 597980 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 9234 154102
rect 9290 154046 9358 154102
rect 9414 154046 9482 154102
rect 9538 154046 9606 154102
rect 9662 154046 39954 154102
rect 40010 154046 40078 154102
rect 40134 154046 40202 154102
rect 40258 154046 40326 154102
rect 40382 154046 59878 154102
rect 59934 154046 60002 154102
rect 60058 154046 90598 154102
rect 90654 154046 90722 154102
rect 90778 154046 121318 154102
rect 121374 154046 121442 154102
rect 121498 154046 152038 154102
rect 152094 154046 152162 154102
rect 152218 154046 182758 154102
rect 182814 154046 182882 154102
rect 182938 154046 213478 154102
rect 213534 154046 213602 154102
rect 213658 154046 244198 154102
rect 244254 154046 244322 154102
rect 244378 154046 285714 154102
rect 285770 154046 285838 154102
rect 285894 154046 285962 154102
rect 286018 154046 286086 154102
rect 286142 154046 316434 154102
rect 316490 154046 316558 154102
rect 316614 154046 316682 154102
rect 316738 154046 316806 154102
rect 316862 154046 347154 154102
rect 347210 154046 347278 154102
rect 347334 154046 347402 154102
rect 347458 154046 347526 154102
rect 347582 154046 377874 154102
rect 377930 154046 377998 154102
rect 378054 154046 378122 154102
rect 378178 154046 378246 154102
rect 378302 154046 408594 154102
rect 408650 154046 408718 154102
rect 408774 154046 408842 154102
rect 408898 154046 408966 154102
rect 409022 154046 439314 154102
rect 439370 154046 439438 154102
rect 439494 154046 439562 154102
rect 439618 154046 439686 154102
rect 439742 154046 470034 154102
rect 470090 154046 470158 154102
rect 470214 154046 470282 154102
rect 470338 154046 470406 154102
rect 470462 154046 500754 154102
rect 500810 154046 500878 154102
rect 500934 154046 501002 154102
rect 501058 154046 501126 154102
rect 501182 154046 531474 154102
rect 531530 154046 531598 154102
rect 531654 154046 531722 154102
rect 531778 154046 531846 154102
rect 531902 154046 562194 154102
rect 562250 154046 562318 154102
rect 562374 154046 562442 154102
rect 562498 154046 562566 154102
rect 562622 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect -1916 153978 597980 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 9234 153978
rect 9290 153922 9358 153978
rect 9414 153922 9482 153978
rect 9538 153922 9606 153978
rect 9662 153922 39954 153978
rect 40010 153922 40078 153978
rect 40134 153922 40202 153978
rect 40258 153922 40326 153978
rect 40382 153922 59878 153978
rect 59934 153922 60002 153978
rect 60058 153922 90598 153978
rect 90654 153922 90722 153978
rect 90778 153922 121318 153978
rect 121374 153922 121442 153978
rect 121498 153922 152038 153978
rect 152094 153922 152162 153978
rect 152218 153922 182758 153978
rect 182814 153922 182882 153978
rect 182938 153922 213478 153978
rect 213534 153922 213602 153978
rect 213658 153922 244198 153978
rect 244254 153922 244322 153978
rect 244378 153922 285714 153978
rect 285770 153922 285838 153978
rect 285894 153922 285962 153978
rect 286018 153922 286086 153978
rect 286142 153922 316434 153978
rect 316490 153922 316558 153978
rect 316614 153922 316682 153978
rect 316738 153922 316806 153978
rect 316862 153922 347154 153978
rect 347210 153922 347278 153978
rect 347334 153922 347402 153978
rect 347458 153922 347526 153978
rect 347582 153922 377874 153978
rect 377930 153922 377998 153978
rect 378054 153922 378122 153978
rect 378178 153922 378246 153978
rect 378302 153922 408594 153978
rect 408650 153922 408718 153978
rect 408774 153922 408842 153978
rect 408898 153922 408966 153978
rect 409022 153922 439314 153978
rect 439370 153922 439438 153978
rect 439494 153922 439562 153978
rect 439618 153922 439686 153978
rect 439742 153922 470034 153978
rect 470090 153922 470158 153978
rect 470214 153922 470282 153978
rect 470338 153922 470406 153978
rect 470462 153922 500754 153978
rect 500810 153922 500878 153978
rect 500934 153922 501002 153978
rect 501058 153922 501126 153978
rect 501182 153922 531474 153978
rect 531530 153922 531598 153978
rect 531654 153922 531722 153978
rect 531778 153922 531846 153978
rect 531902 153922 562194 153978
rect 562250 153922 562318 153978
rect 562374 153922 562442 153978
rect 562498 153922 562566 153978
rect 562622 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect -1916 153826 597980 153922
rect 313388 153658 495924 153674
rect 313388 153602 313404 153658
rect 313460 153602 372428 153658
rect 372484 153602 495852 153658
rect 495908 153602 495924 153658
rect 313388 153586 495924 153602
rect 273740 152938 501412 152954
rect 273740 152882 273756 152938
rect 273812 152882 501340 152938
rect 501396 152882 501412 152938
rect 273740 152866 501412 152882
rect -1916 148350 597980 148446
rect -1916 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 36234 148350
rect 36290 148294 36358 148350
rect 36414 148294 36482 148350
rect 36538 148294 36606 148350
rect 36662 148294 44518 148350
rect 44574 148294 44642 148350
rect 44698 148294 75238 148350
rect 75294 148294 75362 148350
rect 75418 148294 105958 148350
rect 106014 148294 106082 148350
rect 106138 148294 136678 148350
rect 136734 148294 136802 148350
rect 136858 148294 167398 148350
rect 167454 148294 167522 148350
rect 167578 148294 198118 148350
rect 198174 148294 198242 148350
rect 198298 148294 228838 148350
rect 228894 148294 228962 148350
rect 229018 148294 259558 148350
rect 259614 148294 259682 148350
rect 259738 148294 281994 148350
rect 282050 148294 282118 148350
rect 282174 148294 282242 148350
rect 282298 148294 282366 148350
rect 282422 148294 312714 148350
rect 312770 148294 312838 148350
rect 312894 148294 312962 148350
rect 313018 148294 313086 148350
rect 313142 148294 343434 148350
rect 343490 148294 343558 148350
rect 343614 148294 343682 148350
rect 343738 148294 343806 148350
rect 343862 148294 374154 148350
rect 374210 148294 374278 148350
rect 374334 148294 374402 148350
rect 374458 148294 374526 148350
rect 374582 148294 404874 148350
rect 404930 148294 404998 148350
rect 405054 148294 405122 148350
rect 405178 148294 405246 148350
rect 405302 148294 435594 148350
rect 435650 148294 435718 148350
rect 435774 148294 435842 148350
rect 435898 148294 435966 148350
rect 436022 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597980 148350
rect -1916 148226 597980 148294
rect -1916 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 36234 148226
rect 36290 148170 36358 148226
rect 36414 148170 36482 148226
rect 36538 148170 36606 148226
rect 36662 148170 44518 148226
rect 44574 148170 44642 148226
rect 44698 148170 75238 148226
rect 75294 148170 75362 148226
rect 75418 148170 105958 148226
rect 106014 148170 106082 148226
rect 106138 148170 136678 148226
rect 136734 148170 136802 148226
rect 136858 148170 167398 148226
rect 167454 148170 167522 148226
rect 167578 148170 198118 148226
rect 198174 148170 198242 148226
rect 198298 148170 228838 148226
rect 228894 148170 228962 148226
rect 229018 148170 259558 148226
rect 259614 148170 259682 148226
rect 259738 148170 281994 148226
rect 282050 148170 282118 148226
rect 282174 148170 282242 148226
rect 282298 148170 282366 148226
rect 282422 148170 312714 148226
rect 312770 148170 312838 148226
rect 312894 148170 312962 148226
rect 313018 148170 313086 148226
rect 313142 148170 343434 148226
rect 343490 148170 343558 148226
rect 343614 148170 343682 148226
rect 343738 148170 343806 148226
rect 343862 148170 374154 148226
rect 374210 148170 374278 148226
rect 374334 148170 374402 148226
rect 374458 148170 374526 148226
rect 374582 148170 404874 148226
rect 404930 148170 404998 148226
rect 405054 148170 405122 148226
rect 405178 148170 405246 148226
rect 405302 148170 435594 148226
rect 435650 148170 435718 148226
rect 435774 148170 435842 148226
rect 435898 148170 435966 148226
rect 436022 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597980 148226
rect -1916 148102 597980 148170
rect -1916 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 36234 148102
rect 36290 148046 36358 148102
rect 36414 148046 36482 148102
rect 36538 148046 36606 148102
rect 36662 148046 44518 148102
rect 44574 148046 44642 148102
rect 44698 148046 75238 148102
rect 75294 148046 75362 148102
rect 75418 148046 105958 148102
rect 106014 148046 106082 148102
rect 106138 148046 136678 148102
rect 136734 148046 136802 148102
rect 136858 148046 167398 148102
rect 167454 148046 167522 148102
rect 167578 148046 198118 148102
rect 198174 148046 198242 148102
rect 198298 148046 228838 148102
rect 228894 148046 228962 148102
rect 229018 148046 259558 148102
rect 259614 148046 259682 148102
rect 259738 148046 281994 148102
rect 282050 148046 282118 148102
rect 282174 148046 282242 148102
rect 282298 148046 282366 148102
rect 282422 148046 312714 148102
rect 312770 148046 312838 148102
rect 312894 148046 312962 148102
rect 313018 148046 313086 148102
rect 313142 148046 343434 148102
rect 343490 148046 343558 148102
rect 343614 148046 343682 148102
rect 343738 148046 343806 148102
rect 343862 148046 374154 148102
rect 374210 148046 374278 148102
rect 374334 148046 374402 148102
rect 374458 148046 374526 148102
rect 374582 148046 404874 148102
rect 404930 148046 404998 148102
rect 405054 148046 405122 148102
rect 405178 148046 405246 148102
rect 405302 148046 435594 148102
rect 435650 148046 435718 148102
rect 435774 148046 435842 148102
rect 435898 148046 435966 148102
rect 436022 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597980 148102
rect -1916 147978 597980 148046
rect -1916 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 36234 147978
rect 36290 147922 36358 147978
rect 36414 147922 36482 147978
rect 36538 147922 36606 147978
rect 36662 147922 44518 147978
rect 44574 147922 44642 147978
rect 44698 147922 75238 147978
rect 75294 147922 75362 147978
rect 75418 147922 105958 147978
rect 106014 147922 106082 147978
rect 106138 147922 136678 147978
rect 136734 147922 136802 147978
rect 136858 147922 167398 147978
rect 167454 147922 167522 147978
rect 167578 147922 198118 147978
rect 198174 147922 198242 147978
rect 198298 147922 228838 147978
rect 228894 147922 228962 147978
rect 229018 147922 259558 147978
rect 259614 147922 259682 147978
rect 259738 147922 281994 147978
rect 282050 147922 282118 147978
rect 282174 147922 282242 147978
rect 282298 147922 282366 147978
rect 282422 147922 312714 147978
rect 312770 147922 312838 147978
rect 312894 147922 312962 147978
rect 313018 147922 313086 147978
rect 313142 147922 343434 147978
rect 343490 147922 343558 147978
rect 343614 147922 343682 147978
rect 343738 147922 343806 147978
rect 343862 147922 374154 147978
rect 374210 147922 374278 147978
rect 374334 147922 374402 147978
rect 374458 147922 374526 147978
rect 374582 147922 404874 147978
rect 404930 147922 404998 147978
rect 405054 147922 405122 147978
rect 405178 147922 405246 147978
rect 405302 147922 435594 147978
rect 435650 147922 435718 147978
rect 435774 147922 435842 147978
rect 435898 147922 435966 147978
rect 436022 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597980 147978
rect -1916 147826 597980 147922
rect -1916 136350 597980 136446
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 9234 136350
rect 9290 136294 9358 136350
rect 9414 136294 9482 136350
rect 9538 136294 9606 136350
rect 9662 136294 39954 136350
rect 40010 136294 40078 136350
rect 40134 136294 40202 136350
rect 40258 136294 40326 136350
rect 40382 136294 59878 136350
rect 59934 136294 60002 136350
rect 60058 136294 90598 136350
rect 90654 136294 90722 136350
rect 90778 136294 121318 136350
rect 121374 136294 121442 136350
rect 121498 136294 152038 136350
rect 152094 136294 152162 136350
rect 152218 136294 182758 136350
rect 182814 136294 182882 136350
rect 182938 136294 213478 136350
rect 213534 136294 213602 136350
rect 213658 136294 244198 136350
rect 244254 136294 244322 136350
rect 244378 136294 285714 136350
rect 285770 136294 285838 136350
rect 285894 136294 285962 136350
rect 286018 136294 286086 136350
rect 286142 136294 316434 136350
rect 316490 136294 316558 136350
rect 316614 136294 316682 136350
rect 316738 136294 316806 136350
rect 316862 136294 347154 136350
rect 347210 136294 347278 136350
rect 347334 136294 347402 136350
rect 347458 136294 347526 136350
rect 347582 136294 377874 136350
rect 377930 136294 377998 136350
rect 378054 136294 378122 136350
rect 378178 136294 378246 136350
rect 378302 136294 408594 136350
rect 408650 136294 408718 136350
rect 408774 136294 408842 136350
rect 408898 136294 408966 136350
rect 409022 136294 439314 136350
rect 439370 136294 439438 136350
rect 439494 136294 439562 136350
rect 439618 136294 439686 136350
rect 439742 136294 479878 136350
rect 479934 136294 480002 136350
rect 480058 136294 510598 136350
rect 510654 136294 510722 136350
rect 510778 136294 541318 136350
rect 541374 136294 541442 136350
rect 541498 136294 562194 136350
rect 562250 136294 562318 136350
rect 562374 136294 562442 136350
rect 562498 136294 562566 136350
rect 562622 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect -1916 136226 597980 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 9234 136226
rect 9290 136170 9358 136226
rect 9414 136170 9482 136226
rect 9538 136170 9606 136226
rect 9662 136170 39954 136226
rect 40010 136170 40078 136226
rect 40134 136170 40202 136226
rect 40258 136170 40326 136226
rect 40382 136170 59878 136226
rect 59934 136170 60002 136226
rect 60058 136170 90598 136226
rect 90654 136170 90722 136226
rect 90778 136170 121318 136226
rect 121374 136170 121442 136226
rect 121498 136170 152038 136226
rect 152094 136170 152162 136226
rect 152218 136170 182758 136226
rect 182814 136170 182882 136226
rect 182938 136170 213478 136226
rect 213534 136170 213602 136226
rect 213658 136170 244198 136226
rect 244254 136170 244322 136226
rect 244378 136170 285714 136226
rect 285770 136170 285838 136226
rect 285894 136170 285962 136226
rect 286018 136170 286086 136226
rect 286142 136170 316434 136226
rect 316490 136170 316558 136226
rect 316614 136170 316682 136226
rect 316738 136170 316806 136226
rect 316862 136170 347154 136226
rect 347210 136170 347278 136226
rect 347334 136170 347402 136226
rect 347458 136170 347526 136226
rect 347582 136170 377874 136226
rect 377930 136170 377998 136226
rect 378054 136170 378122 136226
rect 378178 136170 378246 136226
rect 378302 136170 408594 136226
rect 408650 136170 408718 136226
rect 408774 136170 408842 136226
rect 408898 136170 408966 136226
rect 409022 136170 439314 136226
rect 439370 136170 439438 136226
rect 439494 136170 439562 136226
rect 439618 136170 439686 136226
rect 439742 136170 479878 136226
rect 479934 136170 480002 136226
rect 480058 136170 510598 136226
rect 510654 136170 510722 136226
rect 510778 136170 541318 136226
rect 541374 136170 541442 136226
rect 541498 136170 562194 136226
rect 562250 136170 562318 136226
rect 562374 136170 562442 136226
rect 562498 136170 562566 136226
rect 562622 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect -1916 136102 597980 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 9234 136102
rect 9290 136046 9358 136102
rect 9414 136046 9482 136102
rect 9538 136046 9606 136102
rect 9662 136046 39954 136102
rect 40010 136046 40078 136102
rect 40134 136046 40202 136102
rect 40258 136046 40326 136102
rect 40382 136046 59878 136102
rect 59934 136046 60002 136102
rect 60058 136046 90598 136102
rect 90654 136046 90722 136102
rect 90778 136046 121318 136102
rect 121374 136046 121442 136102
rect 121498 136046 152038 136102
rect 152094 136046 152162 136102
rect 152218 136046 182758 136102
rect 182814 136046 182882 136102
rect 182938 136046 213478 136102
rect 213534 136046 213602 136102
rect 213658 136046 244198 136102
rect 244254 136046 244322 136102
rect 244378 136046 285714 136102
rect 285770 136046 285838 136102
rect 285894 136046 285962 136102
rect 286018 136046 286086 136102
rect 286142 136046 316434 136102
rect 316490 136046 316558 136102
rect 316614 136046 316682 136102
rect 316738 136046 316806 136102
rect 316862 136046 347154 136102
rect 347210 136046 347278 136102
rect 347334 136046 347402 136102
rect 347458 136046 347526 136102
rect 347582 136046 377874 136102
rect 377930 136046 377998 136102
rect 378054 136046 378122 136102
rect 378178 136046 378246 136102
rect 378302 136046 408594 136102
rect 408650 136046 408718 136102
rect 408774 136046 408842 136102
rect 408898 136046 408966 136102
rect 409022 136046 439314 136102
rect 439370 136046 439438 136102
rect 439494 136046 439562 136102
rect 439618 136046 439686 136102
rect 439742 136046 479878 136102
rect 479934 136046 480002 136102
rect 480058 136046 510598 136102
rect 510654 136046 510722 136102
rect 510778 136046 541318 136102
rect 541374 136046 541442 136102
rect 541498 136046 562194 136102
rect 562250 136046 562318 136102
rect 562374 136046 562442 136102
rect 562498 136046 562566 136102
rect 562622 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect -1916 135978 597980 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 9234 135978
rect 9290 135922 9358 135978
rect 9414 135922 9482 135978
rect 9538 135922 9606 135978
rect 9662 135922 39954 135978
rect 40010 135922 40078 135978
rect 40134 135922 40202 135978
rect 40258 135922 40326 135978
rect 40382 135922 59878 135978
rect 59934 135922 60002 135978
rect 60058 135922 90598 135978
rect 90654 135922 90722 135978
rect 90778 135922 121318 135978
rect 121374 135922 121442 135978
rect 121498 135922 152038 135978
rect 152094 135922 152162 135978
rect 152218 135922 182758 135978
rect 182814 135922 182882 135978
rect 182938 135922 213478 135978
rect 213534 135922 213602 135978
rect 213658 135922 244198 135978
rect 244254 135922 244322 135978
rect 244378 135922 285714 135978
rect 285770 135922 285838 135978
rect 285894 135922 285962 135978
rect 286018 135922 286086 135978
rect 286142 135922 316434 135978
rect 316490 135922 316558 135978
rect 316614 135922 316682 135978
rect 316738 135922 316806 135978
rect 316862 135922 347154 135978
rect 347210 135922 347278 135978
rect 347334 135922 347402 135978
rect 347458 135922 347526 135978
rect 347582 135922 377874 135978
rect 377930 135922 377998 135978
rect 378054 135922 378122 135978
rect 378178 135922 378246 135978
rect 378302 135922 408594 135978
rect 408650 135922 408718 135978
rect 408774 135922 408842 135978
rect 408898 135922 408966 135978
rect 409022 135922 439314 135978
rect 439370 135922 439438 135978
rect 439494 135922 439562 135978
rect 439618 135922 439686 135978
rect 439742 135922 479878 135978
rect 479934 135922 480002 135978
rect 480058 135922 510598 135978
rect 510654 135922 510722 135978
rect 510778 135922 541318 135978
rect 541374 135922 541442 135978
rect 541498 135922 562194 135978
rect 562250 135922 562318 135978
rect 562374 135922 562442 135978
rect 562498 135922 562566 135978
rect 562622 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect -1916 135826 597980 135922
rect -1916 130350 597980 130446
rect -1916 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 36234 130350
rect 36290 130294 36358 130350
rect 36414 130294 36482 130350
rect 36538 130294 36606 130350
rect 36662 130294 44518 130350
rect 44574 130294 44642 130350
rect 44698 130294 75238 130350
rect 75294 130294 75362 130350
rect 75418 130294 105958 130350
rect 106014 130294 106082 130350
rect 106138 130294 136678 130350
rect 136734 130294 136802 130350
rect 136858 130294 167398 130350
rect 167454 130294 167522 130350
rect 167578 130294 198118 130350
rect 198174 130294 198242 130350
rect 198298 130294 228838 130350
rect 228894 130294 228962 130350
rect 229018 130294 259558 130350
rect 259614 130294 259682 130350
rect 259738 130294 281994 130350
rect 282050 130294 282118 130350
rect 282174 130294 282242 130350
rect 282298 130294 282366 130350
rect 282422 130294 312714 130350
rect 312770 130294 312838 130350
rect 312894 130294 312962 130350
rect 313018 130294 313086 130350
rect 313142 130294 343434 130350
rect 343490 130294 343558 130350
rect 343614 130294 343682 130350
rect 343738 130294 343806 130350
rect 343862 130294 374154 130350
rect 374210 130294 374278 130350
rect 374334 130294 374402 130350
rect 374458 130294 374526 130350
rect 374582 130294 404874 130350
rect 404930 130294 404998 130350
rect 405054 130294 405122 130350
rect 405178 130294 405246 130350
rect 405302 130294 435594 130350
rect 435650 130294 435718 130350
rect 435774 130294 435842 130350
rect 435898 130294 435966 130350
rect 436022 130294 464518 130350
rect 464574 130294 464642 130350
rect 464698 130294 495238 130350
rect 495294 130294 495362 130350
rect 495418 130294 525958 130350
rect 526014 130294 526082 130350
rect 526138 130294 556678 130350
rect 556734 130294 556802 130350
rect 556858 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597980 130350
rect -1916 130226 597980 130294
rect -1916 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 36234 130226
rect 36290 130170 36358 130226
rect 36414 130170 36482 130226
rect 36538 130170 36606 130226
rect 36662 130170 44518 130226
rect 44574 130170 44642 130226
rect 44698 130170 75238 130226
rect 75294 130170 75362 130226
rect 75418 130170 105958 130226
rect 106014 130170 106082 130226
rect 106138 130170 136678 130226
rect 136734 130170 136802 130226
rect 136858 130170 167398 130226
rect 167454 130170 167522 130226
rect 167578 130170 198118 130226
rect 198174 130170 198242 130226
rect 198298 130170 228838 130226
rect 228894 130170 228962 130226
rect 229018 130170 259558 130226
rect 259614 130170 259682 130226
rect 259738 130170 281994 130226
rect 282050 130170 282118 130226
rect 282174 130170 282242 130226
rect 282298 130170 282366 130226
rect 282422 130170 312714 130226
rect 312770 130170 312838 130226
rect 312894 130170 312962 130226
rect 313018 130170 313086 130226
rect 313142 130170 343434 130226
rect 343490 130170 343558 130226
rect 343614 130170 343682 130226
rect 343738 130170 343806 130226
rect 343862 130170 374154 130226
rect 374210 130170 374278 130226
rect 374334 130170 374402 130226
rect 374458 130170 374526 130226
rect 374582 130170 404874 130226
rect 404930 130170 404998 130226
rect 405054 130170 405122 130226
rect 405178 130170 405246 130226
rect 405302 130170 435594 130226
rect 435650 130170 435718 130226
rect 435774 130170 435842 130226
rect 435898 130170 435966 130226
rect 436022 130170 464518 130226
rect 464574 130170 464642 130226
rect 464698 130170 495238 130226
rect 495294 130170 495362 130226
rect 495418 130170 525958 130226
rect 526014 130170 526082 130226
rect 526138 130170 556678 130226
rect 556734 130170 556802 130226
rect 556858 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597980 130226
rect -1916 130102 597980 130170
rect -1916 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 36234 130102
rect 36290 130046 36358 130102
rect 36414 130046 36482 130102
rect 36538 130046 36606 130102
rect 36662 130046 44518 130102
rect 44574 130046 44642 130102
rect 44698 130046 75238 130102
rect 75294 130046 75362 130102
rect 75418 130046 105958 130102
rect 106014 130046 106082 130102
rect 106138 130046 136678 130102
rect 136734 130046 136802 130102
rect 136858 130046 167398 130102
rect 167454 130046 167522 130102
rect 167578 130046 198118 130102
rect 198174 130046 198242 130102
rect 198298 130046 228838 130102
rect 228894 130046 228962 130102
rect 229018 130046 259558 130102
rect 259614 130046 259682 130102
rect 259738 130046 281994 130102
rect 282050 130046 282118 130102
rect 282174 130046 282242 130102
rect 282298 130046 282366 130102
rect 282422 130046 312714 130102
rect 312770 130046 312838 130102
rect 312894 130046 312962 130102
rect 313018 130046 313086 130102
rect 313142 130046 343434 130102
rect 343490 130046 343558 130102
rect 343614 130046 343682 130102
rect 343738 130046 343806 130102
rect 343862 130046 374154 130102
rect 374210 130046 374278 130102
rect 374334 130046 374402 130102
rect 374458 130046 374526 130102
rect 374582 130046 404874 130102
rect 404930 130046 404998 130102
rect 405054 130046 405122 130102
rect 405178 130046 405246 130102
rect 405302 130046 435594 130102
rect 435650 130046 435718 130102
rect 435774 130046 435842 130102
rect 435898 130046 435966 130102
rect 436022 130046 464518 130102
rect 464574 130046 464642 130102
rect 464698 130046 495238 130102
rect 495294 130046 495362 130102
rect 495418 130046 525958 130102
rect 526014 130046 526082 130102
rect 526138 130046 556678 130102
rect 556734 130046 556802 130102
rect 556858 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597980 130102
rect -1916 129978 597980 130046
rect -1916 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 36234 129978
rect 36290 129922 36358 129978
rect 36414 129922 36482 129978
rect 36538 129922 36606 129978
rect 36662 129922 44518 129978
rect 44574 129922 44642 129978
rect 44698 129922 75238 129978
rect 75294 129922 75362 129978
rect 75418 129922 105958 129978
rect 106014 129922 106082 129978
rect 106138 129922 136678 129978
rect 136734 129922 136802 129978
rect 136858 129922 167398 129978
rect 167454 129922 167522 129978
rect 167578 129922 198118 129978
rect 198174 129922 198242 129978
rect 198298 129922 228838 129978
rect 228894 129922 228962 129978
rect 229018 129922 259558 129978
rect 259614 129922 259682 129978
rect 259738 129922 281994 129978
rect 282050 129922 282118 129978
rect 282174 129922 282242 129978
rect 282298 129922 282366 129978
rect 282422 129922 312714 129978
rect 312770 129922 312838 129978
rect 312894 129922 312962 129978
rect 313018 129922 313086 129978
rect 313142 129922 343434 129978
rect 343490 129922 343558 129978
rect 343614 129922 343682 129978
rect 343738 129922 343806 129978
rect 343862 129922 374154 129978
rect 374210 129922 374278 129978
rect 374334 129922 374402 129978
rect 374458 129922 374526 129978
rect 374582 129922 404874 129978
rect 404930 129922 404998 129978
rect 405054 129922 405122 129978
rect 405178 129922 405246 129978
rect 405302 129922 435594 129978
rect 435650 129922 435718 129978
rect 435774 129922 435842 129978
rect 435898 129922 435966 129978
rect 436022 129922 464518 129978
rect 464574 129922 464642 129978
rect 464698 129922 495238 129978
rect 495294 129922 495362 129978
rect 495418 129922 525958 129978
rect 526014 129922 526082 129978
rect 526138 129922 556678 129978
rect 556734 129922 556802 129978
rect 556858 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597980 129978
rect -1916 129826 597980 129922
rect -1916 118350 597980 118446
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 9234 118350
rect 9290 118294 9358 118350
rect 9414 118294 9482 118350
rect 9538 118294 9606 118350
rect 9662 118294 39954 118350
rect 40010 118294 40078 118350
rect 40134 118294 40202 118350
rect 40258 118294 40326 118350
rect 40382 118294 59878 118350
rect 59934 118294 60002 118350
rect 60058 118294 90598 118350
rect 90654 118294 90722 118350
rect 90778 118294 121318 118350
rect 121374 118294 121442 118350
rect 121498 118294 152038 118350
rect 152094 118294 152162 118350
rect 152218 118294 182758 118350
rect 182814 118294 182882 118350
rect 182938 118294 213478 118350
rect 213534 118294 213602 118350
rect 213658 118294 244198 118350
rect 244254 118294 244322 118350
rect 244378 118294 285714 118350
rect 285770 118294 285838 118350
rect 285894 118294 285962 118350
rect 286018 118294 286086 118350
rect 286142 118294 316434 118350
rect 316490 118294 316558 118350
rect 316614 118294 316682 118350
rect 316738 118294 316806 118350
rect 316862 118294 347154 118350
rect 347210 118294 347278 118350
rect 347334 118294 347402 118350
rect 347458 118294 347526 118350
rect 347582 118294 377874 118350
rect 377930 118294 377998 118350
rect 378054 118294 378122 118350
rect 378178 118294 378246 118350
rect 378302 118294 408594 118350
rect 408650 118294 408718 118350
rect 408774 118294 408842 118350
rect 408898 118294 408966 118350
rect 409022 118294 439314 118350
rect 439370 118294 439438 118350
rect 439494 118294 439562 118350
rect 439618 118294 439686 118350
rect 439742 118294 479878 118350
rect 479934 118294 480002 118350
rect 480058 118294 510598 118350
rect 510654 118294 510722 118350
rect 510778 118294 541318 118350
rect 541374 118294 541442 118350
rect 541498 118294 562194 118350
rect 562250 118294 562318 118350
rect 562374 118294 562442 118350
rect 562498 118294 562566 118350
rect 562622 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect -1916 118226 597980 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 9234 118226
rect 9290 118170 9358 118226
rect 9414 118170 9482 118226
rect 9538 118170 9606 118226
rect 9662 118170 39954 118226
rect 40010 118170 40078 118226
rect 40134 118170 40202 118226
rect 40258 118170 40326 118226
rect 40382 118170 59878 118226
rect 59934 118170 60002 118226
rect 60058 118170 90598 118226
rect 90654 118170 90722 118226
rect 90778 118170 121318 118226
rect 121374 118170 121442 118226
rect 121498 118170 152038 118226
rect 152094 118170 152162 118226
rect 152218 118170 182758 118226
rect 182814 118170 182882 118226
rect 182938 118170 213478 118226
rect 213534 118170 213602 118226
rect 213658 118170 244198 118226
rect 244254 118170 244322 118226
rect 244378 118170 285714 118226
rect 285770 118170 285838 118226
rect 285894 118170 285962 118226
rect 286018 118170 286086 118226
rect 286142 118170 316434 118226
rect 316490 118170 316558 118226
rect 316614 118170 316682 118226
rect 316738 118170 316806 118226
rect 316862 118170 347154 118226
rect 347210 118170 347278 118226
rect 347334 118170 347402 118226
rect 347458 118170 347526 118226
rect 347582 118170 377874 118226
rect 377930 118170 377998 118226
rect 378054 118170 378122 118226
rect 378178 118170 378246 118226
rect 378302 118170 408594 118226
rect 408650 118170 408718 118226
rect 408774 118170 408842 118226
rect 408898 118170 408966 118226
rect 409022 118170 439314 118226
rect 439370 118170 439438 118226
rect 439494 118170 439562 118226
rect 439618 118170 439686 118226
rect 439742 118170 479878 118226
rect 479934 118170 480002 118226
rect 480058 118170 510598 118226
rect 510654 118170 510722 118226
rect 510778 118170 541318 118226
rect 541374 118170 541442 118226
rect 541498 118170 562194 118226
rect 562250 118170 562318 118226
rect 562374 118170 562442 118226
rect 562498 118170 562566 118226
rect 562622 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect -1916 118102 597980 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 9234 118102
rect 9290 118046 9358 118102
rect 9414 118046 9482 118102
rect 9538 118046 9606 118102
rect 9662 118046 39954 118102
rect 40010 118046 40078 118102
rect 40134 118046 40202 118102
rect 40258 118046 40326 118102
rect 40382 118046 59878 118102
rect 59934 118046 60002 118102
rect 60058 118046 90598 118102
rect 90654 118046 90722 118102
rect 90778 118046 121318 118102
rect 121374 118046 121442 118102
rect 121498 118046 152038 118102
rect 152094 118046 152162 118102
rect 152218 118046 182758 118102
rect 182814 118046 182882 118102
rect 182938 118046 213478 118102
rect 213534 118046 213602 118102
rect 213658 118046 244198 118102
rect 244254 118046 244322 118102
rect 244378 118046 285714 118102
rect 285770 118046 285838 118102
rect 285894 118046 285962 118102
rect 286018 118046 286086 118102
rect 286142 118046 316434 118102
rect 316490 118046 316558 118102
rect 316614 118046 316682 118102
rect 316738 118046 316806 118102
rect 316862 118046 347154 118102
rect 347210 118046 347278 118102
rect 347334 118046 347402 118102
rect 347458 118046 347526 118102
rect 347582 118046 377874 118102
rect 377930 118046 377998 118102
rect 378054 118046 378122 118102
rect 378178 118046 378246 118102
rect 378302 118046 408594 118102
rect 408650 118046 408718 118102
rect 408774 118046 408842 118102
rect 408898 118046 408966 118102
rect 409022 118046 439314 118102
rect 439370 118046 439438 118102
rect 439494 118046 439562 118102
rect 439618 118046 439686 118102
rect 439742 118046 479878 118102
rect 479934 118046 480002 118102
rect 480058 118046 510598 118102
rect 510654 118046 510722 118102
rect 510778 118046 541318 118102
rect 541374 118046 541442 118102
rect 541498 118046 562194 118102
rect 562250 118046 562318 118102
rect 562374 118046 562442 118102
rect 562498 118046 562566 118102
rect 562622 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect -1916 117978 597980 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 9234 117978
rect 9290 117922 9358 117978
rect 9414 117922 9482 117978
rect 9538 117922 9606 117978
rect 9662 117922 39954 117978
rect 40010 117922 40078 117978
rect 40134 117922 40202 117978
rect 40258 117922 40326 117978
rect 40382 117922 59878 117978
rect 59934 117922 60002 117978
rect 60058 117922 90598 117978
rect 90654 117922 90722 117978
rect 90778 117922 121318 117978
rect 121374 117922 121442 117978
rect 121498 117922 152038 117978
rect 152094 117922 152162 117978
rect 152218 117922 182758 117978
rect 182814 117922 182882 117978
rect 182938 117922 213478 117978
rect 213534 117922 213602 117978
rect 213658 117922 244198 117978
rect 244254 117922 244322 117978
rect 244378 117922 285714 117978
rect 285770 117922 285838 117978
rect 285894 117922 285962 117978
rect 286018 117922 286086 117978
rect 286142 117922 316434 117978
rect 316490 117922 316558 117978
rect 316614 117922 316682 117978
rect 316738 117922 316806 117978
rect 316862 117922 347154 117978
rect 347210 117922 347278 117978
rect 347334 117922 347402 117978
rect 347458 117922 347526 117978
rect 347582 117922 377874 117978
rect 377930 117922 377998 117978
rect 378054 117922 378122 117978
rect 378178 117922 378246 117978
rect 378302 117922 408594 117978
rect 408650 117922 408718 117978
rect 408774 117922 408842 117978
rect 408898 117922 408966 117978
rect 409022 117922 439314 117978
rect 439370 117922 439438 117978
rect 439494 117922 439562 117978
rect 439618 117922 439686 117978
rect 439742 117922 479878 117978
rect 479934 117922 480002 117978
rect 480058 117922 510598 117978
rect 510654 117922 510722 117978
rect 510778 117922 541318 117978
rect 541374 117922 541442 117978
rect 541498 117922 562194 117978
rect 562250 117922 562318 117978
rect 562374 117922 562442 117978
rect 562498 117922 562566 117978
rect 562622 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect -1916 117826 597980 117922
rect -1916 112350 597980 112446
rect -1916 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 36234 112350
rect 36290 112294 36358 112350
rect 36414 112294 36482 112350
rect 36538 112294 36606 112350
rect 36662 112294 44518 112350
rect 44574 112294 44642 112350
rect 44698 112294 75238 112350
rect 75294 112294 75362 112350
rect 75418 112294 105958 112350
rect 106014 112294 106082 112350
rect 106138 112294 136678 112350
rect 136734 112294 136802 112350
rect 136858 112294 167398 112350
rect 167454 112294 167522 112350
rect 167578 112294 198118 112350
rect 198174 112294 198242 112350
rect 198298 112294 228838 112350
rect 228894 112294 228962 112350
rect 229018 112294 259558 112350
rect 259614 112294 259682 112350
rect 259738 112294 281994 112350
rect 282050 112294 282118 112350
rect 282174 112294 282242 112350
rect 282298 112294 282366 112350
rect 282422 112294 312714 112350
rect 312770 112294 312838 112350
rect 312894 112294 312962 112350
rect 313018 112294 313086 112350
rect 313142 112294 343434 112350
rect 343490 112294 343558 112350
rect 343614 112294 343682 112350
rect 343738 112294 343806 112350
rect 343862 112294 364518 112350
rect 364574 112294 364642 112350
rect 364698 112294 395238 112350
rect 395294 112294 395362 112350
rect 395418 112294 435594 112350
rect 435650 112294 435718 112350
rect 435774 112294 435842 112350
rect 435898 112294 435966 112350
rect 436022 112294 464518 112350
rect 464574 112294 464642 112350
rect 464698 112294 495238 112350
rect 495294 112294 495362 112350
rect 495418 112294 525958 112350
rect 526014 112294 526082 112350
rect 526138 112294 556678 112350
rect 556734 112294 556802 112350
rect 556858 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597980 112350
rect -1916 112226 597980 112294
rect -1916 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 36234 112226
rect 36290 112170 36358 112226
rect 36414 112170 36482 112226
rect 36538 112170 36606 112226
rect 36662 112170 44518 112226
rect 44574 112170 44642 112226
rect 44698 112170 75238 112226
rect 75294 112170 75362 112226
rect 75418 112170 105958 112226
rect 106014 112170 106082 112226
rect 106138 112170 136678 112226
rect 136734 112170 136802 112226
rect 136858 112170 167398 112226
rect 167454 112170 167522 112226
rect 167578 112170 198118 112226
rect 198174 112170 198242 112226
rect 198298 112170 228838 112226
rect 228894 112170 228962 112226
rect 229018 112170 259558 112226
rect 259614 112170 259682 112226
rect 259738 112170 281994 112226
rect 282050 112170 282118 112226
rect 282174 112170 282242 112226
rect 282298 112170 282366 112226
rect 282422 112170 312714 112226
rect 312770 112170 312838 112226
rect 312894 112170 312962 112226
rect 313018 112170 313086 112226
rect 313142 112170 343434 112226
rect 343490 112170 343558 112226
rect 343614 112170 343682 112226
rect 343738 112170 343806 112226
rect 343862 112170 364518 112226
rect 364574 112170 364642 112226
rect 364698 112170 395238 112226
rect 395294 112170 395362 112226
rect 395418 112170 435594 112226
rect 435650 112170 435718 112226
rect 435774 112170 435842 112226
rect 435898 112170 435966 112226
rect 436022 112170 464518 112226
rect 464574 112170 464642 112226
rect 464698 112170 495238 112226
rect 495294 112170 495362 112226
rect 495418 112170 525958 112226
rect 526014 112170 526082 112226
rect 526138 112170 556678 112226
rect 556734 112170 556802 112226
rect 556858 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597980 112226
rect -1916 112102 597980 112170
rect -1916 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 36234 112102
rect 36290 112046 36358 112102
rect 36414 112046 36482 112102
rect 36538 112046 36606 112102
rect 36662 112046 44518 112102
rect 44574 112046 44642 112102
rect 44698 112046 75238 112102
rect 75294 112046 75362 112102
rect 75418 112046 105958 112102
rect 106014 112046 106082 112102
rect 106138 112046 136678 112102
rect 136734 112046 136802 112102
rect 136858 112046 167398 112102
rect 167454 112046 167522 112102
rect 167578 112046 198118 112102
rect 198174 112046 198242 112102
rect 198298 112046 228838 112102
rect 228894 112046 228962 112102
rect 229018 112046 259558 112102
rect 259614 112046 259682 112102
rect 259738 112046 281994 112102
rect 282050 112046 282118 112102
rect 282174 112046 282242 112102
rect 282298 112046 282366 112102
rect 282422 112046 312714 112102
rect 312770 112046 312838 112102
rect 312894 112046 312962 112102
rect 313018 112046 313086 112102
rect 313142 112046 343434 112102
rect 343490 112046 343558 112102
rect 343614 112046 343682 112102
rect 343738 112046 343806 112102
rect 343862 112046 364518 112102
rect 364574 112046 364642 112102
rect 364698 112046 395238 112102
rect 395294 112046 395362 112102
rect 395418 112046 435594 112102
rect 435650 112046 435718 112102
rect 435774 112046 435842 112102
rect 435898 112046 435966 112102
rect 436022 112046 464518 112102
rect 464574 112046 464642 112102
rect 464698 112046 495238 112102
rect 495294 112046 495362 112102
rect 495418 112046 525958 112102
rect 526014 112046 526082 112102
rect 526138 112046 556678 112102
rect 556734 112046 556802 112102
rect 556858 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597980 112102
rect -1916 111978 597980 112046
rect -1916 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 36234 111978
rect 36290 111922 36358 111978
rect 36414 111922 36482 111978
rect 36538 111922 36606 111978
rect 36662 111922 44518 111978
rect 44574 111922 44642 111978
rect 44698 111922 75238 111978
rect 75294 111922 75362 111978
rect 75418 111922 105958 111978
rect 106014 111922 106082 111978
rect 106138 111922 136678 111978
rect 136734 111922 136802 111978
rect 136858 111922 167398 111978
rect 167454 111922 167522 111978
rect 167578 111922 198118 111978
rect 198174 111922 198242 111978
rect 198298 111922 228838 111978
rect 228894 111922 228962 111978
rect 229018 111922 259558 111978
rect 259614 111922 259682 111978
rect 259738 111922 281994 111978
rect 282050 111922 282118 111978
rect 282174 111922 282242 111978
rect 282298 111922 282366 111978
rect 282422 111922 312714 111978
rect 312770 111922 312838 111978
rect 312894 111922 312962 111978
rect 313018 111922 313086 111978
rect 313142 111922 343434 111978
rect 343490 111922 343558 111978
rect 343614 111922 343682 111978
rect 343738 111922 343806 111978
rect 343862 111922 364518 111978
rect 364574 111922 364642 111978
rect 364698 111922 395238 111978
rect 395294 111922 395362 111978
rect 395418 111922 435594 111978
rect 435650 111922 435718 111978
rect 435774 111922 435842 111978
rect 435898 111922 435966 111978
rect 436022 111922 464518 111978
rect 464574 111922 464642 111978
rect 464698 111922 495238 111978
rect 495294 111922 495362 111978
rect 495418 111922 525958 111978
rect 526014 111922 526082 111978
rect 526138 111922 556678 111978
rect 556734 111922 556802 111978
rect 556858 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597980 111978
rect -1916 111826 597980 111922
rect -1916 100350 597980 100446
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 9234 100350
rect 9290 100294 9358 100350
rect 9414 100294 9482 100350
rect 9538 100294 9606 100350
rect 9662 100294 39954 100350
rect 40010 100294 40078 100350
rect 40134 100294 40202 100350
rect 40258 100294 40326 100350
rect 40382 100294 59878 100350
rect 59934 100294 60002 100350
rect 60058 100294 90598 100350
rect 90654 100294 90722 100350
rect 90778 100294 121318 100350
rect 121374 100294 121442 100350
rect 121498 100294 152038 100350
rect 152094 100294 152162 100350
rect 152218 100294 182758 100350
rect 182814 100294 182882 100350
rect 182938 100294 213478 100350
rect 213534 100294 213602 100350
rect 213658 100294 244198 100350
rect 244254 100294 244322 100350
rect 244378 100294 285714 100350
rect 285770 100294 285838 100350
rect 285894 100294 285962 100350
rect 286018 100294 286086 100350
rect 286142 100294 316434 100350
rect 316490 100294 316558 100350
rect 316614 100294 316682 100350
rect 316738 100294 316806 100350
rect 316862 100294 347154 100350
rect 347210 100294 347278 100350
rect 347334 100294 347402 100350
rect 347458 100294 347526 100350
rect 347582 100294 379878 100350
rect 379934 100294 380002 100350
rect 380058 100294 410598 100350
rect 410654 100294 410722 100350
rect 410778 100294 439314 100350
rect 439370 100294 439438 100350
rect 439494 100294 439562 100350
rect 439618 100294 439686 100350
rect 439742 100294 479878 100350
rect 479934 100294 480002 100350
rect 480058 100294 510598 100350
rect 510654 100294 510722 100350
rect 510778 100294 541318 100350
rect 541374 100294 541442 100350
rect 541498 100294 562194 100350
rect 562250 100294 562318 100350
rect 562374 100294 562442 100350
rect 562498 100294 562566 100350
rect 562622 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect -1916 100226 597980 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 9234 100226
rect 9290 100170 9358 100226
rect 9414 100170 9482 100226
rect 9538 100170 9606 100226
rect 9662 100170 39954 100226
rect 40010 100170 40078 100226
rect 40134 100170 40202 100226
rect 40258 100170 40326 100226
rect 40382 100170 59878 100226
rect 59934 100170 60002 100226
rect 60058 100170 90598 100226
rect 90654 100170 90722 100226
rect 90778 100170 121318 100226
rect 121374 100170 121442 100226
rect 121498 100170 152038 100226
rect 152094 100170 152162 100226
rect 152218 100170 182758 100226
rect 182814 100170 182882 100226
rect 182938 100170 213478 100226
rect 213534 100170 213602 100226
rect 213658 100170 244198 100226
rect 244254 100170 244322 100226
rect 244378 100170 285714 100226
rect 285770 100170 285838 100226
rect 285894 100170 285962 100226
rect 286018 100170 286086 100226
rect 286142 100170 316434 100226
rect 316490 100170 316558 100226
rect 316614 100170 316682 100226
rect 316738 100170 316806 100226
rect 316862 100170 347154 100226
rect 347210 100170 347278 100226
rect 347334 100170 347402 100226
rect 347458 100170 347526 100226
rect 347582 100170 379878 100226
rect 379934 100170 380002 100226
rect 380058 100170 410598 100226
rect 410654 100170 410722 100226
rect 410778 100170 439314 100226
rect 439370 100170 439438 100226
rect 439494 100170 439562 100226
rect 439618 100170 439686 100226
rect 439742 100170 479878 100226
rect 479934 100170 480002 100226
rect 480058 100170 510598 100226
rect 510654 100170 510722 100226
rect 510778 100170 541318 100226
rect 541374 100170 541442 100226
rect 541498 100170 562194 100226
rect 562250 100170 562318 100226
rect 562374 100170 562442 100226
rect 562498 100170 562566 100226
rect 562622 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect -1916 100102 597980 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 9234 100102
rect 9290 100046 9358 100102
rect 9414 100046 9482 100102
rect 9538 100046 9606 100102
rect 9662 100046 39954 100102
rect 40010 100046 40078 100102
rect 40134 100046 40202 100102
rect 40258 100046 40326 100102
rect 40382 100046 59878 100102
rect 59934 100046 60002 100102
rect 60058 100046 90598 100102
rect 90654 100046 90722 100102
rect 90778 100046 121318 100102
rect 121374 100046 121442 100102
rect 121498 100046 152038 100102
rect 152094 100046 152162 100102
rect 152218 100046 182758 100102
rect 182814 100046 182882 100102
rect 182938 100046 213478 100102
rect 213534 100046 213602 100102
rect 213658 100046 244198 100102
rect 244254 100046 244322 100102
rect 244378 100046 285714 100102
rect 285770 100046 285838 100102
rect 285894 100046 285962 100102
rect 286018 100046 286086 100102
rect 286142 100046 316434 100102
rect 316490 100046 316558 100102
rect 316614 100046 316682 100102
rect 316738 100046 316806 100102
rect 316862 100046 347154 100102
rect 347210 100046 347278 100102
rect 347334 100046 347402 100102
rect 347458 100046 347526 100102
rect 347582 100046 379878 100102
rect 379934 100046 380002 100102
rect 380058 100046 410598 100102
rect 410654 100046 410722 100102
rect 410778 100046 439314 100102
rect 439370 100046 439438 100102
rect 439494 100046 439562 100102
rect 439618 100046 439686 100102
rect 439742 100046 479878 100102
rect 479934 100046 480002 100102
rect 480058 100046 510598 100102
rect 510654 100046 510722 100102
rect 510778 100046 541318 100102
rect 541374 100046 541442 100102
rect 541498 100046 562194 100102
rect 562250 100046 562318 100102
rect 562374 100046 562442 100102
rect 562498 100046 562566 100102
rect 562622 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect -1916 99978 597980 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 9234 99978
rect 9290 99922 9358 99978
rect 9414 99922 9482 99978
rect 9538 99922 9606 99978
rect 9662 99922 39954 99978
rect 40010 99922 40078 99978
rect 40134 99922 40202 99978
rect 40258 99922 40326 99978
rect 40382 99922 59878 99978
rect 59934 99922 60002 99978
rect 60058 99922 90598 99978
rect 90654 99922 90722 99978
rect 90778 99922 121318 99978
rect 121374 99922 121442 99978
rect 121498 99922 152038 99978
rect 152094 99922 152162 99978
rect 152218 99922 182758 99978
rect 182814 99922 182882 99978
rect 182938 99922 213478 99978
rect 213534 99922 213602 99978
rect 213658 99922 244198 99978
rect 244254 99922 244322 99978
rect 244378 99922 285714 99978
rect 285770 99922 285838 99978
rect 285894 99922 285962 99978
rect 286018 99922 286086 99978
rect 286142 99922 316434 99978
rect 316490 99922 316558 99978
rect 316614 99922 316682 99978
rect 316738 99922 316806 99978
rect 316862 99922 347154 99978
rect 347210 99922 347278 99978
rect 347334 99922 347402 99978
rect 347458 99922 347526 99978
rect 347582 99922 379878 99978
rect 379934 99922 380002 99978
rect 380058 99922 410598 99978
rect 410654 99922 410722 99978
rect 410778 99922 439314 99978
rect 439370 99922 439438 99978
rect 439494 99922 439562 99978
rect 439618 99922 439686 99978
rect 439742 99922 479878 99978
rect 479934 99922 480002 99978
rect 480058 99922 510598 99978
rect 510654 99922 510722 99978
rect 510778 99922 541318 99978
rect 541374 99922 541442 99978
rect 541498 99922 562194 99978
rect 562250 99922 562318 99978
rect 562374 99922 562442 99978
rect 562498 99922 562566 99978
rect 562622 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect -1916 99826 597980 99922
rect -1916 94350 597980 94446
rect -1916 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 36234 94350
rect 36290 94294 36358 94350
rect 36414 94294 36482 94350
rect 36538 94294 36606 94350
rect 36662 94294 44518 94350
rect 44574 94294 44642 94350
rect 44698 94294 75238 94350
rect 75294 94294 75362 94350
rect 75418 94294 105958 94350
rect 106014 94294 106082 94350
rect 106138 94294 136678 94350
rect 136734 94294 136802 94350
rect 136858 94294 167398 94350
rect 167454 94294 167522 94350
rect 167578 94294 198118 94350
rect 198174 94294 198242 94350
rect 198298 94294 228838 94350
rect 228894 94294 228962 94350
rect 229018 94294 259558 94350
rect 259614 94294 259682 94350
rect 259738 94294 281994 94350
rect 282050 94294 282118 94350
rect 282174 94294 282242 94350
rect 282298 94294 282366 94350
rect 282422 94294 312714 94350
rect 312770 94294 312838 94350
rect 312894 94294 312962 94350
rect 313018 94294 313086 94350
rect 313142 94294 343434 94350
rect 343490 94294 343558 94350
rect 343614 94294 343682 94350
rect 343738 94294 343806 94350
rect 343862 94294 364518 94350
rect 364574 94294 364642 94350
rect 364698 94294 395238 94350
rect 395294 94294 395362 94350
rect 395418 94294 435594 94350
rect 435650 94294 435718 94350
rect 435774 94294 435842 94350
rect 435898 94294 435966 94350
rect 436022 94294 464518 94350
rect 464574 94294 464642 94350
rect 464698 94294 495238 94350
rect 495294 94294 495362 94350
rect 495418 94294 525958 94350
rect 526014 94294 526082 94350
rect 526138 94294 556678 94350
rect 556734 94294 556802 94350
rect 556858 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597980 94350
rect -1916 94226 597980 94294
rect -1916 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 36234 94226
rect 36290 94170 36358 94226
rect 36414 94170 36482 94226
rect 36538 94170 36606 94226
rect 36662 94170 44518 94226
rect 44574 94170 44642 94226
rect 44698 94170 75238 94226
rect 75294 94170 75362 94226
rect 75418 94170 105958 94226
rect 106014 94170 106082 94226
rect 106138 94170 136678 94226
rect 136734 94170 136802 94226
rect 136858 94170 167398 94226
rect 167454 94170 167522 94226
rect 167578 94170 198118 94226
rect 198174 94170 198242 94226
rect 198298 94170 228838 94226
rect 228894 94170 228962 94226
rect 229018 94170 259558 94226
rect 259614 94170 259682 94226
rect 259738 94170 281994 94226
rect 282050 94170 282118 94226
rect 282174 94170 282242 94226
rect 282298 94170 282366 94226
rect 282422 94170 312714 94226
rect 312770 94170 312838 94226
rect 312894 94170 312962 94226
rect 313018 94170 313086 94226
rect 313142 94170 343434 94226
rect 343490 94170 343558 94226
rect 343614 94170 343682 94226
rect 343738 94170 343806 94226
rect 343862 94170 364518 94226
rect 364574 94170 364642 94226
rect 364698 94170 395238 94226
rect 395294 94170 395362 94226
rect 395418 94170 435594 94226
rect 435650 94170 435718 94226
rect 435774 94170 435842 94226
rect 435898 94170 435966 94226
rect 436022 94170 464518 94226
rect 464574 94170 464642 94226
rect 464698 94170 495238 94226
rect 495294 94170 495362 94226
rect 495418 94170 525958 94226
rect 526014 94170 526082 94226
rect 526138 94170 556678 94226
rect 556734 94170 556802 94226
rect 556858 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597980 94226
rect -1916 94102 597980 94170
rect -1916 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 36234 94102
rect 36290 94046 36358 94102
rect 36414 94046 36482 94102
rect 36538 94046 36606 94102
rect 36662 94046 44518 94102
rect 44574 94046 44642 94102
rect 44698 94046 75238 94102
rect 75294 94046 75362 94102
rect 75418 94046 105958 94102
rect 106014 94046 106082 94102
rect 106138 94046 136678 94102
rect 136734 94046 136802 94102
rect 136858 94046 167398 94102
rect 167454 94046 167522 94102
rect 167578 94046 198118 94102
rect 198174 94046 198242 94102
rect 198298 94046 228838 94102
rect 228894 94046 228962 94102
rect 229018 94046 259558 94102
rect 259614 94046 259682 94102
rect 259738 94046 281994 94102
rect 282050 94046 282118 94102
rect 282174 94046 282242 94102
rect 282298 94046 282366 94102
rect 282422 94046 312714 94102
rect 312770 94046 312838 94102
rect 312894 94046 312962 94102
rect 313018 94046 313086 94102
rect 313142 94046 343434 94102
rect 343490 94046 343558 94102
rect 343614 94046 343682 94102
rect 343738 94046 343806 94102
rect 343862 94046 364518 94102
rect 364574 94046 364642 94102
rect 364698 94046 395238 94102
rect 395294 94046 395362 94102
rect 395418 94046 435594 94102
rect 435650 94046 435718 94102
rect 435774 94046 435842 94102
rect 435898 94046 435966 94102
rect 436022 94046 464518 94102
rect 464574 94046 464642 94102
rect 464698 94046 495238 94102
rect 495294 94046 495362 94102
rect 495418 94046 525958 94102
rect 526014 94046 526082 94102
rect 526138 94046 556678 94102
rect 556734 94046 556802 94102
rect 556858 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597980 94102
rect -1916 93978 597980 94046
rect -1916 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 36234 93978
rect 36290 93922 36358 93978
rect 36414 93922 36482 93978
rect 36538 93922 36606 93978
rect 36662 93922 44518 93978
rect 44574 93922 44642 93978
rect 44698 93922 75238 93978
rect 75294 93922 75362 93978
rect 75418 93922 105958 93978
rect 106014 93922 106082 93978
rect 106138 93922 136678 93978
rect 136734 93922 136802 93978
rect 136858 93922 167398 93978
rect 167454 93922 167522 93978
rect 167578 93922 198118 93978
rect 198174 93922 198242 93978
rect 198298 93922 228838 93978
rect 228894 93922 228962 93978
rect 229018 93922 259558 93978
rect 259614 93922 259682 93978
rect 259738 93922 281994 93978
rect 282050 93922 282118 93978
rect 282174 93922 282242 93978
rect 282298 93922 282366 93978
rect 282422 93922 312714 93978
rect 312770 93922 312838 93978
rect 312894 93922 312962 93978
rect 313018 93922 313086 93978
rect 313142 93922 343434 93978
rect 343490 93922 343558 93978
rect 343614 93922 343682 93978
rect 343738 93922 343806 93978
rect 343862 93922 364518 93978
rect 364574 93922 364642 93978
rect 364698 93922 395238 93978
rect 395294 93922 395362 93978
rect 395418 93922 435594 93978
rect 435650 93922 435718 93978
rect 435774 93922 435842 93978
rect 435898 93922 435966 93978
rect 436022 93922 464518 93978
rect 464574 93922 464642 93978
rect 464698 93922 495238 93978
rect 495294 93922 495362 93978
rect 495418 93922 525958 93978
rect 526014 93922 526082 93978
rect 526138 93922 556678 93978
rect 556734 93922 556802 93978
rect 556858 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597980 93978
rect -1916 93826 597980 93922
rect -1916 82350 597980 82446
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 9234 82350
rect 9290 82294 9358 82350
rect 9414 82294 9482 82350
rect 9538 82294 9606 82350
rect 9662 82294 39954 82350
rect 40010 82294 40078 82350
rect 40134 82294 40202 82350
rect 40258 82294 40326 82350
rect 40382 82294 59878 82350
rect 59934 82294 60002 82350
rect 60058 82294 90598 82350
rect 90654 82294 90722 82350
rect 90778 82294 121318 82350
rect 121374 82294 121442 82350
rect 121498 82294 152038 82350
rect 152094 82294 152162 82350
rect 152218 82294 182758 82350
rect 182814 82294 182882 82350
rect 182938 82294 213478 82350
rect 213534 82294 213602 82350
rect 213658 82294 244198 82350
rect 244254 82294 244322 82350
rect 244378 82294 285714 82350
rect 285770 82294 285838 82350
rect 285894 82294 285962 82350
rect 286018 82294 286086 82350
rect 286142 82294 347154 82350
rect 347210 82294 347278 82350
rect 347334 82294 347402 82350
rect 347458 82294 347526 82350
rect 347582 82294 379878 82350
rect 379934 82294 380002 82350
rect 380058 82294 410598 82350
rect 410654 82294 410722 82350
rect 410778 82294 439314 82350
rect 439370 82294 439438 82350
rect 439494 82294 439562 82350
rect 439618 82294 439686 82350
rect 439742 82294 479878 82350
rect 479934 82294 480002 82350
rect 480058 82294 510598 82350
rect 510654 82294 510722 82350
rect 510778 82294 541318 82350
rect 541374 82294 541442 82350
rect 541498 82294 562194 82350
rect 562250 82294 562318 82350
rect 562374 82294 562442 82350
rect 562498 82294 562566 82350
rect 562622 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect -1916 82226 597980 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 9234 82226
rect 9290 82170 9358 82226
rect 9414 82170 9482 82226
rect 9538 82170 9606 82226
rect 9662 82170 39954 82226
rect 40010 82170 40078 82226
rect 40134 82170 40202 82226
rect 40258 82170 40326 82226
rect 40382 82170 59878 82226
rect 59934 82170 60002 82226
rect 60058 82170 90598 82226
rect 90654 82170 90722 82226
rect 90778 82170 121318 82226
rect 121374 82170 121442 82226
rect 121498 82170 152038 82226
rect 152094 82170 152162 82226
rect 152218 82170 182758 82226
rect 182814 82170 182882 82226
rect 182938 82170 213478 82226
rect 213534 82170 213602 82226
rect 213658 82170 244198 82226
rect 244254 82170 244322 82226
rect 244378 82170 285714 82226
rect 285770 82170 285838 82226
rect 285894 82170 285962 82226
rect 286018 82170 286086 82226
rect 286142 82170 347154 82226
rect 347210 82170 347278 82226
rect 347334 82170 347402 82226
rect 347458 82170 347526 82226
rect 347582 82170 379878 82226
rect 379934 82170 380002 82226
rect 380058 82170 410598 82226
rect 410654 82170 410722 82226
rect 410778 82170 439314 82226
rect 439370 82170 439438 82226
rect 439494 82170 439562 82226
rect 439618 82170 439686 82226
rect 439742 82170 479878 82226
rect 479934 82170 480002 82226
rect 480058 82170 510598 82226
rect 510654 82170 510722 82226
rect 510778 82170 541318 82226
rect 541374 82170 541442 82226
rect 541498 82170 562194 82226
rect 562250 82170 562318 82226
rect 562374 82170 562442 82226
rect 562498 82170 562566 82226
rect 562622 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect -1916 82147 597980 82170
rect -1916 82102 299528 82147
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 9234 82102
rect 9290 82046 9358 82102
rect 9414 82046 9482 82102
rect 9538 82046 9606 82102
rect 9662 82046 39954 82102
rect 40010 82046 40078 82102
rect 40134 82046 40202 82102
rect 40258 82046 40326 82102
rect 40382 82046 59878 82102
rect 59934 82046 60002 82102
rect 60058 82046 90598 82102
rect 90654 82046 90722 82102
rect 90778 82046 121318 82102
rect 121374 82046 121442 82102
rect 121498 82046 152038 82102
rect 152094 82046 152162 82102
rect 152218 82046 182758 82102
rect 182814 82046 182882 82102
rect 182938 82046 213478 82102
rect 213534 82046 213602 82102
rect 213658 82046 244198 82102
rect 244254 82046 244322 82102
rect 244378 82046 285714 82102
rect 285770 82046 285838 82102
rect 285894 82046 285962 82102
rect 286018 82046 286086 82102
rect 286142 82091 299528 82102
rect 299584 82091 299632 82147
rect 299688 82091 299736 82147
rect 299792 82091 307844 82147
rect 307900 82091 307948 82147
rect 308004 82091 308052 82147
rect 308108 82091 316160 82147
rect 316216 82091 316264 82147
rect 316320 82091 316368 82147
rect 316424 82091 324476 82147
rect 324532 82091 324580 82147
rect 324636 82091 324684 82147
rect 324740 82102 597980 82147
rect 324740 82091 347154 82102
rect 286142 82046 347154 82091
rect 347210 82046 347278 82102
rect 347334 82046 347402 82102
rect 347458 82046 347526 82102
rect 347582 82046 379878 82102
rect 379934 82046 380002 82102
rect 380058 82046 410598 82102
rect 410654 82046 410722 82102
rect 410778 82046 439314 82102
rect 439370 82046 439438 82102
rect 439494 82046 439562 82102
rect 439618 82046 439686 82102
rect 439742 82046 479878 82102
rect 479934 82046 480002 82102
rect 480058 82046 510598 82102
rect 510654 82046 510722 82102
rect 510778 82046 541318 82102
rect 541374 82046 541442 82102
rect 541498 82046 562194 82102
rect 562250 82046 562318 82102
rect 562374 82046 562442 82102
rect 562498 82046 562566 82102
rect 562622 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect -1916 82043 597980 82046
rect -1916 81987 299528 82043
rect 299584 81987 299632 82043
rect 299688 81987 299736 82043
rect 299792 81987 307844 82043
rect 307900 81987 307948 82043
rect 308004 81987 308052 82043
rect 308108 81987 316160 82043
rect 316216 81987 316264 82043
rect 316320 81987 316368 82043
rect 316424 81987 324476 82043
rect 324532 81987 324580 82043
rect 324636 81987 324684 82043
rect 324740 81987 597980 82043
rect -1916 81978 597980 81987
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 9234 81978
rect 9290 81922 9358 81978
rect 9414 81922 9482 81978
rect 9538 81922 9606 81978
rect 9662 81922 39954 81978
rect 40010 81922 40078 81978
rect 40134 81922 40202 81978
rect 40258 81922 40326 81978
rect 40382 81922 59878 81978
rect 59934 81922 60002 81978
rect 60058 81922 90598 81978
rect 90654 81922 90722 81978
rect 90778 81922 121318 81978
rect 121374 81922 121442 81978
rect 121498 81922 152038 81978
rect 152094 81922 152162 81978
rect 152218 81922 182758 81978
rect 182814 81922 182882 81978
rect 182938 81922 213478 81978
rect 213534 81922 213602 81978
rect 213658 81922 244198 81978
rect 244254 81922 244322 81978
rect 244378 81922 285714 81978
rect 285770 81922 285838 81978
rect 285894 81922 285962 81978
rect 286018 81922 286086 81978
rect 286142 81939 347154 81978
rect 286142 81922 299528 81939
rect -1916 81883 299528 81922
rect 299584 81883 299632 81939
rect 299688 81883 299736 81939
rect 299792 81883 307844 81939
rect 307900 81883 307948 81939
rect 308004 81883 308052 81939
rect 308108 81883 316160 81939
rect 316216 81883 316264 81939
rect 316320 81883 316368 81939
rect 316424 81883 324476 81939
rect 324532 81883 324580 81939
rect 324636 81883 324684 81939
rect 324740 81922 347154 81939
rect 347210 81922 347278 81978
rect 347334 81922 347402 81978
rect 347458 81922 347526 81978
rect 347582 81922 379878 81978
rect 379934 81922 380002 81978
rect 380058 81922 410598 81978
rect 410654 81922 410722 81978
rect 410778 81922 439314 81978
rect 439370 81922 439438 81978
rect 439494 81922 439562 81978
rect 439618 81922 439686 81978
rect 439742 81922 479878 81978
rect 479934 81922 480002 81978
rect 480058 81922 510598 81978
rect 510654 81922 510722 81978
rect 510778 81922 541318 81978
rect 541374 81922 541442 81978
rect 541498 81922 562194 81978
rect 562250 81922 562318 81978
rect 562374 81922 562442 81978
rect 562498 81922 562566 81978
rect 562622 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 324740 81883 597980 81922
rect -1916 81826 597980 81883
rect -1916 76350 597980 76446
rect -1916 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 36234 76350
rect 36290 76294 36358 76350
rect 36414 76294 36482 76350
rect 36538 76294 36606 76350
rect 36662 76294 44518 76350
rect 44574 76294 44642 76350
rect 44698 76294 75238 76350
rect 75294 76294 75362 76350
rect 75418 76294 105958 76350
rect 106014 76294 106082 76350
rect 106138 76294 136678 76350
rect 136734 76294 136802 76350
rect 136858 76294 167398 76350
rect 167454 76294 167522 76350
rect 167578 76294 198118 76350
rect 198174 76294 198242 76350
rect 198298 76294 228838 76350
rect 228894 76294 228962 76350
rect 229018 76294 259558 76350
rect 259614 76294 259682 76350
rect 259738 76294 281994 76350
rect 282050 76294 282118 76350
rect 282174 76294 282242 76350
rect 282298 76294 282366 76350
rect 282422 76294 295412 76350
rect 295468 76294 295536 76350
rect 295592 76294 303728 76350
rect 303784 76294 303852 76350
rect 303908 76294 312044 76350
rect 312100 76294 312168 76350
rect 312224 76294 312714 76350
rect 312770 76294 312838 76350
rect 312894 76294 312962 76350
rect 313018 76294 313086 76350
rect 313142 76294 320360 76350
rect 320416 76294 320484 76350
rect 320540 76294 343434 76350
rect 343490 76294 343558 76350
rect 343614 76294 343682 76350
rect 343738 76294 343806 76350
rect 343862 76294 364518 76350
rect 364574 76294 364642 76350
rect 364698 76294 395238 76350
rect 395294 76294 395362 76350
rect 395418 76294 435594 76350
rect 435650 76294 435718 76350
rect 435774 76294 435842 76350
rect 435898 76294 435966 76350
rect 436022 76294 464518 76350
rect 464574 76294 464642 76350
rect 464698 76294 495238 76350
rect 495294 76294 495362 76350
rect 495418 76294 525958 76350
rect 526014 76294 526082 76350
rect 526138 76294 556678 76350
rect 556734 76294 556802 76350
rect 556858 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597980 76350
rect -1916 76226 597980 76294
rect -1916 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 36234 76226
rect 36290 76170 36358 76226
rect 36414 76170 36482 76226
rect 36538 76170 36606 76226
rect 36662 76170 44518 76226
rect 44574 76170 44642 76226
rect 44698 76170 75238 76226
rect 75294 76170 75362 76226
rect 75418 76170 105958 76226
rect 106014 76170 106082 76226
rect 106138 76170 136678 76226
rect 136734 76170 136802 76226
rect 136858 76170 167398 76226
rect 167454 76170 167522 76226
rect 167578 76170 198118 76226
rect 198174 76170 198242 76226
rect 198298 76170 228838 76226
rect 228894 76170 228962 76226
rect 229018 76170 259558 76226
rect 259614 76170 259682 76226
rect 259738 76170 281994 76226
rect 282050 76170 282118 76226
rect 282174 76170 282242 76226
rect 282298 76170 282366 76226
rect 282422 76170 295412 76226
rect 295468 76170 295536 76226
rect 295592 76170 303728 76226
rect 303784 76170 303852 76226
rect 303908 76170 312044 76226
rect 312100 76170 312168 76226
rect 312224 76170 312714 76226
rect 312770 76170 312838 76226
rect 312894 76170 312962 76226
rect 313018 76170 313086 76226
rect 313142 76170 320360 76226
rect 320416 76170 320484 76226
rect 320540 76170 343434 76226
rect 343490 76170 343558 76226
rect 343614 76170 343682 76226
rect 343738 76170 343806 76226
rect 343862 76170 364518 76226
rect 364574 76170 364642 76226
rect 364698 76170 395238 76226
rect 395294 76170 395362 76226
rect 395418 76170 435594 76226
rect 435650 76170 435718 76226
rect 435774 76170 435842 76226
rect 435898 76170 435966 76226
rect 436022 76170 464518 76226
rect 464574 76170 464642 76226
rect 464698 76170 495238 76226
rect 495294 76170 495362 76226
rect 495418 76170 525958 76226
rect 526014 76170 526082 76226
rect 526138 76170 556678 76226
rect 556734 76170 556802 76226
rect 556858 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597980 76226
rect -1916 76102 597980 76170
rect -1916 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 36234 76102
rect 36290 76046 36358 76102
rect 36414 76046 36482 76102
rect 36538 76046 36606 76102
rect 36662 76046 44518 76102
rect 44574 76046 44642 76102
rect 44698 76046 75238 76102
rect 75294 76046 75362 76102
rect 75418 76046 105958 76102
rect 106014 76046 106082 76102
rect 106138 76046 136678 76102
rect 136734 76046 136802 76102
rect 136858 76046 167398 76102
rect 167454 76046 167522 76102
rect 167578 76046 198118 76102
rect 198174 76046 198242 76102
rect 198298 76046 228838 76102
rect 228894 76046 228962 76102
rect 229018 76046 259558 76102
rect 259614 76046 259682 76102
rect 259738 76046 281994 76102
rect 282050 76046 282118 76102
rect 282174 76046 282242 76102
rect 282298 76046 282366 76102
rect 282422 76046 295412 76102
rect 295468 76046 295536 76102
rect 295592 76046 303728 76102
rect 303784 76046 303852 76102
rect 303908 76046 312044 76102
rect 312100 76046 312168 76102
rect 312224 76046 312714 76102
rect 312770 76046 312838 76102
rect 312894 76046 312962 76102
rect 313018 76046 313086 76102
rect 313142 76046 320360 76102
rect 320416 76046 320484 76102
rect 320540 76046 343434 76102
rect 343490 76046 343558 76102
rect 343614 76046 343682 76102
rect 343738 76046 343806 76102
rect 343862 76046 364518 76102
rect 364574 76046 364642 76102
rect 364698 76046 395238 76102
rect 395294 76046 395362 76102
rect 395418 76046 435594 76102
rect 435650 76046 435718 76102
rect 435774 76046 435842 76102
rect 435898 76046 435966 76102
rect 436022 76046 464518 76102
rect 464574 76046 464642 76102
rect 464698 76046 495238 76102
rect 495294 76046 495362 76102
rect 495418 76046 525958 76102
rect 526014 76046 526082 76102
rect 526138 76046 556678 76102
rect 556734 76046 556802 76102
rect 556858 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597980 76102
rect -1916 75978 597980 76046
rect -1916 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 36234 75978
rect 36290 75922 36358 75978
rect 36414 75922 36482 75978
rect 36538 75922 36606 75978
rect 36662 75922 44518 75978
rect 44574 75922 44642 75978
rect 44698 75922 75238 75978
rect 75294 75922 75362 75978
rect 75418 75922 105958 75978
rect 106014 75922 106082 75978
rect 106138 75922 136678 75978
rect 136734 75922 136802 75978
rect 136858 75922 167398 75978
rect 167454 75922 167522 75978
rect 167578 75922 198118 75978
rect 198174 75922 198242 75978
rect 198298 75922 228838 75978
rect 228894 75922 228962 75978
rect 229018 75922 259558 75978
rect 259614 75922 259682 75978
rect 259738 75922 281994 75978
rect 282050 75922 282118 75978
rect 282174 75922 282242 75978
rect 282298 75922 282366 75978
rect 282422 75922 295412 75978
rect 295468 75922 295536 75978
rect 295592 75922 303728 75978
rect 303784 75922 303852 75978
rect 303908 75922 312044 75978
rect 312100 75922 312168 75978
rect 312224 75922 312714 75978
rect 312770 75922 312838 75978
rect 312894 75922 312962 75978
rect 313018 75922 313086 75978
rect 313142 75922 320360 75978
rect 320416 75922 320484 75978
rect 320540 75922 343434 75978
rect 343490 75922 343558 75978
rect 343614 75922 343682 75978
rect 343738 75922 343806 75978
rect 343862 75922 364518 75978
rect 364574 75922 364642 75978
rect 364698 75922 395238 75978
rect 395294 75922 395362 75978
rect 395418 75922 435594 75978
rect 435650 75922 435718 75978
rect 435774 75922 435842 75978
rect 435898 75922 435966 75978
rect 436022 75922 464518 75978
rect 464574 75922 464642 75978
rect 464698 75922 495238 75978
rect 495294 75922 495362 75978
rect 495418 75922 525958 75978
rect 526014 75922 526082 75978
rect 526138 75922 556678 75978
rect 556734 75922 556802 75978
rect 556858 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597980 75978
rect -1916 75826 597980 75922
rect -1916 64350 597980 64446
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 9234 64350
rect 9290 64294 9358 64350
rect 9414 64294 9482 64350
rect 9538 64294 9606 64350
rect 9662 64294 39954 64350
rect 40010 64294 40078 64350
rect 40134 64294 40202 64350
rect 40258 64294 40326 64350
rect 40382 64294 59878 64350
rect 59934 64294 60002 64350
rect 60058 64294 90598 64350
rect 90654 64294 90722 64350
rect 90778 64294 121318 64350
rect 121374 64294 121442 64350
rect 121498 64294 152038 64350
rect 152094 64294 152162 64350
rect 152218 64294 182758 64350
rect 182814 64294 182882 64350
rect 182938 64294 213478 64350
rect 213534 64294 213602 64350
rect 213658 64294 244198 64350
rect 244254 64294 244322 64350
rect 244378 64294 285714 64350
rect 285770 64294 285838 64350
rect 285894 64294 285962 64350
rect 286018 64294 286086 64350
rect 286142 64294 299570 64350
rect 299626 64294 299694 64350
rect 299750 64294 307886 64350
rect 307942 64294 308010 64350
rect 308066 64294 316202 64350
rect 316258 64294 316326 64350
rect 316382 64294 324518 64350
rect 324574 64294 324642 64350
rect 324698 64294 347154 64350
rect 347210 64294 347278 64350
rect 347334 64294 347402 64350
rect 347458 64294 347526 64350
rect 347582 64294 379878 64350
rect 379934 64294 380002 64350
rect 380058 64294 410598 64350
rect 410654 64294 410722 64350
rect 410778 64294 439314 64350
rect 439370 64294 439438 64350
rect 439494 64294 439562 64350
rect 439618 64294 439686 64350
rect 439742 64294 479878 64350
rect 479934 64294 480002 64350
rect 480058 64294 510598 64350
rect 510654 64294 510722 64350
rect 510778 64294 541318 64350
rect 541374 64294 541442 64350
rect 541498 64294 562194 64350
rect 562250 64294 562318 64350
rect 562374 64294 562442 64350
rect 562498 64294 562566 64350
rect 562622 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect -1916 64226 597980 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 9234 64226
rect 9290 64170 9358 64226
rect 9414 64170 9482 64226
rect 9538 64170 9606 64226
rect 9662 64170 39954 64226
rect 40010 64170 40078 64226
rect 40134 64170 40202 64226
rect 40258 64170 40326 64226
rect 40382 64170 59878 64226
rect 59934 64170 60002 64226
rect 60058 64170 90598 64226
rect 90654 64170 90722 64226
rect 90778 64170 121318 64226
rect 121374 64170 121442 64226
rect 121498 64170 152038 64226
rect 152094 64170 152162 64226
rect 152218 64170 182758 64226
rect 182814 64170 182882 64226
rect 182938 64170 213478 64226
rect 213534 64170 213602 64226
rect 213658 64170 244198 64226
rect 244254 64170 244322 64226
rect 244378 64170 285714 64226
rect 285770 64170 285838 64226
rect 285894 64170 285962 64226
rect 286018 64170 286086 64226
rect 286142 64170 299570 64226
rect 299626 64170 299694 64226
rect 299750 64170 307886 64226
rect 307942 64170 308010 64226
rect 308066 64170 316202 64226
rect 316258 64170 316326 64226
rect 316382 64170 324518 64226
rect 324574 64170 324642 64226
rect 324698 64170 347154 64226
rect 347210 64170 347278 64226
rect 347334 64170 347402 64226
rect 347458 64170 347526 64226
rect 347582 64170 379878 64226
rect 379934 64170 380002 64226
rect 380058 64170 410598 64226
rect 410654 64170 410722 64226
rect 410778 64170 439314 64226
rect 439370 64170 439438 64226
rect 439494 64170 439562 64226
rect 439618 64170 439686 64226
rect 439742 64170 479878 64226
rect 479934 64170 480002 64226
rect 480058 64170 510598 64226
rect 510654 64170 510722 64226
rect 510778 64170 541318 64226
rect 541374 64170 541442 64226
rect 541498 64170 562194 64226
rect 562250 64170 562318 64226
rect 562374 64170 562442 64226
rect 562498 64170 562566 64226
rect 562622 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect -1916 64102 597980 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 9234 64102
rect 9290 64046 9358 64102
rect 9414 64046 9482 64102
rect 9538 64046 9606 64102
rect 9662 64046 39954 64102
rect 40010 64046 40078 64102
rect 40134 64046 40202 64102
rect 40258 64046 40326 64102
rect 40382 64046 59878 64102
rect 59934 64046 60002 64102
rect 60058 64046 90598 64102
rect 90654 64046 90722 64102
rect 90778 64046 121318 64102
rect 121374 64046 121442 64102
rect 121498 64046 152038 64102
rect 152094 64046 152162 64102
rect 152218 64046 182758 64102
rect 182814 64046 182882 64102
rect 182938 64046 213478 64102
rect 213534 64046 213602 64102
rect 213658 64046 244198 64102
rect 244254 64046 244322 64102
rect 244378 64046 285714 64102
rect 285770 64046 285838 64102
rect 285894 64046 285962 64102
rect 286018 64046 286086 64102
rect 286142 64046 299570 64102
rect 299626 64046 299694 64102
rect 299750 64046 307886 64102
rect 307942 64046 308010 64102
rect 308066 64046 316202 64102
rect 316258 64046 316326 64102
rect 316382 64046 324518 64102
rect 324574 64046 324642 64102
rect 324698 64046 347154 64102
rect 347210 64046 347278 64102
rect 347334 64046 347402 64102
rect 347458 64046 347526 64102
rect 347582 64046 379878 64102
rect 379934 64046 380002 64102
rect 380058 64046 410598 64102
rect 410654 64046 410722 64102
rect 410778 64046 439314 64102
rect 439370 64046 439438 64102
rect 439494 64046 439562 64102
rect 439618 64046 439686 64102
rect 439742 64046 479878 64102
rect 479934 64046 480002 64102
rect 480058 64046 510598 64102
rect 510654 64046 510722 64102
rect 510778 64046 541318 64102
rect 541374 64046 541442 64102
rect 541498 64046 562194 64102
rect 562250 64046 562318 64102
rect 562374 64046 562442 64102
rect 562498 64046 562566 64102
rect 562622 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect -1916 63978 597980 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 9234 63978
rect 9290 63922 9358 63978
rect 9414 63922 9482 63978
rect 9538 63922 9606 63978
rect 9662 63922 39954 63978
rect 40010 63922 40078 63978
rect 40134 63922 40202 63978
rect 40258 63922 40326 63978
rect 40382 63922 59878 63978
rect 59934 63922 60002 63978
rect 60058 63922 90598 63978
rect 90654 63922 90722 63978
rect 90778 63922 121318 63978
rect 121374 63922 121442 63978
rect 121498 63922 152038 63978
rect 152094 63922 152162 63978
rect 152218 63922 182758 63978
rect 182814 63922 182882 63978
rect 182938 63922 213478 63978
rect 213534 63922 213602 63978
rect 213658 63922 244198 63978
rect 244254 63922 244322 63978
rect 244378 63922 285714 63978
rect 285770 63922 285838 63978
rect 285894 63922 285962 63978
rect 286018 63922 286086 63978
rect 286142 63922 299570 63978
rect 299626 63922 299694 63978
rect 299750 63922 307886 63978
rect 307942 63922 308010 63978
rect 308066 63922 316202 63978
rect 316258 63922 316326 63978
rect 316382 63922 324518 63978
rect 324574 63922 324642 63978
rect 324698 63922 347154 63978
rect 347210 63922 347278 63978
rect 347334 63922 347402 63978
rect 347458 63922 347526 63978
rect 347582 63922 379878 63978
rect 379934 63922 380002 63978
rect 380058 63922 410598 63978
rect 410654 63922 410722 63978
rect 410778 63922 439314 63978
rect 439370 63922 439438 63978
rect 439494 63922 439562 63978
rect 439618 63922 439686 63978
rect 439742 63922 479878 63978
rect 479934 63922 480002 63978
rect 480058 63922 510598 63978
rect 510654 63922 510722 63978
rect 510778 63922 541318 63978
rect 541374 63922 541442 63978
rect 541498 63922 562194 63978
rect 562250 63922 562318 63978
rect 562374 63922 562442 63978
rect 562498 63922 562566 63978
rect 562622 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect -1916 63826 597980 63922
rect -1916 58350 597980 58446
rect -1916 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 36234 58350
rect 36290 58294 36358 58350
rect 36414 58294 36482 58350
rect 36538 58294 36606 58350
rect 36662 58294 44518 58350
rect 44574 58294 44642 58350
rect 44698 58294 75238 58350
rect 75294 58294 75362 58350
rect 75418 58294 105958 58350
rect 106014 58294 106082 58350
rect 106138 58294 136678 58350
rect 136734 58294 136802 58350
rect 136858 58294 167398 58350
rect 167454 58294 167522 58350
rect 167578 58294 198118 58350
rect 198174 58294 198242 58350
rect 198298 58294 228838 58350
rect 228894 58294 228962 58350
rect 229018 58294 259558 58350
rect 259614 58294 259682 58350
rect 259738 58294 281994 58350
rect 282050 58294 282118 58350
rect 282174 58294 282242 58350
rect 282298 58294 282366 58350
rect 282422 58294 295412 58350
rect 295468 58294 295536 58350
rect 295592 58294 303728 58350
rect 303784 58294 303852 58350
rect 303908 58294 312044 58350
rect 312100 58294 312168 58350
rect 312224 58294 312714 58350
rect 312770 58294 312838 58350
rect 312894 58294 312962 58350
rect 313018 58294 313086 58350
rect 313142 58294 320360 58350
rect 320416 58294 320484 58350
rect 320540 58294 343434 58350
rect 343490 58294 343558 58350
rect 343614 58294 343682 58350
rect 343738 58294 343806 58350
rect 343862 58294 364518 58350
rect 364574 58294 364642 58350
rect 364698 58294 395238 58350
rect 395294 58294 395362 58350
rect 395418 58294 435594 58350
rect 435650 58294 435718 58350
rect 435774 58294 435842 58350
rect 435898 58294 435966 58350
rect 436022 58294 464518 58350
rect 464574 58294 464642 58350
rect 464698 58294 495238 58350
rect 495294 58294 495362 58350
rect 495418 58294 525958 58350
rect 526014 58294 526082 58350
rect 526138 58294 556678 58350
rect 556734 58294 556802 58350
rect 556858 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597980 58350
rect -1916 58226 597980 58294
rect -1916 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 36234 58226
rect 36290 58170 36358 58226
rect 36414 58170 36482 58226
rect 36538 58170 36606 58226
rect 36662 58170 44518 58226
rect 44574 58170 44642 58226
rect 44698 58170 75238 58226
rect 75294 58170 75362 58226
rect 75418 58170 105958 58226
rect 106014 58170 106082 58226
rect 106138 58170 136678 58226
rect 136734 58170 136802 58226
rect 136858 58170 167398 58226
rect 167454 58170 167522 58226
rect 167578 58170 198118 58226
rect 198174 58170 198242 58226
rect 198298 58170 228838 58226
rect 228894 58170 228962 58226
rect 229018 58170 259558 58226
rect 259614 58170 259682 58226
rect 259738 58170 281994 58226
rect 282050 58170 282118 58226
rect 282174 58170 282242 58226
rect 282298 58170 282366 58226
rect 282422 58170 295412 58226
rect 295468 58170 295536 58226
rect 295592 58170 303728 58226
rect 303784 58170 303852 58226
rect 303908 58170 312044 58226
rect 312100 58170 312168 58226
rect 312224 58170 312714 58226
rect 312770 58170 312838 58226
rect 312894 58170 312962 58226
rect 313018 58170 313086 58226
rect 313142 58170 320360 58226
rect 320416 58170 320484 58226
rect 320540 58170 343434 58226
rect 343490 58170 343558 58226
rect 343614 58170 343682 58226
rect 343738 58170 343806 58226
rect 343862 58170 364518 58226
rect 364574 58170 364642 58226
rect 364698 58170 395238 58226
rect 395294 58170 395362 58226
rect 395418 58170 435594 58226
rect 435650 58170 435718 58226
rect 435774 58170 435842 58226
rect 435898 58170 435966 58226
rect 436022 58170 464518 58226
rect 464574 58170 464642 58226
rect 464698 58170 495238 58226
rect 495294 58170 495362 58226
rect 495418 58170 525958 58226
rect 526014 58170 526082 58226
rect 526138 58170 556678 58226
rect 556734 58170 556802 58226
rect 556858 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597980 58226
rect -1916 58102 597980 58170
rect -1916 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 36234 58102
rect 36290 58046 36358 58102
rect 36414 58046 36482 58102
rect 36538 58046 36606 58102
rect 36662 58046 44518 58102
rect 44574 58046 44642 58102
rect 44698 58046 75238 58102
rect 75294 58046 75362 58102
rect 75418 58046 105958 58102
rect 106014 58046 106082 58102
rect 106138 58046 136678 58102
rect 136734 58046 136802 58102
rect 136858 58046 167398 58102
rect 167454 58046 167522 58102
rect 167578 58046 198118 58102
rect 198174 58046 198242 58102
rect 198298 58046 228838 58102
rect 228894 58046 228962 58102
rect 229018 58046 259558 58102
rect 259614 58046 259682 58102
rect 259738 58046 281994 58102
rect 282050 58046 282118 58102
rect 282174 58046 282242 58102
rect 282298 58046 282366 58102
rect 282422 58046 295412 58102
rect 295468 58046 295536 58102
rect 295592 58046 303728 58102
rect 303784 58046 303852 58102
rect 303908 58046 312044 58102
rect 312100 58046 312168 58102
rect 312224 58046 312714 58102
rect 312770 58046 312838 58102
rect 312894 58046 312962 58102
rect 313018 58046 313086 58102
rect 313142 58046 320360 58102
rect 320416 58046 320484 58102
rect 320540 58046 343434 58102
rect 343490 58046 343558 58102
rect 343614 58046 343682 58102
rect 343738 58046 343806 58102
rect 343862 58046 364518 58102
rect 364574 58046 364642 58102
rect 364698 58046 395238 58102
rect 395294 58046 395362 58102
rect 395418 58046 435594 58102
rect 435650 58046 435718 58102
rect 435774 58046 435842 58102
rect 435898 58046 435966 58102
rect 436022 58046 464518 58102
rect 464574 58046 464642 58102
rect 464698 58046 495238 58102
rect 495294 58046 495362 58102
rect 495418 58046 525958 58102
rect 526014 58046 526082 58102
rect 526138 58046 556678 58102
rect 556734 58046 556802 58102
rect 556858 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597980 58102
rect -1916 57978 597980 58046
rect -1916 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 36234 57978
rect 36290 57922 36358 57978
rect 36414 57922 36482 57978
rect 36538 57922 36606 57978
rect 36662 57922 44518 57978
rect 44574 57922 44642 57978
rect 44698 57922 75238 57978
rect 75294 57922 75362 57978
rect 75418 57922 105958 57978
rect 106014 57922 106082 57978
rect 106138 57922 136678 57978
rect 136734 57922 136802 57978
rect 136858 57922 167398 57978
rect 167454 57922 167522 57978
rect 167578 57922 198118 57978
rect 198174 57922 198242 57978
rect 198298 57922 228838 57978
rect 228894 57922 228962 57978
rect 229018 57922 259558 57978
rect 259614 57922 259682 57978
rect 259738 57922 281994 57978
rect 282050 57922 282118 57978
rect 282174 57922 282242 57978
rect 282298 57922 282366 57978
rect 282422 57922 295412 57978
rect 295468 57922 295536 57978
rect 295592 57922 303728 57978
rect 303784 57922 303852 57978
rect 303908 57922 312044 57978
rect 312100 57922 312168 57978
rect 312224 57922 312714 57978
rect 312770 57922 312838 57978
rect 312894 57922 312962 57978
rect 313018 57922 313086 57978
rect 313142 57922 320360 57978
rect 320416 57922 320484 57978
rect 320540 57922 343434 57978
rect 343490 57922 343558 57978
rect 343614 57922 343682 57978
rect 343738 57922 343806 57978
rect 343862 57922 364518 57978
rect 364574 57922 364642 57978
rect 364698 57922 395238 57978
rect 395294 57922 395362 57978
rect 395418 57922 435594 57978
rect 435650 57922 435718 57978
rect 435774 57922 435842 57978
rect 435898 57922 435966 57978
rect 436022 57922 464518 57978
rect 464574 57922 464642 57978
rect 464698 57922 495238 57978
rect 495294 57922 495362 57978
rect 495418 57922 525958 57978
rect 526014 57922 526082 57978
rect 526138 57922 556678 57978
rect 556734 57922 556802 57978
rect 556858 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597980 57978
rect -1916 57826 597980 57922
rect -1916 46350 597980 46446
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 9234 46350
rect 9290 46294 9358 46350
rect 9414 46294 9482 46350
rect 9538 46294 9606 46350
rect 9662 46294 39954 46350
rect 40010 46294 40078 46350
rect 40134 46294 40202 46350
rect 40258 46294 40326 46350
rect 40382 46294 70674 46350
rect 70730 46294 70798 46350
rect 70854 46294 70922 46350
rect 70978 46294 71046 46350
rect 71102 46294 101394 46350
rect 101450 46294 101518 46350
rect 101574 46294 101642 46350
rect 101698 46294 101766 46350
rect 101822 46294 132114 46350
rect 132170 46294 132238 46350
rect 132294 46294 132362 46350
rect 132418 46294 132486 46350
rect 132542 46294 162834 46350
rect 162890 46294 162958 46350
rect 163014 46294 163082 46350
rect 163138 46294 163206 46350
rect 163262 46294 193554 46350
rect 193610 46294 193678 46350
rect 193734 46294 193802 46350
rect 193858 46294 193926 46350
rect 193982 46294 224274 46350
rect 224330 46294 224398 46350
rect 224454 46294 224522 46350
rect 224578 46294 224646 46350
rect 224702 46294 254994 46350
rect 255050 46294 255118 46350
rect 255174 46294 255242 46350
rect 255298 46294 255366 46350
rect 255422 46294 285714 46350
rect 285770 46294 285838 46350
rect 285894 46294 285962 46350
rect 286018 46294 286086 46350
rect 286142 46294 316434 46350
rect 316490 46294 316558 46350
rect 316614 46294 316682 46350
rect 316738 46294 316806 46350
rect 316862 46294 347154 46350
rect 347210 46294 347278 46350
rect 347334 46294 347402 46350
rect 347458 46294 347526 46350
rect 347582 46294 377874 46350
rect 377930 46294 377998 46350
rect 378054 46294 378122 46350
rect 378178 46294 378246 46350
rect 378302 46294 408594 46350
rect 408650 46294 408718 46350
rect 408774 46294 408842 46350
rect 408898 46294 408966 46350
rect 409022 46294 439314 46350
rect 439370 46294 439438 46350
rect 439494 46294 439562 46350
rect 439618 46294 439686 46350
rect 439742 46294 470034 46350
rect 470090 46294 470158 46350
rect 470214 46294 470282 46350
rect 470338 46294 470406 46350
rect 470462 46294 500754 46350
rect 500810 46294 500878 46350
rect 500934 46294 501002 46350
rect 501058 46294 501126 46350
rect 501182 46294 531474 46350
rect 531530 46294 531598 46350
rect 531654 46294 531722 46350
rect 531778 46294 531846 46350
rect 531902 46294 562194 46350
rect 562250 46294 562318 46350
rect 562374 46294 562442 46350
rect 562498 46294 562566 46350
rect 562622 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect -1916 46226 597980 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 9234 46226
rect 9290 46170 9358 46226
rect 9414 46170 9482 46226
rect 9538 46170 9606 46226
rect 9662 46170 39954 46226
rect 40010 46170 40078 46226
rect 40134 46170 40202 46226
rect 40258 46170 40326 46226
rect 40382 46170 70674 46226
rect 70730 46170 70798 46226
rect 70854 46170 70922 46226
rect 70978 46170 71046 46226
rect 71102 46170 101394 46226
rect 101450 46170 101518 46226
rect 101574 46170 101642 46226
rect 101698 46170 101766 46226
rect 101822 46170 132114 46226
rect 132170 46170 132238 46226
rect 132294 46170 132362 46226
rect 132418 46170 132486 46226
rect 132542 46170 162834 46226
rect 162890 46170 162958 46226
rect 163014 46170 163082 46226
rect 163138 46170 163206 46226
rect 163262 46170 193554 46226
rect 193610 46170 193678 46226
rect 193734 46170 193802 46226
rect 193858 46170 193926 46226
rect 193982 46170 224274 46226
rect 224330 46170 224398 46226
rect 224454 46170 224522 46226
rect 224578 46170 224646 46226
rect 224702 46170 254994 46226
rect 255050 46170 255118 46226
rect 255174 46170 255242 46226
rect 255298 46170 255366 46226
rect 255422 46170 285714 46226
rect 285770 46170 285838 46226
rect 285894 46170 285962 46226
rect 286018 46170 286086 46226
rect 286142 46170 316434 46226
rect 316490 46170 316558 46226
rect 316614 46170 316682 46226
rect 316738 46170 316806 46226
rect 316862 46170 347154 46226
rect 347210 46170 347278 46226
rect 347334 46170 347402 46226
rect 347458 46170 347526 46226
rect 347582 46170 377874 46226
rect 377930 46170 377998 46226
rect 378054 46170 378122 46226
rect 378178 46170 378246 46226
rect 378302 46170 408594 46226
rect 408650 46170 408718 46226
rect 408774 46170 408842 46226
rect 408898 46170 408966 46226
rect 409022 46170 439314 46226
rect 439370 46170 439438 46226
rect 439494 46170 439562 46226
rect 439618 46170 439686 46226
rect 439742 46170 470034 46226
rect 470090 46170 470158 46226
rect 470214 46170 470282 46226
rect 470338 46170 470406 46226
rect 470462 46170 500754 46226
rect 500810 46170 500878 46226
rect 500934 46170 501002 46226
rect 501058 46170 501126 46226
rect 501182 46170 531474 46226
rect 531530 46170 531598 46226
rect 531654 46170 531722 46226
rect 531778 46170 531846 46226
rect 531902 46170 562194 46226
rect 562250 46170 562318 46226
rect 562374 46170 562442 46226
rect 562498 46170 562566 46226
rect 562622 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect -1916 46102 597980 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 9234 46102
rect 9290 46046 9358 46102
rect 9414 46046 9482 46102
rect 9538 46046 9606 46102
rect 9662 46046 39954 46102
rect 40010 46046 40078 46102
rect 40134 46046 40202 46102
rect 40258 46046 40326 46102
rect 40382 46046 70674 46102
rect 70730 46046 70798 46102
rect 70854 46046 70922 46102
rect 70978 46046 71046 46102
rect 71102 46046 101394 46102
rect 101450 46046 101518 46102
rect 101574 46046 101642 46102
rect 101698 46046 101766 46102
rect 101822 46046 132114 46102
rect 132170 46046 132238 46102
rect 132294 46046 132362 46102
rect 132418 46046 132486 46102
rect 132542 46046 162834 46102
rect 162890 46046 162958 46102
rect 163014 46046 163082 46102
rect 163138 46046 163206 46102
rect 163262 46046 193554 46102
rect 193610 46046 193678 46102
rect 193734 46046 193802 46102
rect 193858 46046 193926 46102
rect 193982 46046 224274 46102
rect 224330 46046 224398 46102
rect 224454 46046 224522 46102
rect 224578 46046 224646 46102
rect 224702 46046 254994 46102
rect 255050 46046 255118 46102
rect 255174 46046 255242 46102
rect 255298 46046 255366 46102
rect 255422 46046 285714 46102
rect 285770 46046 285838 46102
rect 285894 46046 285962 46102
rect 286018 46046 286086 46102
rect 286142 46046 316434 46102
rect 316490 46046 316558 46102
rect 316614 46046 316682 46102
rect 316738 46046 316806 46102
rect 316862 46046 347154 46102
rect 347210 46046 347278 46102
rect 347334 46046 347402 46102
rect 347458 46046 347526 46102
rect 347582 46046 377874 46102
rect 377930 46046 377998 46102
rect 378054 46046 378122 46102
rect 378178 46046 378246 46102
rect 378302 46046 408594 46102
rect 408650 46046 408718 46102
rect 408774 46046 408842 46102
rect 408898 46046 408966 46102
rect 409022 46046 439314 46102
rect 439370 46046 439438 46102
rect 439494 46046 439562 46102
rect 439618 46046 439686 46102
rect 439742 46046 470034 46102
rect 470090 46046 470158 46102
rect 470214 46046 470282 46102
rect 470338 46046 470406 46102
rect 470462 46046 500754 46102
rect 500810 46046 500878 46102
rect 500934 46046 501002 46102
rect 501058 46046 501126 46102
rect 501182 46046 531474 46102
rect 531530 46046 531598 46102
rect 531654 46046 531722 46102
rect 531778 46046 531846 46102
rect 531902 46046 562194 46102
rect 562250 46046 562318 46102
rect 562374 46046 562442 46102
rect 562498 46046 562566 46102
rect 562622 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect -1916 45978 597980 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 9234 45978
rect 9290 45922 9358 45978
rect 9414 45922 9482 45978
rect 9538 45922 9606 45978
rect 9662 45922 39954 45978
rect 40010 45922 40078 45978
rect 40134 45922 40202 45978
rect 40258 45922 40326 45978
rect 40382 45922 70674 45978
rect 70730 45922 70798 45978
rect 70854 45922 70922 45978
rect 70978 45922 71046 45978
rect 71102 45922 101394 45978
rect 101450 45922 101518 45978
rect 101574 45922 101642 45978
rect 101698 45922 101766 45978
rect 101822 45922 132114 45978
rect 132170 45922 132238 45978
rect 132294 45922 132362 45978
rect 132418 45922 132486 45978
rect 132542 45922 162834 45978
rect 162890 45922 162958 45978
rect 163014 45922 163082 45978
rect 163138 45922 163206 45978
rect 163262 45922 193554 45978
rect 193610 45922 193678 45978
rect 193734 45922 193802 45978
rect 193858 45922 193926 45978
rect 193982 45922 224274 45978
rect 224330 45922 224398 45978
rect 224454 45922 224522 45978
rect 224578 45922 224646 45978
rect 224702 45922 254994 45978
rect 255050 45922 255118 45978
rect 255174 45922 255242 45978
rect 255298 45922 255366 45978
rect 255422 45922 285714 45978
rect 285770 45922 285838 45978
rect 285894 45922 285962 45978
rect 286018 45922 286086 45978
rect 286142 45922 316434 45978
rect 316490 45922 316558 45978
rect 316614 45922 316682 45978
rect 316738 45922 316806 45978
rect 316862 45922 347154 45978
rect 347210 45922 347278 45978
rect 347334 45922 347402 45978
rect 347458 45922 347526 45978
rect 347582 45922 377874 45978
rect 377930 45922 377998 45978
rect 378054 45922 378122 45978
rect 378178 45922 378246 45978
rect 378302 45922 408594 45978
rect 408650 45922 408718 45978
rect 408774 45922 408842 45978
rect 408898 45922 408966 45978
rect 409022 45922 439314 45978
rect 439370 45922 439438 45978
rect 439494 45922 439562 45978
rect 439618 45922 439686 45978
rect 439742 45922 470034 45978
rect 470090 45922 470158 45978
rect 470214 45922 470282 45978
rect 470338 45922 470406 45978
rect 470462 45922 500754 45978
rect 500810 45922 500878 45978
rect 500934 45922 501002 45978
rect 501058 45922 501126 45978
rect 501182 45922 531474 45978
rect 531530 45922 531598 45978
rect 531654 45922 531722 45978
rect 531778 45922 531846 45978
rect 531902 45922 562194 45978
rect 562250 45922 562318 45978
rect 562374 45922 562442 45978
rect 562498 45922 562566 45978
rect 562622 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect -1916 45826 597980 45922
rect -1916 40350 597980 40446
rect -1916 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 36234 40350
rect 36290 40294 36358 40350
rect 36414 40294 36482 40350
rect 36538 40294 36606 40350
rect 36662 40294 66954 40350
rect 67010 40294 67078 40350
rect 67134 40294 67202 40350
rect 67258 40294 67326 40350
rect 67382 40294 97674 40350
rect 97730 40294 97798 40350
rect 97854 40294 97922 40350
rect 97978 40294 98046 40350
rect 98102 40294 128394 40350
rect 128450 40294 128518 40350
rect 128574 40294 128642 40350
rect 128698 40294 128766 40350
rect 128822 40294 159114 40350
rect 159170 40294 159238 40350
rect 159294 40294 159362 40350
rect 159418 40294 159486 40350
rect 159542 40294 189834 40350
rect 189890 40294 189958 40350
rect 190014 40294 190082 40350
rect 190138 40294 190206 40350
rect 190262 40294 220554 40350
rect 220610 40294 220678 40350
rect 220734 40294 220802 40350
rect 220858 40294 220926 40350
rect 220982 40294 251274 40350
rect 251330 40294 251398 40350
rect 251454 40294 251522 40350
rect 251578 40294 251646 40350
rect 251702 40294 281994 40350
rect 282050 40294 282118 40350
rect 282174 40294 282242 40350
rect 282298 40294 282366 40350
rect 282422 40294 312714 40350
rect 312770 40294 312838 40350
rect 312894 40294 312962 40350
rect 313018 40294 313086 40350
rect 313142 40294 343434 40350
rect 343490 40294 343558 40350
rect 343614 40294 343682 40350
rect 343738 40294 343806 40350
rect 343862 40294 374154 40350
rect 374210 40294 374278 40350
rect 374334 40294 374402 40350
rect 374458 40294 374526 40350
rect 374582 40294 404874 40350
rect 404930 40294 404998 40350
rect 405054 40294 405122 40350
rect 405178 40294 405246 40350
rect 405302 40294 435594 40350
rect 435650 40294 435718 40350
rect 435774 40294 435842 40350
rect 435898 40294 435966 40350
rect 436022 40294 466314 40350
rect 466370 40294 466438 40350
rect 466494 40294 466562 40350
rect 466618 40294 466686 40350
rect 466742 40294 497034 40350
rect 497090 40294 497158 40350
rect 497214 40294 497282 40350
rect 497338 40294 497406 40350
rect 497462 40294 527754 40350
rect 527810 40294 527878 40350
rect 527934 40294 528002 40350
rect 528058 40294 528126 40350
rect 528182 40294 558474 40350
rect 558530 40294 558598 40350
rect 558654 40294 558722 40350
rect 558778 40294 558846 40350
rect 558902 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597980 40350
rect -1916 40226 597980 40294
rect -1916 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 36234 40226
rect 36290 40170 36358 40226
rect 36414 40170 36482 40226
rect 36538 40170 36606 40226
rect 36662 40170 66954 40226
rect 67010 40170 67078 40226
rect 67134 40170 67202 40226
rect 67258 40170 67326 40226
rect 67382 40170 97674 40226
rect 97730 40170 97798 40226
rect 97854 40170 97922 40226
rect 97978 40170 98046 40226
rect 98102 40170 128394 40226
rect 128450 40170 128518 40226
rect 128574 40170 128642 40226
rect 128698 40170 128766 40226
rect 128822 40170 159114 40226
rect 159170 40170 159238 40226
rect 159294 40170 159362 40226
rect 159418 40170 159486 40226
rect 159542 40170 189834 40226
rect 189890 40170 189958 40226
rect 190014 40170 190082 40226
rect 190138 40170 190206 40226
rect 190262 40170 220554 40226
rect 220610 40170 220678 40226
rect 220734 40170 220802 40226
rect 220858 40170 220926 40226
rect 220982 40170 251274 40226
rect 251330 40170 251398 40226
rect 251454 40170 251522 40226
rect 251578 40170 251646 40226
rect 251702 40170 281994 40226
rect 282050 40170 282118 40226
rect 282174 40170 282242 40226
rect 282298 40170 282366 40226
rect 282422 40170 312714 40226
rect 312770 40170 312838 40226
rect 312894 40170 312962 40226
rect 313018 40170 313086 40226
rect 313142 40170 343434 40226
rect 343490 40170 343558 40226
rect 343614 40170 343682 40226
rect 343738 40170 343806 40226
rect 343862 40170 374154 40226
rect 374210 40170 374278 40226
rect 374334 40170 374402 40226
rect 374458 40170 374526 40226
rect 374582 40170 404874 40226
rect 404930 40170 404998 40226
rect 405054 40170 405122 40226
rect 405178 40170 405246 40226
rect 405302 40170 435594 40226
rect 435650 40170 435718 40226
rect 435774 40170 435842 40226
rect 435898 40170 435966 40226
rect 436022 40170 466314 40226
rect 466370 40170 466438 40226
rect 466494 40170 466562 40226
rect 466618 40170 466686 40226
rect 466742 40170 497034 40226
rect 497090 40170 497158 40226
rect 497214 40170 497282 40226
rect 497338 40170 497406 40226
rect 497462 40170 527754 40226
rect 527810 40170 527878 40226
rect 527934 40170 528002 40226
rect 528058 40170 528126 40226
rect 528182 40170 558474 40226
rect 558530 40170 558598 40226
rect 558654 40170 558722 40226
rect 558778 40170 558846 40226
rect 558902 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597980 40226
rect -1916 40102 597980 40170
rect -1916 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 36234 40102
rect 36290 40046 36358 40102
rect 36414 40046 36482 40102
rect 36538 40046 36606 40102
rect 36662 40046 66954 40102
rect 67010 40046 67078 40102
rect 67134 40046 67202 40102
rect 67258 40046 67326 40102
rect 67382 40046 97674 40102
rect 97730 40046 97798 40102
rect 97854 40046 97922 40102
rect 97978 40046 98046 40102
rect 98102 40046 128394 40102
rect 128450 40046 128518 40102
rect 128574 40046 128642 40102
rect 128698 40046 128766 40102
rect 128822 40046 159114 40102
rect 159170 40046 159238 40102
rect 159294 40046 159362 40102
rect 159418 40046 159486 40102
rect 159542 40046 189834 40102
rect 189890 40046 189958 40102
rect 190014 40046 190082 40102
rect 190138 40046 190206 40102
rect 190262 40046 220554 40102
rect 220610 40046 220678 40102
rect 220734 40046 220802 40102
rect 220858 40046 220926 40102
rect 220982 40046 251274 40102
rect 251330 40046 251398 40102
rect 251454 40046 251522 40102
rect 251578 40046 251646 40102
rect 251702 40046 281994 40102
rect 282050 40046 282118 40102
rect 282174 40046 282242 40102
rect 282298 40046 282366 40102
rect 282422 40046 312714 40102
rect 312770 40046 312838 40102
rect 312894 40046 312962 40102
rect 313018 40046 313086 40102
rect 313142 40046 343434 40102
rect 343490 40046 343558 40102
rect 343614 40046 343682 40102
rect 343738 40046 343806 40102
rect 343862 40046 374154 40102
rect 374210 40046 374278 40102
rect 374334 40046 374402 40102
rect 374458 40046 374526 40102
rect 374582 40046 404874 40102
rect 404930 40046 404998 40102
rect 405054 40046 405122 40102
rect 405178 40046 405246 40102
rect 405302 40046 435594 40102
rect 435650 40046 435718 40102
rect 435774 40046 435842 40102
rect 435898 40046 435966 40102
rect 436022 40046 466314 40102
rect 466370 40046 466438 40102
rect 466494 40046 466562 40102
rect 466618 40046 466686 40102
rect 466742 40046 497034 40102
rect 497090 40046 497158 40102
rect 497214 40046 497282 40102
rect 497338 40046 497406 40102
rect 497462 40046 527754 40102
rect 527810 40046 527878 40102
rect 527934 40046 528002 40102
rect 528058 40046 528126 40102
rect 528182 40046 558474 40102
rect 558530 40046 558598 40102
rect 558654 40046 558722 40102
rect 558778 40046 558846 40102
rect 558902 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597980 40102
rect -1916 39978 597980 40046
rect -1916 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 36234 39978
rect 36290 39922 36358 39978
rect 36414 39922 36482 39978
rect 36538 39922 36606 39978
rect 36662 39922 66954 39978
rect 67010 39922 67078 39978
rect 67134 39922 67202 39978
rect 67258 39922 67326 39978
rect 67382 39922 97674 39978
rect 97730 39922 97798 39978
rect 97854 39922 97922 39978
rect 97978 39922 98046 39978
rect 98102 39922 128394 39978
rect 128450 39922 128518 39978
rect 128574 39922 128642 39978
rect 128698 39922 128766 39978
rect 128822 39922 159114 39978
rect 159170 39922 159238 39978
rect 159294 39922 159362 39978
rect 159418 39922 159486 39978
rect 159542 39922 189834 39978
rect 189890 39922 189958 39978
rect 190014 39922 190082 39978
rect 190138 39922 190206 39978
rect 190262 39922 220554 39978
rect 220610 39922 220678 39978
rect 220734 39922 220802 39978
rect 220858 39922 220926 39978
rect 220982 39922 251274 39978
rect 251330 39922 251398 39978
rect 251454 39922 251522 39978
rect 251578 39922 251646 39978
rect 251702 39922 281994 39978
rect 282050 39922 282118 39978
rect 282174 39922 282242 39978
rect 282298 39922 282366 39978
rect 282422 39922 312714 39978
rect 312770 39922 312838 39978
rect 312894 39922 312962 39978
rect 313018 39922 313086 39978
rect 313142 39922 343434 39978
rect 343490 39922 343558 39978
rect 343614 39922 343682 39978
rect 343738 39922 343806 39978
rect 343862 39922 374154 39978
rect 374210 39922 374278 39978
rect 374334 39922 374402 39978
rect 374458 39922 374526 39978
rect 374582 39922 404874 39978
rect 404930 39922 404998 39978
rect 405054 39922 405122 39978
rect 405178 39922 405246 39978
rect 405302 39922 435594 39978
rect 435650 39922 435718 39978
rect 435774 39922 435842 39978
rect 435898 39922 435966 39978
rect 436022 39922 466314 39978
rect 466370 39922 466438 39978
rect 466494 39922 466562 39978
rect 466618 39922 466686 39978
rect 466742 39922 497034 39978
rect 497090 39922 497158 39978
rect 497214 39922 497282 39978
rect 497338 39922 497406 39978
rect 497462 39922 527754 39978
rect 527810 39922 527878 39978
rect 527934 39922 528002 39978
rect 528058 39922 528126 39978
rect 528182 39922 558474 39978
rect 558530 39922 558598 39978
rect 558654 39922 558722 39978
rect 558778 39922 558846 39978
rect 558902 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597980 39978
rect -1916 39826 597980 39922
rect -1916 28350 597980 28446
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 9234 28350
rect 9290 28294 9358 28350
rect 9414 28294 9482 28350
rect 9538 28294 9606 28350
rect 9662 28294 39954 28350
rect 40010 28294 40078 28350
rect 40134 28294 40202 28350
rect 40258 28294 40326 28350
rect 40382 28294 70674 28350
rect 70730 28294 70798 28350
rect 70854 28294 70922 28350
rect 70978 28294 71046 28350
rect 71102 28294 101394 28350
rect 101450 28294 101518 28350
rect 101574 28294 101642 28350
rect 101698 28294 101766 28350
rect 101822 28294 132114 28350
rect 132170 28294 132238 28350
rect 132294 28294 132362 28350
rect 132418 28294 132486 28350
rect 132542 28294 162834 28350
rect 162890 28294 162958 28350
rect 163014 28294 163082 28350
rect 163138 28294 163206 28350
rect 163262 28294 193554 28350
rect 193610 28294 193678 28350
rect 193734 28294 193802 28350
rect 193858 28294 193926 28350
rect 193982 28294 224274 28350
rect 224330 28294 224398 28350
rect 224454 28294 224522 28350
rect 224578 28294 224646 28350
rect 224702 28294 254994 28350
rect 255050 28294 255118 28350
rect 255174 28294 255242 28350
rect 255298 28294 255366 28350
rect 255422 28294 285714 28350
rect 285770 28294 285838 28350
rect 285894 28294 285962 28350
rect 286018 28294 286086 28350
rect 286142 28294 316434 28350
rect 316490 28294 316558 28350
rect 316614 28294 316682 28350
rect 316738 28294 316806 28350
rect 316862 28294 347154 28350
rect 347210 28294 347278 28350
rect 347334 28294 347402 28350
rect 347458 28294 347526 28350
rect 347582 28294 377874 28350
rect 377930 28294 377998 28350
rect 378054 28294 378122 28350
rect 378178 28294 378246 28350
rect 378302 28294 408594 28350
rect 408650 28294 408718 28350
rect 408774 28294 408842 28350
rect 408898 28294 408966 28350
rect 409022 28294 439314 28350
rect 439370 28294 439438 28350
rect 439494 28294 439562 28350
rect 439618 28294 439686 28350
rect 439742 28294 470034 28350
rect 470090 28294 470158 28350
rect 470214 28294 470282 28350
rect 470338 28294 470406 28350
rect 470462 28294 500754 28350
rect 500810 28294 500878 28350
rect 500934 28294 501002 28350
rect 501058 28294 501126 28350
rect 501182 28294 531474 28350
rect 531530 28294 531598 28350
rect 531654 28294 531722 28350
rect 531778 28294 531846 28350
rect 531902 28294 562194 28350
rect 562250 28294 562318 28350
rect 562374 28294 562442 28350
rect 562498 28294 562566 28350
rect 562622 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect -1916 28226 597980 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 9234 28226
rect 9290 28170 9358 28226
rect 9414 28170 9482 28226
rect 9538 28170 9606 28226
rect 9662 28170 39954 28226
rect 40010 28170 40078 28226
rect 40134 28170 40202 28226
rect 40258 28170 40326 28226
rect 40382 28170 70674 28226
rect 70730 28170 70798 28226
rect 70854 28170 70922 28226
rect 70978 28170 71046 28226
rect 71102 28170 101394 28226
rect 101450 28170 101518 28226
rect 101574 28170 101642 28226
rect 101698 28170 101766 28226
rect 101822 28170 132114 28226
rect 132170 28170 132238 28226
rect 132294 28170 132362 28226
rect 132418 28170 132486 28226
rect 132542 28170 162834 28226
rect 162890 28170 162958 28226
rect 163014 28170 163082 28226
rect 163138 28170 163206 28226
rect 163262 28170 193554 28226
rect 193610 28170 193678 28226
rect 193734 28170 193802 28226
rect 193858 28170 193926 28226
rect 193982 28170 224274 28226
rect 224330 28170 224398 28226
rect 224454 28170 224522 28226
rect 224578 28170 224646 28226
rect 224702 28170 254994 28226
rect 255050 28170 255118 28226
rect 255174 28170 255242 28226
rect 255298 28170 255366 28226
rect 255422 28170 285714 28226
rect 285770 28170 285838 28226
rect 285894 28170 285962 28226
rect 286018 28170 286086 28226
rect 286142 28170 316434 28226
rect 316490 28170 316558 28226
rect 316614 28170 316682 28226
rect 316738 28170 316806 28226
rect 316862 28170 347154 28226
rect 347210 28170 347278 28226
rect 347334 28170 347402 28226
rect 347458 28170 347526 28226
rect 347582 28170 377874 28226
rect 377930 28170 377998 28226
rect 378054 28170 378122 28226
rect 378178 28170 378246 28226
rect 378302 28170 408594 28226
rect 408650 28170 408718 28226
rect 408774 28170 408842 28226
rect 408898 28170 408966 28226
rect 409022 28170 439314 28226
rect 439370 28170 439438 28226
rect 439494 28170 439562 28226
rect 439618 28170 439686 28226
rect 439742 28170 470034 28226
rect 470090 28170 470158 28226
rect 470214 28170 470282 28226
rect 470338 28170 470406 28226
rect 470462 28170 500754 28226
rect 500810 28170 500878 28226
rect 500934 28170 501002 28226
rect 501058 28170 501126 28226
rect 501182 28170 531474 28226
rect 531530 28170 531598 28226
rect 531654 28170 531722 28226
rect 531778 28170 531846 28226
rect 531902 28170 562194 28226
rect 562250 28170 562318 28226
rect 562374 28170 562442 28226
rect 562498 28170 562566 28226
rect 562622 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect -1916 28102 597980 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 9234 28102
rect 9290 28046 9358 28102
rect 9414 28046 9482 28102
rect 9538 28046 9606 28102
rect 9662 28046 39954 28102
rect 40010 28046 40078 28102
rect 40134 28046 40202 28102
rect 40258 28046 40326 28102
rect 40382 28046 70674 28102
rect 70730 28046 70798 28102
rect 70854 28046 70922 28102
rect 70978 28046 71046 28102
rect 71102 28046 101394 28102
rect 101450 28046 101518 28102
rect 101574 28046 101642 28102
rect 101698 28046 101766 28102
rect 101822 28046 132114 28102
rect 132170 28046 132238 28102
rect 132294 28046 132362 28102
rect 132418 28046 132486 28102
rect 132542 28046 162834 28102
rect 162890 28046 162958 28102
rect 163014 28046 163082 28102
rect 163138 28046 163206 28102
rect 163262 28046 193554 28102
rect 193610 28046 193678 28102
rect 193734 28046 193802 28102
rect 193858 28046 193926 28102
rect 193982 28046 224274 28102
rect 224330 28046 224398 28102
rect 224454 28046 224522 28102
rect 224578 28046 224646 28102
rect 224702 28046 254994 28102
rect 255050 28046 255118 28102
rect 255174 28046 255242 28102
rect 255298 28046 255366 28102
rect 255422 28046 285714 28102
rect 285770 28046 285838 28102
rect 285894 28046 285962 28102
rect 286018 28046 286086 28102
rect 286142 28046 316434 28102
rect 316490 28046 316558 28102
rect 316614 28046 316682 28102
rect 316738 28046 316806 28102
rect 316862 28046 347154 28102
rect 347210 28046 347278 28102
rect 347334 28046 347402 28102
rect 347458 28046 347526 28102
rect 347582 28046 377874 28102
rect 377930 28046 377998 28102
rect 378054 28046 378122 28102
rect 378178 28046 378246 28102
rect 378302 28046 408594 28102
rect 408650 28046 408718 28102
rect 408774 28046 408842 28102
rect 408898 28046 408966 28102
rect 409022 28046 439314 28102
rect 439370 28046 439438 28102
rect 439494 28046 439562 28102
rect 439618 28046 439686 28102
rect 439742 28046 470034 28102
rect 470090 28046 470158 28102
rect 470214 28046 470282 28102
rect 470338 28046 470406 28102
rect 470462 28046 500754 28102
rect 500810 28046 500878 28102
rect 500934 28046 501002 28102
rect 501058 28046 501126 28102
rect 501182 28046 531474 28102
rect 531530 28046 531598 28102
rect 531654 28046 531722 28102
rect 531778 28046 531846 28102
rect 531902 28046 562194 28102
rect 562250 28046 562318 28102
rect 562374 28046 562442 28102
rect 562498 28046 562566 28102
rect 562622 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect -1916 27978 597980 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 9234 27978
rect 9290 27922 9358 27978
rect 9414 27922 9482 27978
rect 9538 27922 9606 27978
rect 9662 27922 39954 27978
rect 40010 27922 40078 27978
rect 40134 27922 40202 27978
rect 40258 27922 40326 27978
rect 40382 27922 70674 27978
rect 70730 27922 70798 27978
rect 70854 27922 70922 27978
rect 70978 27922 71046 27978
rect 71102 27922 101394 27978
rect 101450 27922 101518 27978
rect 101574 27922 101642 27978
rect 101698 27922 101766 27978
rect 101822 27922 132114 27978
rect 132170 27922 132238 27978
rect 132294 27922 132362 27978
rect 132418 27922 132486 27978
rect 132542 27922 162834 27978
rect 162890 27922 162958 27978
rect 163014 27922 163082 27978
rect 163138 27922 163206 27978
rect 163262 27922 193554 27978
rect 193610 27922 193678 27978
rect 193734 27922 193802 27978
rect 193858 27922 193926 27978
rect 193982 27922 224274 27978
rect 224330 27922 224398 27978
rect 224454 27922 224522 27978
rect 224578 27922 224646 27978
rect 224702 27922 254994 27978
rect 255050 27922 255118 27978
rect 255174 27922 255242 27978
rect 255298 27922 255366 27978
rect 255422 27922 285714 27978
rect 285770 27922 285838 27978
rect 285894 27922 285962 27978
rect 286018 27922 286086 27978
rect 286142 27922 316434 27978
rect 316490 27922 316558 27978
rect 316614 27922 316682 27978
rect 316738 27922 316806 27978
rect 316862 27922 347154 27978
rect 347210 27922 347278 27978
rect 347334 27922 347402 27978
rect 347458 27922 347526 27978
rect 347582 27922 377874 27978
rect 377930 27922 377998 27978
rect 378054 27922 378122 27978
rect 378178 27922 378246 27978
rect 378302 27922 408594 27978
rect 408650 27922 408718 27978
rect 408774 27922 408842 27978
rect 408898 27922 408966 27978
rect 409022 27922 439314 27978
rect 439370 27922 439438 27978
rect 439494 27922 439562 27978
rect 439618 27922 439686 27978
rect 439742 27922 470034 27978
rect 470090 27922 470158 27978
rect 470214 27922 470282 27978
rect 470338 27922 470406 27978
rect 470462 27922 500754 27978
rect 500810 27922 500878 27978
rect 500934 27922 501002 27978
rect 501058 27922 501126 27978
rect 501182 27922 531474 27978
rect 531530 27922 531598 27978
rect 531654 27922 531722 27978
rect 531778 27922 531846 27978
rect 531902 27922 562194 27978
rect 562250 27922 562318 27978
rect 562374 27922 562442 27978
rect 562498 27922 562566 27978
rect 562622 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect -1916 27826 597980 27922
rect -1916 22350 597980 22446
rect -1916 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 36234 22350
rect 36290 22294 36358 22350
rect 36414 22294 36482 22350
rect 36538 22294 36606 22350
rect 36662 22294 66954 22350
rect 67010 22294 67078 22350
rect 67134 22294 67202 22350
rect 67258 22294 67326 22350
rect 67382 22294 97674 22350
rect 97730 22294 97798 22350
rect 97854 22294 97922 22350
rect 97978 22294 98046 22350
rect 98102 22294 128394 22350
rect 128450 22294 128518 22350
rect 128574 22294 128642 22350
rect 128698 22294 128766 22350
rect 128822 22294 159114 22350
rect 159170 22294 159238 22350
rect 159294 22294 159362 22350
rect 159418 22294 159486 22350
rect 159542 22294 189834 22350
rect 189890 22294 189958 22350
rect 190014 22294 190082 22350
rect 190138 22294 190206 22350
rect 190262 22294 220554 22350
rect 220610 22294 220678 22350
rect 220734 22294 220802 22350
rect 220858 22294 220926 22350
rect 220982 22294 251274 22350
rect 251330 22294 251398 22350
rect 251454 22294 251522 22350
rect 251578 22294 251646 22350
rect 251702 22294 281994 22350
rect 282050 22294 282118 22350
rect 282174 22294 282242 22350
rect 282298 22294 282366 22350
rect 282422 22294 312714 22350
rect 312770 22294 312838 22350
rect 312894 22294 312962 22350
rect 313018 22294 313086 22350
rect 313142 22294 343434 22350
rect 343490 22294 343558 22350
rect 343614 22294 343682 22350
rect 343738 22294 343806 22350
rect 343862 22294 374154 22350
rect 374210 22294 374278 22350
rect 374334 22294 374402 22350
rect 374458 22294 374526 22350
rect 374582 22294 404874 22350
rect 404930 22294 404998 22350
rect 405054 22294 405122 22350
rect 405178 22294 405246 22350
rect 405302 22294 435594 22350
rect 435650 22294 435718 22350
rect 435774 22294 435842 22350
rect 435898 22294 435966 22350
rect 436022 22294 466314 22350
rect 466370 22294 466438 22350
rect 466494 22294 466562 22350
rect 466618 22294 466686 22350
rect 466742 22294 497034 22350
rect 497090 22294 497158 22350
rect 497214 22294 497282 22350
rect 497338 22294 497406 22350
rect 497462 22294 527754 22350
rect 527810 22294 527878 22350
rect 527934 22294 528002 22350
rect 528058 22294 528126 22350
rect 528182 22294 558474 22350
rect 558530 22294 558598 22350
rect 558654 22294 558722 22350
rect 558778 22294 558846 22350
rect 558902 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597980 22350
rect -1916 22226 597980 22294
rect -1916 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 36234 22226
rect 36290 22170 36358 22226
rect 36414 22170 36482 22226
rect 36538 22170 36606 22226
rect 36662 22170 66954 22226
rect 67010 22170 67078 22226
rect 67134 22170 67202 22226
rect 67258 22170 67326 22226
rect 67382 22170 97674 22226
rect 97730 22170 97798 22226
rect 97854 22170 97922 22226
rect 97978 22170 98046 22226
rect 98102 22170 128394 22226
rect 128450 22170 128518 22226
rect 128574 22170 128642 22226
rect 128698 22170 128766 22226
rect 128822 22170 159114 22226
rect 159170 22170 159238 22226
rect 159294 22170 159362 22226
rect 159418 22170 159486 22226
rect 159542 22170 189834 22226
rect 189890 22170 189958 22226
rect 190014 22170 190082 22226
rect 190138 22170 190206 22226
rect 190262 22170 220554 22226
rect 220610 22170 220678 22226
rect 220734 22170 220802 22226
rect 220858 22170 220926 22226
rect 220982 22170 251274 22226
rect 251330 22170 251398 22226
rect 251454 22170 251522 22226
rect 251578 22170 251646 22226
rect 251702 22170 281994 22226
rect 282050 22170 282118 22226
rect 282174 22170 282242 22226
rect 282298 22170 282366 22226
rect 282422 22170 312714 22226
rect 312770 22170 312838 22226
rect 312894 22170 312962 22226
rect 313018 22170 313086 22226
rect 313142 22170 343434 22226
rect 343490 22170 343558 22226
rect 343614 22170 343682 22226
rect 343738 22170 343806 22226
rect 343862 22170 374154 22226
rect 374210 22170 374278 22226
rect 374334 22170 374402 22226
rect 374458 22170 374526 22226
rect 374582 22170 404874 22226
rect 404930 22170 404998 22226
rect 405054 22170 405122 22226
rect 405178 22170 405246 22226
rect 405302 22170 435594 22226
rect 435650 22170 435718 22226
rect 435774 22170 435842 22226
rect 435898 22170 435966 22226
rect 436022 22170 466314 22226
rect 466370 22170 466438 22226
rect 466494 22170 466562 22226
rect 466618 22170 466686 22226
rect 466742 22170 497034 22226
rect 497090 22170 497158 22226
rect 497214 22170 497282 22226
rect 497338 22170 497406 22226
rect 497462 22170 527754 22226
rect 527810 22170 527878 22226
rect 527934 22170 528002 22226
rect 528058 22170 528126 22226
rect 528182 22170 558474 22226
rect 558530 22170 558598 22226
rect 558654 22170 558722 22226
rect 558778 22170 558846 22226
rect 558902 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597980 22226
rect -1916 22102 597980 22170
rect -1916 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 36234 22102
rect 36290 22046 36358 22102
rect 36414 22046 36482 22102
rect 36538 22046 36606 22102
rect 36662 22046 66954 22102
rect 67010 22046 67078 22102
rect 67134 22046 67202 22102
rect 67258 22046 67326 22102
rect 67382 22046 97674 22102
rect 97730 22046 97798 22102
rect 97854 22046 97922 22102
rect 97978 22046 98046 22102
rect 98102 22046 128394 22102
rect 128450 22046 128518 22102
rect 128574 22046 128642 22102
rect 128698 22046 128766 22102
rect 128822 22046 159114 22102
rect 159170 22046 159238 22102
rect 159294 22046 159362 22102
rect 159418 22046 159486 22102
rect 159542 22046 189834 22102
rect 189890 22046 189958 22102
rect 190014 22046 190082 22102
rect 190138 22046 190206 22102
rect 190262 22046 220554 22102
rect 220610 22046 220678 22102
rect 220734 22046 220802 22102
rect 220858 22046 220926 22102
rect 220982 22046 251274 22102
rect 251330 22046 251398 22102
rect 251454 22046 251522 22102
rect 251578 22046 251646 22102
rect 251702 22046 281994 22102
rect 282050 22046 282118 22102
rect 282174 22046 282242 22102
rect 282298 22046 282366 22102
rect 282422 22046 312714 22102
rect 312770 22046 312838 22102
rect 312894 22046 312962 22102
rect 313018 22046 313086 22102
rect 313142 22046 343434 22102
rect 343490 22046 343558 22102
rect 343614 22046 343682 22102
rect 343738 22046 343806 22102
rect 343862 22046 374154 22102
rect 374210 22046 374278 22102
rect 374334 22046 374402 22102
rect 374458 22046 374526 22102
rect 374582 22046 404874 22102
rect 404930 22046 404998 22102
rect 405054 22046 405122 22102
rect 405178 22046 405246 22102
rect 405302 22046 435594 22102
rect 435650 22046 435718 22102
rect 435774 22046 435842 22102
rect 435898 22046 435966 22102
rect 436022 22046 466314 22102
rect 466370 22046 466438 22102
rect 466494 22046 466562 22102
rect 466618 22046 466686 22102
rect 466742 22046 497034 22102
rect 497090 22046 497158 22102
rect 497214 22046 497282 22102
rect 497338 22046 497406 22102
rect 497462 22046 527754 22102
rect 527810 22046 527878 22102
rect 527934 22046 528002 22102
rect 528058 22046 528126 22102
rect 528182 22046 558474 22102
rect 558530 22046 558598 22102
rect 558654 22046 558722 22102
rect 558778 22046 558846 22102
rect 558902 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597980 22102
rect -1916 21978 597980 22046
rect -1916 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 36234 21978
rect 36290 21922 36358 21978
rect 36414 21922 36482 21978
rect 36538 21922 36606 21978
rect 36662 21922 66954 21978
rect 67010 21922 67078 21978
rect 67134 21922 67202 21978
rect 67258 21922 67326 21978
rect 67382 21922 97674 21978
rect 97730 21922 97798 21978
rect 97854 21922 97922 21978
rect 97978 21922 98046 21978
rect 98102 21922 128394 21978
rect 128450 21922 128518 21978
rect 128574 21922 128642 21978
rect 128698 21922 128766 21978
rect 128822 21922 159114 21978
rect 159170 21922 159238 21978
rect 159294 21922 159362 21978
rect 159418 21922 159486 21978
rect 159542 21922 189834 21978
rect 189890 21922 189958 21978
rect 190014 21922 190082 21978
rect 190138 21922 190206 21978
rect 190262 21922 220554 21978
rect 220610 21922 220678 21978
rect 220734 21922 220802 21978
rect 220858 21922 220926 21978
rect 220982 21922 251274 21978
rect 251330 21922 251398 21978
rect 251454 21922 251522 21978
rect 251578 21922 251646 21978
rect 251702 21922 281994 21978
rect 282050 21922 282118 21978
rect 282174 21922 282242 21978
rect 282298 21922 282366 21978
rect 282422 21922 312714 21978
rect 312770 21922 312838 21978
rect 312894 21922 312962 21978
rect 313018 21922 313086 21978
rect 313142 21922 343434 21978
rect 343490 21922 343558 21978
rect 343614 21922 343682 21978
rect 343738 21922 343806 21978
rect 343862 21922 374154 21978
rect 374210 21922 374278 21978
rect 374334 21922 374402 21978
rect 374458 21922 374526 21978
rect 374582 21922 404874 21978
rect 404930 21922 404998 21978
rect 405054 21922 405122 21978
rect 405178 21922 405246 21978
rect 405302 21922 435594 21978
rect 435650 21922 435718 21978
rect 435774 21922 435842 21978
rect 435898 21922 435966 21978
rect 436022 21922 466314 21978
rect 466370 21922 466438 21978
rect 466494 21922 466562 21978
rect 466618 21922 466686 21978
rect 466742 21922 497034 21978
rect 497090 21922 497158 21978
rect 497214 21922 497282 21978
rect 497338 21922 497406 21978
rect 497462 21922 527754 21978
rect 527810 21922 527878 21978
rect 527934 21922 528002 21978
rect 528058 21922 528126 21978
rect 528182 21922 558474 21978
rect 558530 21922 558598 21978
rect 558654 21922 558722 21978
rect 558778 21922 558846 21978
rect 558902 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597980 21978
rect -1916 21826 597980 21922
rect -1916 10350 597980 10446
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 9234 10350
rect 9290 10294 9358 10350
rect 9414 10294 9482 10350
rect 9538 10294 9606 10350
rect 9662 10294 39954 10350
rect 40010 10294 40078 10350
rect 40134 10294 40202 10350
rect 40258 10294 40326 10350
rect 40382 10294 70674 10350
rect 70730 10294 70798 10350
rect 70854 10294 70922 10350
rect 70978 10294 71046 10350
rect 71102 10294 101394 10350
rect 101450 10294 101518 10350
rect 101574 10294 101642 10350
rect 101698 10294 101766 10350
rect 101822 10294 132114 10350
rect 132170 10294 132238 10350
rect 132294 10294 132362 10350
rect 132418 10294 132486 10350
rect 132542 10294 162834 10350
rect 162890 10294 162958 10350
rect 163014 10294 163082 10350
rect 163138 10294 163206 10350
rect 163262 10294 193554 10350
rect 193610 10294 193678 10350
rect 193734 10294 193802 10350
rect 193858 10294 193926 10350
rect 193982 10294 224274 10350
rect 224330 10294 224398 10350
rect 224454 10294 224522 10350
rect 224578 10294 224646 10350
rect 224702 10294 254994 10350
rect 255050 10294 255118 10350
rect 255174 10294 255242 10350
rect 255298 10294 255366 10350
rect 255422 10294 285714 10350
rect 285770 10294 285838 10350
rect 285894 10294 285962 10350
rect 286018 10294 286086 10350
rect 286142 10294 316434 10350
rect 316490 10294 316558 10350
rect 316614 10294 316682 10350
rect 316738 10294 316806 10350
rect 316862 10294 347154 10350
rect 347210 10294 347278 10350
rect 347334 10294 347402 10350
rect 347458 10294 347526 10350
rect 347582 10294 377874 10350
rect 377930 10294 377998 10350
rect 378054 10294 378122 10350
rect 378178 10294 378246 10350
rect 378302 10294 408594 10350
rect 408650 10294 408718 10350
rect 408774 10294 408842 10350
rect 408898 10294 408966 10350
rect 409022 10294 439314 10350
rect 439370 10294 439438 10350
rect 439494 10294 439562 10350
rect 439618 10294 439686 10350
rect 439742 10294 470034 10350
rect 470090 10294 470158 10350
rect 470214 10294 470282 10350
rect 470338 10294 470406 10350
rect 470462 10294 500754 10350
rect 500810 10294 500878 10350
rect 500934 10294 501002 10350
rect 501058 10294 501126 10350
rect 501182 10294 531474 10350
rect 531530 10294 531598 10350
rect 531654 10294 531722 10350
rect 531778 10294 531846 10350
rect 531902 10294 562194 10350
rect 562250 10294 562318 10350
rect 562374 10294 562442 10350
rect 562498 10294 562566 10350
rect 562622 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect -1916 10226 597980 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 9234 10226
rect 9290 10170 9358 10226
rect 9414 10170 9482 10226
rect 9538 10170 9606 10226
rect 9662 10170 39954 10226
rect 40010 10170 40078 10226
rect 40134 10170 40202 10226
rect 40258 10170 40326 10226
rect 40382 10170 70674 10226
rect 70730 10170 70798 10226
rect 70854 10170 70922 10226
rect 70978 10170 71046 10226
rect 71102 10170 101394 10226
rect 101450 10170 101518 10226
rect 101574 10170 101642 10226
rect 101698 10170 101766 10226
rect 101822 10170 132114 10226
rect 132170 10170 132238 10226
rect 132294 10170 132362 10226
rect 132418 10170 132486 10226
rect 132542 10170 162834 10226
rect 162890 10170 162958 10226
rect 163014 10170 163082 10226
rect 163138 10170 163206 10226
rect 163262 10170 193554 10226
rect 193610 10170 193678 10226
rect 193734 10170 193802 10226
rect 193858 10170 193926 10226
rect 193982 10170 224274 10226
rect 224330 10170 224398 10226
rect 224454 10170 224522 10226
rect 224578 10170 224646 10226
rect 224702 10170 254994 10226
rect 255050 10170 255118 10226
rect 255174 10170 255242 10226
rect 255298 10170 255366 10226
rect 255422 10170 285714 10226
rect 285770 10170 285838 10226
rect 285894 10170 285962 10226
rect 286018 10170 286086 10226
rect 286142 10170 316434 10226
rect 316490 10170 316558 10226
rect 316614 10170 316682 10226
rect 316738 10170 316806 10226
rect 316862 10170 347154 10226
rect 347210 10170 347278 10226
rect 347334 10170 347402 10226
rect 347458 10170 347526 10226
rect 347582 10170 377874 10226
rect 377930 10170 377998 10226
rect 378054 10170 378122 10226
rect 378178 10170 378246 10226
rect 378302 10170 408594 10226
rect 408650 10170 408718 10226
rect 408774 10170 408842 10226
rect 408898 10170 408966 10226
rect 409022 10170 439314 10226
rect 439370 10170 439438 10226
rect 439494 10170 439562 10226
rect 439618 10170 439686 10226
rect 439742 10170 470034 10226
rect 470090 10170 470158 10226
rect 470214 10170 470282 10226
rect 470338 10170 470406 10226
rect 470462 10170 500754 10226
rect 500810 10170 500878 10226
rect 500934 10170 501002 10226
rect 501058 10170 501126 10226
rect 501182 10170 531474 10226
rect 531530 10170 531598 10226
rect 531654 10170 531722 10226
rect 531778 10170 531846 10226
rect 531902 10170 562194 10226
rect 562250 10170 562318 10226
rect 562374 10170 562442 10226
rect 562498 10170 562566 10226
rect 562622 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect -1916 10102 597980 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 9234 10102
rect 9290 10046 9358 10102
rect 9414 10046 9482 10102
rect 9538 10046 9606 10102
rect 9662 10046 39954 10102
rect 40010 10046 40078 10102
rect 40134 10046 40202 10102
rect 40258 10046 40326 10102
rect 40382 10046 70674 10102
rect 70730 10046 70798 10102
rect 70854 10046 70922 10102
rect 70978 10046 71046 10102
rect 71102 10046 101394 10102
rect 101450 10046 101518 10102
rect 101574 10046 101642 10102
rect 101698 10046 101766 10102
rect 101822 10046 132114 10102
rect 132170 10046 132238 10102
rect 132294 10046 132362 10102
rect 132418 10046 132486 10102
rect 132542 10046 162834 10102
rect 162890 10046 162958 10102
rect 163014 10046 163082 10102
rect 163138 10046 163206 10102
rect 163262 10046 193554 10102
rect 193610 10046 193678 10102
rect 193734 10046 193802 10102
rect 193858 10046 193926 10102
rect 193982 10046 224274 10102
rect 224330 10046 224398 10102
rect 224454 10046 224522 10102
rect 224578 10046 224646 10102
rect 224702 10046 254994 10102
rect 255050 10046 255118 10102
rect 255174 10046 255242 10102
rect 255298 10046 255366 10102
rect 255422 10046 285714 10102
rect 285770 10046 285838 10102
rect 285894 10046 285962 10102
rect 286018 10046 286086 10102
rect 286142 10046 316434 10102
rect 316490 10046 316558 10102
rect 316614 10046 316682 10102
rect 316738 10046 316806 10102
rect 316862 10046 347154 10102
rect 347210 10046 347278 10102
rect 347334 10046 347402 10102
rect 347458 10046 347526 10102
rect 347582 10046 377874 10102
rect 377930 10046 377998 10102
rect 378054 10046 378122 10102
rect 378178 10046 378246 10102
rect 378302 10046 408594 10102
rect 408650 10046 408718 10102
rect 408774 10046 408842 10102
rect 408898 10046 408966 10102
rect 409022 10046 439314 10102
rect 439370 10046 439438 10102
rect 439494 10046 439562 10102
rect 439618 10046 439686 10102
rect 439742 10046 470034 10102
rect 470090 10046 470158 10102
rect 470214 10046 470282 10102
rect 470338 10046 470406 10102
rect 470462 10046 500754 10102
rect 500810 10046 500878 10102
rect 500934 10046 501002 10102
rect 501058 10046 501126 10102
rect 501182 10046 531474 10102
rect 531530 10046 531598 10102
rect 531654 10046 531722 10102
rect 531778 10046 531846 10102
rect 531902 10046 562194 10102
rect 562250 10046 562318 10102
rect 562374 10046 562442 10102
rect 562498 10046 562566 10102
rect 562622 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect -1916 9978 597980 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 9234 9978
rect 9290 9922 9358 9978
rect 9414 9922 9482 9978
rect 9538 9922 9606 9978
rect 9662 9922 39954 9978
rect 40010 9922 40078 9978
rect 40134 9922 40202 9978
rect 40258 9922 40326 9978
rect 40382 9922 70674 9978
rect 70730 9922 70798 9978
rect 70854 9922 70922 9978
rect 70978 9922 71046 9978
rect 71102 9922 101394 9978
rect 101450 9922 101518 9978
rect 101574 9922 101642 9978
rect 101698 9922 101766 9978
rect 101822 9922 132114 9978
rect 132170 9922 132238 9978
rect 132294 9922 132362 9978
rect 132418 9922 132486 9978
rect 132542 9922 162834 9978
rect 162890 9922 162958 9978
rect 163014 9922 163082 9978
rect 163138 9922 163206 9978
rect 163262 9922 193554 9978
rect 193610 9922 193678 9978
rect 193734 9922 193802 9978
rect 193858 9922 193926 9978
rect 193982 9922 224274 9978
rect 224330 9922 224398 9978
rect 224454 9922 224522 9978
rect 224578 9922 224646 9978
rect 224702 9922 254994 9978
rect 255050 9922 255118 9978
rect 255174 9922 255242 9978
rect 255298 9922 255366 9978
rect 255422 9922 285714 9978
rect 285770 9922 285838 9978
rect 285894 9922 285962 9978
rect 286018 9922 286086 9978
rect 286142 9922 316434 9978
rect 316490 9922 316558 9978
rect 316614 9922 316682 9978
rect 316738 9922 316806 9978
rect 316862 9922 347154 9978
rect 347210 9922 347278 9978
rect 347334 9922 347402 9978
rect 347458 9922 347526 9978
rect 347582 9922 377874 9978
rect 377930 9922 377998 9978
rect 378054 9922 378122 9978
rect 378178 9922 378246 9978
rect 378302 9922 408594 9978
rect 408650 9922 408718 9978
rect 408774 9922 408842 9978
rect 408898 9922 408966 9978
rect 409022 9922 439314 9978
rect 439370 9922 439438 9978
rect 439494 9922 439562 9978
rect 439618 9922 439686 9978
rect 439742 9922 470034 9978
rect 470090 9922 470158 9978
rect 470214 9922 470282 9978
rect 470338 9922 470406 9978
rect 470462 9922 500754 9978
rect 500810 9922 500878 9978
rect 500934 9922 501002 9978
rect 501058 9922 501126 9978
rect 501182 9922 531474 9978
rect 531530 9922 531598 9978
rect 531654 9922 531722 9978
rect 531778 9922 531846 9978
rect 531902 9922 562194 9978
rect 562250 9922 562318 9978
rect 562374 9922 562442 9978
rect 562498 9922 562566 9978
rect 562622 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect -1916 9826 597980 9922
rect -1916 4350 597980 4446
rect -1916 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597980 4350
rect -1916 4226 597980 4294
rect -1916 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597980 4226
rect -1916 4102 597980 4170
rect -1916 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597980 4102
rect -1916 3978 597980 4046
rect -1916 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597980 3978
rect -1916 3826 597980 3922
rect -956 -160 597020 -64
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect -956 -284 597020 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect -956 -408 597020 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect -956 -532 597020 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect -956 -684 597020 -588
rect -1916 -1120 597980 -1024
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 9234 -1120
rect 9290 -1176 9358 -1120
rect 9414 -1176 9482 -1120
rect 9538 -1176 9606 -1120
rect 9662 -1176 39954 -1120
rect 40010 -1176 40078 -1120
rect 40134 -1176 40202 -1120
rect 40258 -1176 40326 -1120
rect 40382 -1176 70674 -1120
rect 70730 -1176 70798 -1120
rect 70854 -1176 70922 -1120
rect 70978 -1176 71046 -1120
rect 71102 -1176 101394 -1120
rect 101450 -1176 101518 -1120
rect 101574 -1176 101642 -1120
rect 101698 -1176 101766 -1120
rect 101822 -1176 132114 -1120
rect 132170 -1176 132238 -1120
rect 132294 -1176 132362 -1120
rect 132418 -1176 132486 -1120
rect 132542 -1176 162834 -1120
rect 162890 -1176 162958 -1120
rect 163014 -1176 163082 -1120
rect 163138 -1176 163206 -1120
rect 163262 -1176 193554 -1120
rect 193610 -1176 193678 -1120
rect 193734 -1176 193802 -1120
rect 193858 -1176 193926 -1120
rect 193982 -1176 224274 -1120
rect 224330 -1176 224398 -1120
rect 224454 -1176 224522 -1120
rect 224578 -1176 224646 -1120
rect 224702 -1176 254994 -1120
rect 255050 -1176 255118 -1120
rect 255174 -1176 255242 -1120
rect 255298 -1176 255366 -1120
rect 255422 -1176 285714 -1120
rect 285770 -1176 285838 -1120
rect 285894 -1176 285962 -1120
rect 286018 -1176 286086 -1120
rect 286142 -1176 316434 -1120
rect 316490 -1176 316558 -1120
rect 316614 -1176 316682 -1120
rect 316738 -1176 316806 -1120
rect 316862 -1176 347154 -1120
rect 347210 -1176 347278 -1120
rect 347334 -1176 347402 -1120
rect 347458 -1176 347526 -1120
rect 347582 -1176 377874 -1120
rect 377930 -1176 377998 -1120
rect 378054 -1176 378122 -1120
rect 378178 -1176 378246 -1120
rect 378302 -1176 408594 -1120
rect 408650 -1176 408718 -1120
rect 408774 -1176 408842 -1120
rect 408898 -1176 408966 -1120
rect 409022 -1176 439314 -1120
rect 439370 -1176 439438 -1120
rect 439494 -1176 439562 -1120
rect 439618 -1176 439686 -1120
rect 439742 -1176 470034 -1120
rect 470090 -1176 470158 -1120
rect 470214 -1176 470282 -1120
rect 470338 -1176 470406 -1120
rect 470462 -1176 500754 -1120
rect 500810 -1176 500878 -1120
rect 500934 -1176 501002 -1120
rect 501058 -1176 501126 -1120
rect 501182 -1176 531474 -1120
rect 531530 -1176 531598 -1120
rect 531654 -1176 531722 -1120
rect 531778 -1176 531846 -1120
rect 531902 -1176 562194 -1120
rect 562250 -1176 562318 -1120
rect 562374 -1176 562442 -1120
rect 562498 -1176 562566 -1120
rect 562622 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect -1916 -1244 597980 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 9234 -1244
rect 9290 -1300 9358 -1244
rect 9414 -1300 9482 -1244
rect 9538 -1300 9606 -1244
rect 9662 -1300 39954 -1244
rect 40010 -1300 40078 -1244
rect 40134 -1300 40202 -1244
rect 40258 -1300 40326 -1244
rect 40382 -1300 70674 -1244
rect 70730 -1300 70798 -1244
rect 70854 -1300 70922 -1244
rect 70978 -1300 71046 -1244
rect 71102 -1300 101394 -1244
rect 101450 -1300 101518 -1244
rect 101574 -1300 101642 -1244
rect 101698 -1300 101766 -1244
rect 101822 -1300 132114 -1244
rect 132170 -1300 132238 -1244
rect 132294 -1300 132362 -1244
rect 132418 -1300 132486 -1244
rect 132542 -1300 162834 -1244
rect 162890 -1300 162958 -1244
rect 163014 -1300 163082 -1244
rect 163138 -1300 163206 -1244
rect 163262 -1300 193554 -1244
rect 193610 -1300 193678 -1244
rect 193734 -1300 193802 -1244
rect 193858 -1300 193926 -1244
rect 193982 -1300 224274 -1244
rect 224330 -1300 224398 -1244
rect 224454 -1300 224522 -1244
rect 224578 -1300 224646 -1244
rect 224702 -1300 254994 -1244
rect 255050 -1300 255118 -1244
rect 255174 -1300 255242 -1244
rect 255298 -1300 255366 -1244
rect 255422 -1300 285714 -1244
rect 285770 -1300 285838 -1244
rect 285894 -1300 285962 -1244
rect 286018 -1300 286086 -1244
rect 286142 -1300 316434 -1244
rect 316490 -1300 316558 -1244
rect 316614 -1300 316682 -1244
rect 316738 -1300 316806 -1244
rect 316862 -1300 347154 -1244
rect 347210 -1300 347278 -1244
rect 347334 -1300 347402 -1244
rect 347458 -1300 347526 -1244
rect 347582 -1300 377874 -1244
rect 377930 -1300 377998 -1244
rect 378054 -1300 378122 -1244
rect 378178 -1300 378246 -1244
rect 378302 -1300 408594 -1244
rect 408650 -1300 408718 -1244
rect 408774 -1300 408842 -1244
rect 408898 -1300 408966 -1244
rect 409022 -1300 439314 -1244
rect 439370 -1300 439438 -1244
rect 439494 -1300 439562 -1244
rect 439618 -1300 439686 -1244
rect 439742 -1300 470034 -1244
rect 470090 -1300 470158 -1244
rect 470214 -1300 470282 -1244
rect 470338 -1300 470406 -1244
rect 470462 -1300 500754 -1244
rect 500810 -1300 500878 -1244
rect 500934 -1300 501002 -1244
rect 501058 -1300 501126 -1244
rect 501182 -1300 531474 -1244
rect 531530 -1300 531598 -1244
rect 531654 -1300 531722 -1244
rect 531778 -1300 531846 -1244
rect 531902 -1300 562194 -1244
rect 562250 -1300 562318 -1244
rect 562374 -1300 562442 -1244
rect 562498 -1300 562566 -1244
rect 562622 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect -1916 -1368 597980 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 9234 -1368
rect 9290 -1424 9358 -1368
rect 9414 -1424 9482 -1368
rect 9538 -1424 9606 -1368
rect 9662 -1424 39954 -1368
rect 40010 -1424 40078 -1368
rect 40134 -1424 40202 -1368
rect 40258 -1424 40326 -1368
rect 40382 -1424 70674 -1368
rect 70730 -1424 70798 -1368
rect 70854 -1424 70922 -1368
rect 70978 -1424 71046 -1368
rect 71102 -1424 101394 -1368
rect 101450 -1424 101518 -1368
rect 101574 -1424 101642 -1368
rect 101698 -1424 101766 -1368
rect 101822 -1424 132114 -1368
rect 132170 -1424 132238 -1368
rect 132294 -1424 132362 -1368
rect 132418 -1424 132486 -1368
rect 132542 -1424 162834 -1368
rect 162890 -1424 162958 -1368
rect 163014 -1424 163082 -1368
rect 163138 -1424 163206 -1368
rect 163262 -1424 193554 -1368
rect 193610 -1424 193678 -1368
rect 193734 -1424 193802 -1368
rect 193858 -1424 193926 -1368
rect 193982 -1424 224274 -1368
rect 224330 -1424 224398 -1368
rect 224454 -1424 224522 -1368
rect 224578 -1424 224646 -1368
rect 224702 -1424 254994 -1368
rect 255050 -1424 255118 -1368
rect 255174 -1424 255242 -1368
rect 255298 -1424 255366 -1368
rect 255422 -1424 285714 -1368
rect 285770 -1424 285838 -1368
rect 285894 -1424 285962 -1368
rect 286018 -1424 286086 -1368
rect 286142 -1424 316434 -1368
rect 316490 -1424 316558 -1368
rect 316614 -1424 316682 -1368
rect 316738 -1424 316806 -1368
rect 316862 -1424 347154 -1368
rect 347210 -1424 347278 -1368
rect 347334 -1424 347402 -1368
rect 347458 -1424 347526 -1368
rect 347582 -1424 377874 -1368
rect 377930 -1424 377998 -1368
rect 378054 -1424 378122 -1368
rect 378178 -1424 378246 -1368
rect 378302 -1424 408594 -1368
rect 408650 -1424 408718 -1368
rect 408774 -1424 408842 -1368
rect 408898 -1424 408966 -1368
rect 409022 -1424 439314 -1368
rect 439370 -1424 439438 -1368
rect 439494 -1424 439562 -1368
rect 439618 -1424 439686 -1368
rect 439742 -1424 470034 -1368
rect 470090 -1424 470158 -1368
rect 470214 -1424 470282 -1368
rect 470338 -1424 470406 -1368
rect 470462 -1424 500754 -1368
rect 500810 -1424 500878 -1368
rect 500934 -1424 501002 -1368
rect 501058 -1424 501126 -1368
rect 501182 -1424 531474 -1368
rect 531530 -1424 531598 -1368
rect 531654 -1424 531722 -1368
rect 531778 -1424 531846 -1368
rect 531902 -1424 562194 -1368
rect 562250 -1424 562318 -1368
rect 562374 -1424 562442 -1368
rect 562498 -1424 562566 -1368
rect 562622 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect -1916 -1492 597980 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 9234 -1492
rect 9290 -1548 9358 -1492
rect 9414 -1548 9482 -1492
rect 9538 -1548 9606 -1492
rect 9662 -1548 39954 -1492
rect 40010 -1548 40078 -1492
rect 40134 -1548 40202 -1492
rect 40258 -1548 40326 -1492
rect 40382 -1548 70674 -1492
rect 70730 -1548 70798 -1492
rect 70854 -1548 70922 -1492
rect 70978 -1548 71046 -1492
rect 71102 -1548 101394 -1492
rect 101450 -1548 101518 -1492
rect 101574 -1548 101642 -1492
rect 101698 -1548 101766 -1492
rect 101822 -1548 132114 -1492
rect 132170 -1548 132238 -1492
rect 132294 -1548 132362 -1492
rect 132418 -1548 132486 -1492
rect 132542 -1548 162834 -1492
rect 162890 -1548 162958 -1492
rect 163014 -1548 163082 -1492
rect 163138 -1548 163206 -1492
rect 163262 -1548 193554 -1492
rect 193610 -1548 193678 -1492
rect 193734 -1548 193802 -1492
rect 193858 -1548 193926 -1492
rect 193982 -1548 224274 -1492
rect 224330 -1548 224398 -1492
rect 224454 -1548 224522 -1492
rect 224578 -1548 224646 -1492
rect 224702 -1548 254994 -1492
rect 255050 -1548 255118 -1492
rect 255174 -1548 255242 -1492
rect 255298 -1548 255366 -1492
rect 255422 -1548 285714 -1492
rect 285770 -1548 285838 -1492
rect 285894 -1548 285962 -1492
rect 286018 -1548 286086 -1492
rect 286142 -1548 316434 -1492
rect 316490 -1548 316558 -1492
rect 316614 -1548 316682 -1492
rect 316738 -1548 316806 -1492
rect 316862 -1548 347154 -1492
rect 347210 -1548 347278 -1492
rect 347334 -1548 347402 -1492
rect 347458 -1548 347526 -1492
rect 347582 -1548 377874 -1492
rect 377930 -1548 377998 -1492
rect 378054 -1548 378122 -1492
rect 378178 -1548 378246 -1492
rect 378302 -1548 408594 -1492
rect 408650 -1548 408718 -1492
rect 408774 -1548 408842 -1492
rect 408898 -1548 408966 -1492
rect 409022 -1548 439314 -1492
rect 439370 -1548 439438 -1492
rect 439494 -1548 439562 -1492
rect 439618 -1548 439686 -1492
rect 439742 -1548 470034 -1492
rect 470090 -1548 470158 -1492
rect 470214 -1548 470282 -1492
rect 470338 -1548 470406 -1492
rect 470462 -1548 500754 -1492
rect 500810 -1548 500878 -1492
rect 500934 -1548 501002 -1492
rect 501058 -1548 501126 -1492
rect 501182 -1548 531474 -1492
rect 531530 -1548 531598 -1492
rect 531654 -1548 531722 -1492
rect 531778 -1548 531846 -1492
rect 531902 -1548 562194 -1492
rect 562250 -1548 562318 -1492
rect 562374 -1548 562442 -1492
rect 562498 -1548 562566 -1492
rect 562622 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect -1916 -1644 597980 -1548
use avali_logo  avali_logo
timestamp 0
transform 1 0 60000 0 1 480000
box 0 0 75000 88050
use wrapped_ay8913  ay8913
timestamp 0
transform 1 0 40000 0 1 240000
box 1258 0 60000 60000
use blinker  blinker
timestamp 0
transform 1 0 290000 0 1 50000
box 1258 0 34768 32230
use hellorld  hellorld
timestamp 0
transform 1 0 160000 0 1 260000
box 1258 1792 26000 26000
use wrapped_mc14500  mc14500
timestamp 0
transform 1 0 480000 0 1 200000
box 1258 0 37000 37000
use multiplexer  multiplexer
timestamp 0
transform 1 0 236000 0 1 256000
box 0 0 140000 130000
use wrapped_sid  sid
timestamp 0
transform 1 0 40000 0 1 50000
box 1258 0 230000 160000
use tholin_avalonsemi_tbb1143  tbb1143
timestamp 0
transform 1 0 150000 0 1 320000
box 1258 2688 46000 43120
use wrapped_pdp11  wrapped_pdp11
timestamp 0
transform 1 0 190000 0 1 410000
box 0 0 360000 158686
use wrapped_qcpu  wrapped_qcpu
timestamp 0
transform 1 0 460000 0 1 50000
box 0 802 100000 100000
use wrapped_sn76489  wrapped_sn76489
timestamp 0
transform 1 0 360000 0 1 50000
box 0 3076 60000 70000
<< labels >>
flabel metal3 s 595560 7112 597000 7336 0 FreeSans 896 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 595560 403592 597000 403816 0 FreeSans 896 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 595560 443240 597000 443464 0 FreeSans 896 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 595560 482888 597000 483112 0 FreeSans 896 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 595560 522536 597000 522760 0 FreeSans 896 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 595560 562184 597000 562408 0 FreeSans 896 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 584696 595560 584920 597000 0 FreeSans 896 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 518504 595560 518728 597000 0 FreeSans 896 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 452312 595560 452536 597000 0 FreeSans 896 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 386120 595560 386344 597000 0 FreeSans 896 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 319928 595560 320152 597000 0 FreeSans 896 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 595560 46760 597000 46984 0 FreeSans 896 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 253736 595560 253960 597000 0 FreeSans 896 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 187544 595560 187768 597000 0 FreeSans 896 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 121352 595560 121576 597000 0 FreeSans 896 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 55160 595560 55384 597000 0 FreeSans 896 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -960 587160 480 587384 0 FreeSans 896 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -960 544824 480 545048 0 FreeSans 896 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -960 502488 480 502712 0 FreeSans 896 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -960 460152 480 460376 0 FreeSans 896 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -960 417816 480 418040 0 FreeSans 896 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -960 375480 480 375704 0 FreeSans 896 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 595560 86408 597000 86632 0 FreeSans 896 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -960 333144 480 333368 0 FreeSans 896 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -960 290808 480 291032 0 FreeSans 896 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -960 248472 480 248696 0 FreeSans 896 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -960 206136 480 206360 0 FreeSans 896 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -960 163800 480 164024 0 FreeSans 896 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -960 121464 480 121688 0 FreeSans 896 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -960 79128 480 79352 0 FreeSans 896 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -960 36792 480 37016 0 FreeSans 896 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 595560 126056 597000 126280 0 FreeSans 896 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 595560 165704 597000 165928 0 FreeSans 896 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 595560 205352 597000 205576 0 FreeSans 896 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 595560 245000 597000 245224 0 FreeSans 896 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 595560 284648 597000 284872 0 FreeSans 896 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 595560 324296 597000 324520 0 FreeSans 896 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 595560 363944 597000 364168 0 FreeSans 896 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 595560 33544 597000 33768 0 FreeSans 896 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 595560 430024 597000 430248 0 FreeSans 896 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 595560 469672 597000 469896 0 FreeSans 896 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 595560 509320 597000 509544 0 FreeSans 896 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 595560 548968 597000 549192 0 FreeSans 896 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 595560 588616 597000 588840 0 FreeSans 896 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 540568 595560 540792 597000 0 FreeSans 896 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 474376 595560 474600 597000 0 FreeSans 896 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 408184 595560 408408 597000 0 FreeSans 896 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 341992 595560 342216 597000 0 FreeSans 896 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 275800 595560 276024 597000 0 FreeSans 896 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 595560 73192 597000 73416 0 FreeSans 896 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 209608 595560 209832 597000 0 FreeSans 896 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 143416 595560 143640 597000 0 FreeSans 896 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 77224 595560 77448 597000 0 FreeSans 896 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 11032 595560 11256 597000 0 FreeSans 896 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -960 558936 480 559160 0 FreeSans 896 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -960 516600 480 516824 0 FreeSans 896 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -960 474264 480 474488 0 FreeSans 896 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -960 431928 480 432152 0 FreeSans 896 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -960 389592 480 389816 0 FreeSans 896 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -960 347256 480 347480 0 FreeSans 896 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 595560 112840 597000 113064 0 FreeSans 896 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -960 304920 480 305144 0 FreeSans 896 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -960 262584 480 262808 0 FreeSans 896 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -960 220248 480 220472 0 FreeSans 896 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -960 177912 480 178136 0 FreeSans 896 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -960 135576 480 135800 0 FreeSans 896 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -960 93240 480 93464 0 FreeSans 896 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -960 50904 480 51128 0 FreeSans 896 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -960 8568 480 8792 0 FreeSans 896 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 595560 152488 597000 152712 0 FreeSans 896 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 595560 192136 597000 192360 0 FreeSans 896 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 595560 231784 597000 232008 0 FreeSans 896 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 595560 271432 597000 271656 0 FreeSans 896 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 595560 311080 597000 311304 0 FreeSans 896 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 595560 350728 597000 350952 0 FreeSans 896 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 595560 390376 597000 390600 0 FreeSans 896 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 595560 20328 597000 20552 0 FreeSans 896 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 595560 416808 597000 417032 0 FreeSans 896 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 595560 456456 597000 456680 0 FreeSans 896 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 595560 496104 597000 496328 0 FreeSans 896 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 595560 535752 597000 535976 0 FreeSans 896 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 595560 575400 597000 575624 0 FreeSans 896 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 562632 595560 562856 597000 0 FreeSans 896 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 496440 595560 496664 597000 0 FreeSans 896 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 430248 595560 430472 597000 0 FreeSans 896 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 364056 595560 364280 597000 0 FreeSans 896 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 297864 595560 298088 597000 0 FreeSans 896 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 595560 59976 597000 60200 0 FreeSans 896 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 231672 595560 231896 597000 0 FreeSans 896 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 165480 595560 165704 597000 0 FreeSans 896 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 99288 595560 99512 597000 0 FreeSans 896 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 33096 595560 33320 597000 0 FreeSans 896 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -960 573048 480 573272 0 FreeSans 896 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -960 530712 480 530936 0 FreeSans 896 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -960 488376 480 488600 0 FreeSans 896 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -960 446040 480 446264 0 FreeSans 896 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -960 403704 480 403928 0 FreeSans 896 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -960 361368 480 361592 0 FreeSans 896 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 595560 99624 597000 99848 0 FreeSans 896 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -960 319032 480 319256 0 FreeSans 896 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -960 276696 480 276920 0 FreeSans 896 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -960 234360 480 234584 0 FreeSans 896 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -960 192024 480 192248 0 FreeSans 896 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -960 149688 480 149912 0 FreeSans 896 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -960 107352 480 107576 0 FreeSans 896 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -960 65016 480 65240 0 FreeSans 896 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -960 22680 480 22904 0 FreeSans 896 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 595560 139272 597000 139496 0 FreeSans 896 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 595560 178920 597000 179144 0 FreeSans 896 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 595560 218568 597000 218792 0 FreeSans 896 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 595560 258216 597000 258440 0 FreeSans 896 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 595560 297864 597000 298088 0 FreeSans 896 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 595560 337512 597000 337736 0 FreeSans 896 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 595560 377160 597000 377384 0 FreeSans 896 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 213192 -960 213416 480 0 FreeSans 896 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 270312 -960 270536 480 0 FreeSans 896 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 276024 -960 276248 480 0 FreeSans 896 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 281736 -960 281960 480 0 FreeSans 896 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 287448 -960 287672 480 0 FreeSans 896 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 293160 -960 293384 480 0 FreeSans 896 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 298872 -960 299096 480 0 FreeSans 896 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 304584 -960 304808 480 0 FreeSans 896 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 310296 -960 310520 480 0 FreeSans 896 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 316008 -960 316232 480 0 FreeSans 896 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 321720 -960 321944 480 0 FreeSans 896 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 218904 -960 219128 480 0 FreeSans 896 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 327432 -960 327656 480 0 FreeSans 896 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 333144 -960 333368 480 0 FreeSans 896 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 338856 -960 339080 480 0 FreeSans 896 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 344568 -960 344792 480 0 FreeSans 896 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 350280 -960 350504 480 0 FreeSans 896 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 355992 -960 356216 480 0 FreeSans 896 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 361704 -960 361928 480 0 FreeSans 896 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 367416 -960 367640 480 0 FreeSans 896 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 373128 -960 373352 480 0 FreeSans 896 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 378840 -960 379064 480 0 FreeSans 896 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 224616 -960 224840 480 0 FreeSans 896 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 384552 -960 384776 480 0 FreeSans 896 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 390264 -960 390488 480 0 FreeSans 896 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 395976 -960 396200 480 0 FreeSans 896 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 401688 -960 401912 480 0 FreeSans 896 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 407400 -960 407624 480 0 FreeSans 896 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 413112 -960 413336 480 0 FreeSans 896 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 418824 -960 419048 480 0 FreeSans 896 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 424536 -960 424760 480 0 FreeSans 896 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 430248 -960 430472 480 0 FreeSans 896 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 435960 -960 436184 480 0 FreeSans 896 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 230328 -960 230552 480 0 FreeSans 896 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 441672 -960 441896 480 0 FreeSans 896 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 447384 -960 447608 480 0 FreeSans 896 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 453096 -960 453320 480 0 FreeSans 896 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 458808 -960 459032 480 0 FreeSans 896 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 464520 -960 464744 480 0 FreeSans 896 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 470232 -960 470456 480 0 FreeSans 896 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 475944 -960 476168 480 0 FreeSans 896 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 481656 -960 481880 480 0 FreeSans 896 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 487368 -960 487592 480 0 FreeSans 896 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 493080 -960 493304 480 0 FreeSans 896 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 236040 -960 236264 480 0 FreeSans 896 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 498792 -960 499016 480 0 FreeSans 896 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 504504 -960 504728 480 0 FreeSans 896 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 510216 -960 510440 480 0 FreeSans 896 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 515928 -960 516152 480 0 FreeSans 896 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 521640 -960 521864 480 0 FreeSans 896 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 527352 -960 527576 480 0 FreeSans 896 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 533064 -960 533288 480 0 FreeSans 896 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 538776 -960 539000 480 0 FreeSans 896 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 544488 -960 544712 480 0 FreeSans 896 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 550200 -960 550424 480 0 FreeSans 896 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 241752 -960 241976 480 0 FreeSans 896 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 555912 -960 556136 480 0 FreeSans 896 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 561624 -960 561848 480 0 FreeSans 896 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 567336 -960 567560 480 0 FreeSans 896 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 573048 -960 573272 480 0 FreeSans 896 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 247464 -960 247688 480 0 FreeSans 896 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 253176 -960 253400 480 0 FreeSans 896 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 258888 -960 259112 480 0 FreeSans 896 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 264600 -960 264824 480 0 FreeSans 896 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 215096 -960 215320 480 0 FreeSans 896 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal2 s 272216 -960 272440 480 0 FreeSans 896 90 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal2 s 277928 -960 278152 480 0 FreeSans 896 90 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal2 s 283640 -960 283864 480 0 FreeSans 896 90 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 289352 -960 289576 480 0 FreeSans 896 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal2 s 295064 -960 295288 480 0 FreeSans 896 90 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal2 s 300776 -960 301000 480 0 FreeSans 896 90 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal2 s 306488 -960 306712 480 0 FreeSans 896 90 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 312200 -960 312424 480 0 FreeSans 896 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal2 s 317912 -960 318136 480 0 FreeSans 896 90 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 323624 -960 323848 480 0 FreeSans 896 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal2 s 220808 -960 221032 480 0 FreeSans 896 90 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal2 s 329336 -960 329560 480 0 FreeSans 896 90 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal2 s 335048 -960 335272 480 0 FreeSans 896 90 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal2 s 340760 -960 340984 480 0 FreeSans 896 90 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 346472 -960 346696 480 0 FreeSans 896 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal2 s 352184 -960 352408 480 0 FreeSans 896 90 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 357896 -960 358120 480 0 FreeSans 896 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal2 s 363608 -960 363832 480 0 FreeSans 896 90 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 369320 -960 369544 480 0 FreeSans 896 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal2 s 375032 -960 375256 480 0 FreeSans 896 90 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 380744 -960 380968 480 0 FreeSans 896 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal2 s 226520 -960 226744 480 0 FreeSans 896 90 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal2 s 386456 -960 386680 480 0 FreeSans 896 90 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal2 s 392168 -960 392392 480 0 FreeSans 896 90 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 397880 -960 398104 480 0 FreeSans 896 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal2 s 403592 -960 403816 480 0 FreeSans 896 90 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 409304 -960 409528 480 0 FreeSans 896 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 415016 -960 415240 480 0 FreeSans 896 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal2 s 420728 -960 420952 480 0 FreeSans 896 90 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal2 s 426440 -960 426664 480 0 FreeSans 896 90 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal2 s 432152 -960 432376 480 0 FreeSans 896 90 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal2 s 437864 -960 438088 480 0 FreeSans 896 90 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal2 s 232232 -960 232456 480 0 FreeSans 896 90 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal2 s 443576 -960 443800 480 0 FreeSans 896 90 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal2 s 449288 -960 449512 480 0 FreeSans 896 90 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal2 s 455000 -960 455224 480 0 FreeSans 896 90 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 460712 -960 460936 480 0 FreeSans 896 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 466424 -960 466648 480 0 FreeSans 896 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 472136 -960 472360 480 0 FreeSans 896 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 477848 -960 478072 480 0 FreeSans 896 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal2 s 483560 -960 483784 480 0 FreeSans 896 90 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 489272 -960 489496 480 0 FreeSans 896 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 494984 -960 495208 480 0 FreeSans 896 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 237944 -960 238168 480 0 FreeSans 896 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 500696 -960 500920 480 0 FreeSans 896 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal2 s 506408 -960 506632 480 0 FreeSans 896 90 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal2 s 512120 -960 512344 480 0 FreeSans 896 90 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal2 s 517832 -960 518056 480 0 FreeSans 896 90 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal2 s 523544 -960 523768 480 0 FreeSans 896 90 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 529256 -960 529480 480 0 FreeSans 896 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal2 s 534968 -960 535192 480 0 FreeSans 896 90 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 540680 -960 540904 480 0 FreeSans 896 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal2 s 546392 -960 546616 480 0 FreeSans 896 90 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal2 s 552104 -960 552328 480 0 FreeSans 896 90 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal2 s 243656 -960 243880 480 0 FreeSans 896 90 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 557816 -960 558040 480 0 FreeSans 896 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 563528 -960 563752 480 0 FreeSans 896 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 569240 -960 569464 480 0 FreeSans 896 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal2 s 574952 -960 575176 480 0 FreeSans 896 90 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal2 s 249368 -960 249592 480 0 FreeSans 896 90 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 255080 -960 255304 480 0 FreeSans 896 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal2 s 260792 -960 261016 480 0 FreeSans 896 90 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal2 s 266504 -960 266728 480 0 FreeSans 896 90 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal2 s 217000 -960 217224 480 0 FreeSans 896 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 274120 -960 274344 480 0 FreeSans 896 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 279832 -960 280056 480 0 FreeSans 896 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 285544 -960 285768 480 0 FreeSans 896 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 291256 -960 291480 480 0 FreeSans 896 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 296968 -960 297192 480 0 FreeSans 896 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 302680 -960 302904 480 0 FreeSans 896 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 308392 -960 308616 480 0 FreeSans 896 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 314104 -960 314328 480 0 FreeSans 896 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 319816 -960 320040 480 0 FreeSans 896 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 325528 -960 325752 480 0 FreeSans 896 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 222712 -960 222936 480 0 FreeSans 896 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 331240 -960 331464 480 0 FreeSans 896 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 336952 -960 337176 480 0 FreeSans 896 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 342664 -960 342888 480 0 FreeSans 896 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 348376 -960 348600 480 0 FreeSans 896 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 354088 -960 354312 480 0 FreeSans 896 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 359800 -960 360024 480 0 FreeSans 896 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 365512 -960 365736 480 0 FreeSans 896 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 371224 -960 371448 480 0 FreeSans 896 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 376936 -960 377160 480 0 FreeSans 896 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 382648 -960 382872 480 0 FreeSans 896 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 228424 -960 228648 480 0 FreeSans 896 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 388360 -960 388584 480 0 FreeSans 896 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 394072 -960 394296 480 0 FreeSans 896 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 399784 -960 400008 480 0 FreeSans 896 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 405496 -960 405720 480 0 FreeSans 896 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 411208 -960 411432 480 0 FreeSans 896 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 416920 -960 417144 480 0 FreeSans 896 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 422632 -960 422856 480 0 FreeSans 896 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 428344 -960 428568 480 0 FreeSans 896 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 434056 -960 434280 480 0 FreeSans 896 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 439768 -960 439992 480 0 FreeSans 896 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 234136 -960 234360 480 0 FreeSans 896 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 445480 -960 445704 480 0 FreeSans 896 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 451192 -960 451416 480 0 FreeSans 896 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 456904 -960 457128 480 0 FreeSans 896 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 462616 -960 462840 480 0 FreeSans 896 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 468328 -960 468552 480 0 FreeSans 896 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 474040 -960 474264 480 0 FreeSans 896 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 479752 -960 479976 480 0 FreeSans 896 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 485464 -960 485688 480 0 FreeSans 896 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 491176 -960 491400 480 0 FreeSans 896 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 496888 -960 497112 480 0 FreeSans 896 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 239848 -960 240072 480 0 FreeSans 896 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 502600 -960 502824 480 0 FreeSans 896 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 508312 -960 508536 480 0 FreeSans 896 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 514024 -960 514248 480 0 FreeSans 896 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 519736 -960 519960 480 0 FreeSans 896 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 525448 -960 525672 480 0 FreeSans 896 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 531160 -960 531384 480 0 FreeSans 896 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 536872 -960 537096 480 0 FreeSans 896 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 542584 -960 542808 480 0 FreeSans 896 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 548296 -960 548520 480 0 FreeSans 896 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 554008 -960 554232 480 0 FreeSans 896 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 245560 -960 245784 480 0 FreeSans 896 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 559720 -960 559944 480 0 FreeSans 896 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 565432 -960 565656 480 0 FreeSans 896 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 571144 -960 571368 480 0 FreeSans 896 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 576856 -960 577080 480 0 FreeSans 896 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 251272 -960 251496 480 0 FreeSans 896 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 256984 -960 257208 480 0 FreeSans 896 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 262696 -960 262920 480 0 FreeSans 896 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 268408 -960 268632 480 0 FreeSans 896 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 578760 -960 578984 480 0 FreeSans 896 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 580664 -960 580888 480 0 FreeSans 896 90 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 582568 -960 582792 480 0 FreeSans 896 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal2 s 584472 -960 584696 480 0 FreeSans 896 90 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s -956 -684 -336 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 -684 597020 -64 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 596688 597020 597308 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 596400 -684 597020 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 5418 -1644 6038 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 36138 -1644 36758 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 -1644 67478 48802 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 210462 67478 245074 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 298094 67478 488238 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 532362 67478 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 -1644 98198 48802 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 210462 98198 478338 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 542112 98198 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128298 -1644 128918 48802 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128298 210462 128918 497538 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128298 543612 128918 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 -1644 159638 48802 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 210462 159638 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 -1644 190358 48802 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 210462 190358 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 -1644 221078 48802 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 210462 221078 408578 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 569342 221078 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 -1644 251798 48802 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 210462 251798 257490 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 569342 251798 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 -1644 282518 257490 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 569342 282518 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 -1644 313238 257490 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 569342 313238 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 -1644 343958 257490 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 569342 343958 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 -1644 374678 53730 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 115262 374678 257490 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 569342 374678 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 -1644 405398 53730 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 115262 405398 408578 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 569342 405398 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 -1644 436118 408578 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 569342 436118 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 466218 -1644 466838 48690 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 466218 149870 466838 408578 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 466218 569342 466838 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 -1644 497558 48690 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 149870 497558 203170 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 233230 497558 408578 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 569342 497558 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 527658 -1644 528278 48690 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 527658 149870 528278 408578 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 527658 569342 528278 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 558378 -1644 558998 48690 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 558378 149870 558998 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 589098 -1644 589718 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 3826 597980 4446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 21826 597980 22446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 39826 597980 40446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 57826 597980 58446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 75826 597980 76446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 93826 597980 94446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 111826 597980 112446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 129826 597980 130446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 147826 597980 148446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 165826 597980 166446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 183826 597980 184446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 201826 597980 202446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 219826 597980 220446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 237826 597980 238446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 255826 597980 256446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 273826 597980 274446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 291826 597980 292446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 309826 597980 310446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 327826 597980 328446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 345826 597980 346446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 363826 597980 364446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 381826 597980 382446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 399826 597980 400446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 417826 597980 418446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 435826 597980 436446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 453826 597980 454446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 471826 597980 472446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 489826 597980 490446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 507826 597980 508446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 525826 597980 526446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 543826 597980 544446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 561826 597980 562446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 579826 597980 580446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -1916 -1644 -1296 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 -1644 597980 -1024 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 597648 597980 598268 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 597360 -1644 597980 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 9138 -1644 9758 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 39858 -1644 40478 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 -1644 71198 48802 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 210462 71198 245074 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 298094 71198 484638 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 535962 71198 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 -1644 101918 48802 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 210462 101918 479238 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 547962 101918 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 -1644 132638 48802 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 210462 132638 500388 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 544962 132638 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 -1644 163358 48802 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 210462 163358 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 -1644 194078 48802 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 210462 194078 408578 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 569342 194078 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 -1644 224798 48802 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 210462 224798 408578 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 569342 224798 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 -1644 255518 48802 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 210462 255518 257490 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 383870 255518 408578 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 569342 255518 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 -1644 286238 257490 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 383870 286238 408578 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 569342 286238 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 -1644 316958 50964 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 84316 316958 257490 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 383870 316958 408578 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 569342 316958 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 -1644 347678 257490 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 383870 347678 408578 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 569342 347678 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 -1644 378398 53730 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 115262 378398 408578 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 569342 378398 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 -1644 409118 53730 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 115262 409118 408578 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 569342 409118 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 439218 -1644 439838 408578 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 439218 569342 439838 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 469938 -1644 470558 48690 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 469938 149870 470558 408578 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 469938 569342 470558 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 -1644 501278 48690 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 149870 501278 203170 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 233230 501278 408578 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 569342 501278 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 531378 -1644 531998 48690 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 531378 149870 531998 408578 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 531378 569342 531998 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 562098 -1644 562718 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 592818 -1644 593438 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 9826 597980 10446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 27826 597980 28446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 45826 597980 46446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 63826 597980 64446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 81826 597980 82446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 99826 597980 100446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 117826 597980 118446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 135826 597980 136446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 153826 597980 154446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 171826 597980 172446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 189826 597980 190446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 207826 597980 208446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 225826 597980 226446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 243826 597980 244446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 261826 597980 262446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 279826 597980 280446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 297826 597980 298446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 315826 597980 316446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 333826 597980 334446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 351826 597980 352446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 369826 597980 370446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 387826 597980 388446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 405826 597980 406446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 423826 597980 424446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 441826 597980 442446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 459826 597980 460446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 477826 597980 478446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 495826 597980 496446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 513826 597980 514446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 531826 597980 532446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 549826 597980 550446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 567826 597980 568446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 585826 597980 586446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 11368 -960 11592 480 0 FreeSans 896 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 13272 -960 13496 480 0 FreeSans 896 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 15176 -960 15400 480 0 FreeSans 896 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 22792 -960 23016 480 0 FreeSans 896 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 87528 -960 87752 480 0 FreeSans 896 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 93240 -960 93464 480 0 FreeSans 896 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 98952 -960 99176 480 0 FreeSans 896 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 104664 -960 104888 480 0 FreeSans 896 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 110376 -960 110600 480 0 FreeSans 896 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 116088 -960 116312 480 0 FreeSans 896 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 121800 -960 122024 480 0 FreeSans 896 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 127512 -960 127736 480 0 FreeSans 896 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 133224 -960 133448 480 0 FreeSans 896 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 138936 -960 139160 480 0 FreeSans 896 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 30408 -960 30632 480 0 FreeSans 896 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 144648 -960 144872 480 0 FreeSans 896 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 150360 -960 150584 480 0 FreeSans 896 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 156072 -960 156296 480 0 FreeSans 896 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 161784 -960 162008 480 0 FreeSans 896 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 167496 -960 167720 480 0 FreeSans 896 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 173208 -960 173432 480 0 FreeSans 896 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 178920 -960 179144 480 0 FreeSans 896 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 184632 -960 184856 480 0 FreeSans 896 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 190344 -960 190568 480 0 FreeSans 896 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 196056 -960 196280 480 0 FreeSans 896 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 38024 -960 38248 480 0 FreeSans 896 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 201768 -960 201992 480 0 FreeSans 896 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 207480 -960 207704 480 0 FreeSans 896 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 45640 -960 45864 480 0 FreeSans 896 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 53256 -960 53480 480 0 FreeSans 896 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 58968 -960 59192 480 0 FreeSans 896 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 64680 -960 64904 480 0 FreeSans 896 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 70392 -960 70616 480 0 FreeSans 896 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 76104 -960 76328 480 0 FreeSans 896 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 81816 -960 82040 480 0 FreeSans 896 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 17080 -960 17304 480 0 FreeSans 896 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 24696 -960 24920 480 0 FreeSans 896 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 89432 -960 89656 480 0 FreeSans 896 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 95144 -960 95368 480 0 FreeSans 896 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 100856 -960 101080 480 0 FreeSans 896 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 106568 -960 106792 480 0 FreeSans 896 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 112280 -960 112504 480 0 FreeSans 896 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 117992 -960 118216 480 0 FreeSans 896 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 123704 -960 123928 480 0 FreeSans 896 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 129416 -960 129640 480 0 FreeSans 896 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 135128 -960 135352 480 0 FreeSans 896 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 140840 -960 141064 480 0 FreeSans 896 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 32312 -960 32536 480 0 FreeSans 896 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 146552 -960 146776 480 0 FreeSans 896 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 152264 -960 152488 480 0 FreeSans 896 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 157976 -960 158200 480 0 FreeSans 896 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 163688 -960 163912 480 0 FreeSans 896 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 169400 -960 169624 480 0 FreeSans 896 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 175112 -960 175336 480 0 FreeSans 896 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 180824 -960 181048 480 0 FreeSans 896 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 186536 -960 186760 480 0 FreeSans 896 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 192248 -960 192472 480 0 FreeSans 896 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 197960 -960 198184 480 0 FreeSans 896 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 39928 -960 40152 480 0 FreeSans 896 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 203672 -960 203896 480 0 FreeSans 896 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 209384 -960 209608 480 0 FreeSans 896 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 47544 -960 47768 480 0 FreeSans 896 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 55160 -960 55384 480 0 FreeSans 896 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 60872 -960 61096 480 0 FreeSans 896 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 66584 -960 66808 480 0 FreeSans 896 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 72296 -960 72520 480 0 FreeSans 896 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 78008 -960 78232 480 0 FreeSans 896 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 83720 -960 83944 480 0 FreeSans 896 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 26600 -960 26824 480 0 FreeSans 896 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 91336 -960 91560 480 0 FreeSans 896 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 97048 -960 97272 480 0 FreeSans 896 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 102760 -960 102984 480 0 FreeSans 896 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 108472 -960 108696 480 0 FreeSans 896 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 114184 -960 114408 480 0 FreeSans 896 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 119896 -960 120120 480 0 FreeSans 896 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 125608 -960 125832 480 0 FreeSans 896 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 131320 -960 131544 480 0 FreeSans 896 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 137032 -960 137256 480 0 FreeSans 896 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 142744 -960 142968 480 0 FreeSans 896 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 34216 -960 34440 480 0 FreeSans 896 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 148456 -960 148680 480 0 FreeSans 896 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 154168 -960 154392 480 0 FreeSans 896 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 159880 -960 160104 480 0 FreeSans 896 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 165592 -960 165816 480 0 FreeSans 896 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 171304 -960 171528 480 0 FreeSans 896 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 177016 -960 177240 480 0 FreeSans 896 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 182728 -960 182952 480 0 FreeSans 896 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 188440 -960 188664 480 0 FreeSans 896 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 194152 -960 194376 480 0 FreeSans 896 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 199864 -960 200088 480 0 FreeSans 896 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 41832 -960 42056 480 0 FreeSans 896 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 205576 -960 205800 480 0 FreeSans 896 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 211288 -960 211512 480 0 FreeSans 896 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 49448 -960 49672 480 0 FreeSans 896 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 57064 -960 57288 480 0 FreeSans 896 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 62776 -960 63000 480 0 FreeSans 896 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 68488 -960 68712 480 0 FreeSans 896 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 74200 -960 74424 480 0 FreeSans 896 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 79912 -960 80136 480 0 FreeSans 896 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 85624 -960 85848 480 0 FreeSans 896 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 28504 -960 28728 480 0 FreeSans 896 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 36120 -960 36344 480 0 FreeSans 896 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 43736 -960 43960 480 0 FreeSans 896 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 51352 -960 51576 480 0 FreeSans 896 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 18984 -960 19208 480 0 FreeSans 896 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 20888 -960 21112 480 0 FreeSans 896 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel via4 395390 112322 395390 112322 0 vdd
rlabel via4 410750 100322 410750 100322 0 vss
rlabel metal2 42210 240520 42210 240520 0 ay8913_do\[0\]
rlabel metal2 219240 314720 219240 314720 0 ay8913_do\[10\]
rlabel metal2 116760 314496 116760 314496 0 ay8913_do\[11\]
rlabel metal2 234584 311472 234584 311472 0 ay8913_do\[12\]
rlabel metal2 68936 237594 68936 237594 0 ay8913_do\[13\]
rlabel metal2 70952 238322 70952 238322 0 ay8913_do\[14\]
rlabel metal2 72968 237538 72968 237538 0 ay8913_do\[15\]
rlabel metal4 74984 238007 74984 238007 0 ay8913_do\[16\]
rlabel metal4 77000 238097 77000 238097 0 ay8913_do\[17\]
rlabel metal2 217784 314216 217784 314216 0 ay8913_do\[18\]
rlabel metal4 309064 384832 309064 384832 0 ay8913_do\[19\]
rlabel metal2 44450 240520 44450 240520 0 ay8913_do\[1\]
rlabel metal2 100408 313824 100408 313824 0 ay8913_do\[20\]
rlabel metal2 120120 314888 120120 314888 0 ay8913_do\[21\]
rlabel metal2 311752 388038 311752 388038 0 ay8913_do\[22\]
rlabel metal4 95480 237944 95480 237944 0 ay8913_do\[23\]
rlabel metal2 91112 239274 91112 239274 0 ay8913_do\[24\]
rlabel metal3 100184 238560 100184 238560 0 ay8913_do\[25\]
rlabel metal3 100072 238336 100072 238336 0 ay8913_do\[26\]
rlabel metal2 97160 239106 97160 239106 0 ay8913_do\[27\]
rlabel metal2 46760 239274 46760 239274 0 ay8913_do\[2\]
rlabel metal2 48776 239162 48776 239162 0 ay8913_do\[3\]
rlabel metal3 88816 240744 88816 240744 0 ay8913_do\[4\]
rlabel metal2 210840 314384 210840 314384 0 ay8913_do\[5\]
rlabel metal4 212520 314705 212520 314705 0 ay8913_do\[6\]
rlabel metal3 56840 240016 56840 240016 0 ay8913_do\[7\]
rlabel metal2 215880 314608 215880 314608 0 ay8913_do\[8\]
rlabel metal2 217560 314552 217560 314552 0 ay8913_do\[9\]
rlabel metal2 307706 50232 307706 50232 0 blinker_do\[0\]
rlabel metal2 235704 298592 235704 298592 0 blinker_do\[1\]
rlabel metal2 235872 385560 235872 385560 0 blinker_do\[2\]
rlabel metal3 187558 261800 187558 261800 0 custom_settings\[0\]
rlabel metal3 185864 281666 185864 281666 0 custom_settings\[10\]
rlabel metal3 185864 284102 185864 284102 0 custom_settings\[11\]
rlabel metal3 188146 514920 188146 514920 0 custom_settings\[12\]
rlabel metal3 188874 522088 188874 522088 0 custom_settings\[13\]
rlabel metal3 188930 529256 188930 529256 0 custom_settings\[14\]
rlabel metal3 188202 536424 188202 536424 0 custom_settings\[15\]
rlabel metal3 188818 543592 188818 543592 0 custom_settings\[16\]
rlabel metal3 188258 550760 188258 550760 0 custom_settings\[17\]
rlabel metal3 188986 557928 188986 557928 0 custom_settings\[18\]
rlabel metal3 375928 320418 375928 320418 0 custom_settings\[19\]
rlabel metal3 185864 264222 185864 264222 0 custom_settings\[1\]
rlabel metal3 459368 115892 459368 115892 0 custom_settings\[20\]
rlabel metal3 457744 118888 457744 118888 0 custom_settings\[21\]
rlabel metal3 379918 324184 379918 324184 0 custom_settings\[22\]
rlabel metal3 459368 124684 459368 124684 0 custom_settings\[23\]
rlabel metal3 379078 326424 379078 326424 0 custom_settings\[24\]
rlabel metal4 451080 229040 451080 229040 0 custom_settings\[25\]
rlabel metal3 380758 328664 380758 328664 0 custom_settings\[26\]
rlabel metal3 381598 329784 381598 329784 0 custom_settings\[27\]
rlabel metal3 378238 330904 378238 330904 0 custom_settings\[28\]
rlabel metal3 382438 332024 382438 332024 0 custom_settings\[29\]
rlabel metal3 185864 266070 185864 266070 0 custom_settings\[2\]
rlabel metal3 383278 333144 383278 333144 0 custom_settings\[30\]
rlabel metal3 384958 334264 384958 334264 0 custom_settings\[31\]
rlabel metal4 235592 264870 235592 264870 0 custom_settings\[3\]
rlabel metal3 377622 304024 377622 304024 0 custom_settings\[4\]
rlabel metal3 377678 305144 377678 305144 0 custom_settings\[5\]
rlabel metal3 189042 471912 189042 471912 0 custom_settings\[6\]
rlabel metal3 377398 307384 377398 307384 0 custom_settings\[7\]
rlabel metal3 185864 277998 185864 277998 0 custom_settings\[8\]
rlabel metal3 187446 279944 187446 279944 0 custom_settings\[9\]
rlabel metal2 214200 342048 214200 342048 0 hellorld_do
rlabel metal2 236306 385336 236306 385336 0 io_in[0]
rlabel metal3 195944 346598 195944 346598 0 io_in[10]
rlabel metal2 519736 407232 519736 407232 0 io_in[11]
rlabel metal2 232792 404656 232792 404656 0 io_in[12]
rlabel metal4 238168 407583 238168 407583 0 io_in[13]
rlabel metal2 243544 407120 243544 407120 0 io_in[14]
rlabel metal2 233464 298816 233464 298816 0 io_in[15]
rlabel metal2 309960 118048 309960 118048 0 io_in[16]
rlabel metal2 451976 407176 451976 407176 0 io_in[17]
rlabel metal4 190568 498568 190568 498568 0 io_in[18]
rlabel metal2 237720 406280 237720 406280 0 io_in[19]
rlabel metal2 92456 300734 92456 300734 0 io_in[20]
rlabel metal3 188384 590184 188384 590184 0 io_in[21]
rlabel metal2 121576 593138 121576 593138 0 io_in[22]
rlabel metal2 55160 502754 55160 502754 0 io_in[23]
rlabel metal4 237944 301631 237944 301631 0 io_in[24]
rlabel metal3 3990 544824 3990 544824 0 io_in[25]
rlabel metal3 309624 154504 309624 154504 0 io_in[26]
rlabel metal2 4256 420000 4256 420000 0 io_in[27]
rlabel metal2 4200 416808 4200 416808 0 io_in[28]
rlabel metal2 236040 383880 236040 383880 0 io_in[29]
rlabel metal3 2310 333144 2310 333144 0 io_in[30]
rlabel metal3 2310 291032 2310 291032 0 io_in[31]
rlabel metal4 4088 247761 4088 247761 0 io_in[32]
rlabel metal3 2310 206360 2310 206360 0 io_in[33]
rlabel metal3 2310 164024 2310 164024 0 io_in[34]
rlabel metal3 2310 121688 2310 121688 0 io_in[35]
rlabel metal3 2310 79128 2310 79128 0 io_in[36]
rlabel metal3 2422 36904 2422 36904 0 io_in[37]
rlabel metal2 195160 408338 195160 408338 0 io_in[5]
rlabel metal3 195944 333158 195944 333158 0 io_in[6]
rlabel metal3 195944 336518 195944 336518 0 io_in[7]
rlabel metal3 518294 215768 518294 215768 0 io_in[8]
rlabel metal3 518182 218456 518182 218456 0 io_in[9]
rlabel metal3 234682 264376 234682 264376 0 io_oeb[0]
rlabel metal3 593306 430136 593306 430136 0 io_oeb[10]
rlabel metal3 593250 469672 593250 469672 0 io_oeb[11]
rlabel metal3 593194 509320 593194 509320 0 io_oeb[12]
rlabel metal3 593138 548968 593138 548968 0 io_oeb[13]
rlabel metal3 235466 280056 235466 280056 0 io_oeb[14]
rlabel metal3 234682 281176 234682 281176 0 io_oeb[15]
rlabel metal4 474376 590537 474376 590537 0 io_oeb[16]
rlabel metal4 190680 436683 190680 436683 0 io_oeb[17]
rlabel metal3 214522 284536 214522 284536 0 io_oeb[18]
rlabel metal2 190568 499744 190568 499744 0 io_oeb[19]
rlabel metal3 235410 265496 235410 265496 0 io_oeb[1]
rlabel metal2 209608 593026 209608 593026 0 io_oeb[20]
rlabel metal2 143416 441770 143416 441770 0 io_oeb[21]
rlabel metal2 77336 583002 77336 583002 0 io_oeb[22]
rlabel metal2 215992 300888 215992 300888 0 io_oeb[23]
rlabel metal3 2310 558936 2310 558936 0 io_oeb[24]
rlabel metal3 2366 516600 2366 516600 0 io_oeb[25]
rlabel metal4 141960 383880 141960 383880 0 io_oeb[26]
rlabel metal4 140280 363272 140280 363272 0 io_oeb[27]
rlabel metal3 2310 389592 2310 389592 0 io_oeb[28]
rlabel metal4 4200 346248 4200 346248 0 io_oeb[29]
rlabel metal3 235298 266616 235298 266616 0 io_oeb[2]
rlabel metal3 114366 304920 114366 304920 0 io_oeb[30]
rlabel metal3 236040 299222 236040 299222 0 io_oeb[31]
rlabel metal3 6510 220248 6510 220248 0 io_oeb[32]
rlabel metal4 27832 239624 27832 239624 0 io_oeb[33]
rlabel metal3 236040 302526 236040 302526 0 io_oeb[34]
rlabel metal4 29400 198408 29400 198408 0 io_oeb[35]
rlabel metal3 2366 51128 2366 51128 0 io_oeb[36]
rlabel metal3 2310 8792 2310 8792 0 io_oeb[37]
rlabel metal3 235466 267736 235466 267736 0 io_oeb[3]
rlabel metal3 593250 192360 593250 192360 0 io_oeb[4]
rlabel metal4 590184 235760 590184 235760 0 io_oeb[5]
rlabel metal3 235578 271096 235578 271096 0 io_oeb[6]
rlabel metal3 593138 311080 593138 311080 0 io_oeb[7]
rlabel metal3 593082 350728 593082 350728 0 io_oeb[8]
rlabel metal3 235410 274456 235410 274456 0 io_oeb[9]
rlabel metal2 237384 386470 237384 386470 0 io_out[0]
rlabel metal3 401632 399112 401632 399112 0 io_out[10]
rlabel metal2 565320 430248 565320 430248 0 io_out[11]
rlabel metal3 415968 402584 415968 402584 0 io_out[12]
rlabel metal2 563640 466648 563640 466648 0 io_out[13]
rlabel metal2 567000 490560 567000 490560 0 io_out[14]
rlabel metal2 562632 593474 562632 593474 0 io_out[15]
rlabel metal2 496664 593138 496664 593138 0 io_out[16]
rlabel metal2 430248 593082 430248 593082 0 io_out[17]
rlabel metal2 190344 499912 190344 499912 0 io_out[18]
rlabel metal4 192808 500192 192808 500192 0 io_out[19]
rlabel metal2 238280 387030 238280 387030 0 io_out[1]
rlabel metal2 190456 483000 190456 483000 0 io_out[20]
rlabel metal3 167272 590184 167272 590184 0 io_out[21]
rlabel metal2 99512 593082 99512 593082 0 io_out[22]
rlabel metal2 257992 388262 257992 388262 0 io_out[23]
rlabel metal2 258888 388318 258888 388318 0 io_out[24]
rlabel metal2 259784 395038 259784 395038 0 io_out[25]
rlabel metal2 260680 394310 260680 394310 0 io_out[26]
rlabel metal2 261576 393302 261576 393302 0 io_out[27]
rlabel metal2 262472 394814 262472 394814 0 io_out[28]
rlabel metal2 138600 373856 138600 373856 0 io_out[29]
rlabel metal3 590562 99848 590562 99848 0 io_out[2]
rlabel metal2 212520 352632 212520 352632 0 io_out[30]
rlabel metal3 17430 276696 17430 276696 0 io_out[31]
rlabel metal4 266056 384776 266056 384776 0 io_out[32]
rlabel metal2 266952 386302 266952 386302 0 io_out[33]
rlabel metal3 3990 149912 3990 149912 0 io_out[34]
rlabel metal2 31080 247072 31080 247072 0 io_out[35]
rlabel metal4 27720 225153 27720 225153 0 io_out[36]
rlabel metal3 5670 22904 5670 22904 0 io_out[37]
rlabel metal2 240072 387870 240072 387870 0 io_out[3]
rlabel metal2 240968 388094 240968 388094 0 io_out[4]
rlabel metal2 241864 386246 241864 386246 0 io_out[5]
rlabel metal2 242760 388150 242760 388150 0 io_out[6]
rlabel metal2 383880 342496 383880 342496 0 io_out[7]
rlabel metal2 380632 361648 380632 361648 0 io_out[8]
rlabel metal2 245448 388206 245448 388206 0 io_out[9]
rlabel metal3 235410 334936 235410 334936 0 mc14500_do\[0\]
rlabel metal3 236152 346010 236152 346010 0 mc14500_do\[10\]
rlabel metal2 493976 240030 493976 240030 0 mc14500_do\[11\]
rlabel metal2 495096 243390 495096 243390 0 mc14500_do\[12\]
rlabel metal2 496216 239190 496216 239190 0 mc14500_do\[13\]
rlabel metal2 497336 244174 497336 244174 0 mc14500_do\[14\]
rlabel metal3 235466 351736 235466 351736 0 mc14500_do\[15\]
rlabel metal2 499576 239974 499576 239974 0 mc14500_do\[16\]
rlabel metal2 500696 238406 500696 238406 0 mc14500_do\[17\]
rlabel metal2 501816 239134 501816 239134 0 mc14500_do\[18\]
rlabel metal3 236040 356090 236040 356090 0 mc14500_do\[19\]
rlabel metal3 233674 336056 233674 336056 0 mc14500_do\[1\]
rlabel metal3 231210 357336 231210 357336 0 mc14500_do\[20\]
rlabel metal3 232162 358456 232162 358456 0 mc14500_do\[21\]
rlabel metal3 231266 359576 231266 359576 0 mc14500_do\[22\]
rlabel metal3 234346 360696 234346 360696 0 mc14500_do\[23\]
rlabel metal2 223160 305648 223160 305648 0 mc14500_do\[24\]
rlabel metal2 228424 304528 228424 304528 0 mc14500_do\[25\]
rlabel metal2 510776 239078 510776 239078 0 mc14500_do\[26\]
rlabel metal2 225064 306488 225064 306488 0 mc14500_do\[27\]
rlabel metal3 233856 331800 233856 331800 0 mc14500_do\[28\]
rlabel metal2 514136 239862 514136 239862 0 mc14500_do\[29\]
rlabel metal3 233730 337176 233730 337176 0 mc14500_do\[2\]
rlabel metal2 515256 244062 515256 244062 0 mc14500_do\[30\]
rlabel metal3 236264 338114 236264 338114 0 mc14500_do\[3\]
rlabel metal2 486136 239246 486136 239246 0 mc14500_do\[4\]
rlabel metal2 229768 293384 229768 293384 0 mc14500_do\[5\]
rlabel metal2 224952 294896 224952 294896 0 mc14500_do\[6\]
rlabel metal3 234402 342776 234402 342776 0 mc14500_do\[7\]
rlabel metal2 490616 237342 490616 237342 0 mc14500_do\[8\]
rlabel metal2 491736 240702 491736 240702 0 mc14500_do\[9\]
rlabel metal2 278600 386358 278600 386358 0 mc14500_sram_addr\[0\]
rlabel metal2 279496 386078 279496 386078 0 mc14500_sram_addr\[1\]
rlabel metal2 280392 386134 280392 386134 0 mc14500_sram_addr\[2\]
rlabel metal4 281288 384944 281288 384944 0 mc14500_sram_addr\[3\]
rlabel metal2 282184 387030 282184 387030 0 mc14500_sram_addr\[4\]
rlabel metal4 283080 384888 283080 384888 0 mc14500_sram_addr\[5\]
rlabel metal3 517230 231896 517230 231896 0 mc14500_sram_gwe
rlabel metal2 283976 386302 283976 386302 0 mc14500_sram_in\[0\]
rlabel metal2 472920 291592 472920 291592 0 mc14500_sram_in\[1\]
rlabel metal2 494424 199122 494424 199122 0 mc14500_sram_in\[2\]
rlabel metal2 477960 291760 477960 291760 0 mc14500_sram_in\[3\]
rlabel metal4 287560 384863 287560 384863 0 mc14500_sram_in\[4\]
rlabel metal4 288456 384773 288456 384773 0 mc14500_sram_in\[5\]
rlabel metal4 289352 384593 289352 384593 0 mc14500_sram_in\[6\]
rlabel metal4 290248 384683 290248 384683 0 mc14500_sram_in\[7\]
rlabel metal2 326760 395024 326760 395024 0 pdp11_do\[0\]
rlabel metal2 335048 390334 335048 390334 0 pdp11_do\[10\]
rlabel metal2 336840 392798 336840 392798 0 pdp11_do\[11\]
rlabel metal3 387856 404600 387856 404600 0 pdp11_do\[12\]
rlabel metal3 391440 403144 391440 403144 0 pdp11_do\[13\]
rlabel metal2 447832 405482 447832 405482 0 pdp11_do\[14\]
rlabel metal2 453208 404082 453208 404082 0 pdp11_do\[15\]
rlabel metal3 402192 399560 402192 399560 0 pdp11_do\[16\]
rlabel metal2 347592 387534 347592 387534 0 pdp11_do\[17\]
rlabel metal2 468664 406364 468664 406364 0 pdp11_do\[18\]
rlabel metal2 351176 396046 351176 396046 0 pdp11_do\[19\]
rlabel metal2 377944 409010 377944 409010 0 pdp11_do\[1\]
rlabel metal2 352968 394478 352968 394478 0 pdp11_do\[20\]
rlabel metal2 354760 389438 354760 389438 0 pdp11_do\[21\]
rlabel metal2 356552 389326 356552 389326 0 pdp11_do\[22\]
rlabel metal2 358344 389382 358344 389382 0 pdp11_do\[23\]
rlabel metal3 500696 406840 500696 406840 0 pdp11_do\[24\]
rlabel metal2 361928 389214 361928 389214 0 pdp11_do\[25\]
rlabel metal3 438032 400792 438032 400792 0 pdp11_do\[26\]
rlabel metal2 517720 404026 517720 404026 0 pdp11_do\[27\]
rlabel metal2 523096 404754 523096 404754 0 pdp11_do\[28\]
rlabel metal3 448280 404376 448280 404376 0 pdp11_do\[29\]
rlabel metal2 383320 401114 383320 401114 0 pdp11_do\[2\]
rlabel metal3 452368 402920 452368 402920 0 pdp11_do\[30\]
rlabel metal2 539224 401226 539224 401226 0 pdp11_do\[31\]
rlabel metal2 374472 395990 374472 395990 0 pdp11_do\[32\]
rlabel metal3 355600 402248 355600 402248 0 pdp11_do\[3\]
rlabel metal3 359184 406280 359184 406280 0 pdp11_do\[4\]
rlabel metal2 326088 389494 326088 389494 0 pdp11_do\[5\]
rlabel metal2 327880 395318 327880 395318 0 pdp11_do\[6\]
rlabel metal2 329672 389102 329672 389102 0 pdp11_do\[7\]
rlabel metal2 331464 393470 331464 393470 0 pdp11_do\[8\]
rlabel metal2 333256 388374 333256 388374 0 pdp11_do\[9\]
rlabel metal3 434560 397768 434560 397768 0 pdp11_oeb\[0\]
rlabel metal2 335944 392574 335944 392574 0 pdp11_oeb\[10\]
rlabel metal2 337736 389942 337736 389942 0 pdp11_oeb\[11\]
rlabel metal3 550662 471016 550662 471016 0 pdp11_oeb\[12\]
rlabel metal3 549752 475594 549752 475594 0 pdp11_oeb\[13\]
rlabel metal2 343112 390110 343112 390110 0 pdp11_oeb\[14\]
rlabel metal2 344904 390222 344904 390222 0 pdp11_oeb\[15\]
rlabel metal2 346696 390166 346696 390166 0 pdp11_oeb\[16\]
rlabel metal3 452536 402696 452536 402696 0 pdp11_oeb\[17\]
rlabel metal2 350280 390950 350280 390950 0 pdp11_oeb\[18\]
rlabel metal2 352072 391006 352072 391006 0 pdp11_oeb\[19\]
rlabel metal3 435008 400680 435008 400680 0 pdp11_oeb\[1\]
rlabel metal2 353864 395038 353864 395038 0 pdp11_oeb\[20\]
rlabel metal2 355656 397782 355656 397782 0 pdp11_oeb\[21\]
rlabel metal2 357448 388262 357448 388262 0 pdp11_oeb\[22\]
rlabel metal2 359240 395878 359240 395878 0 pdp11_oeb\[23\]
rlabel metal2 361032 390278 361032 390278 0 pdp11_oeb\[24\]
rlabel metal2 362824 397838 362824 397838 0 pdp11_oeb\[25\]
rlabel metal2 364616 389102 364616 389102 0 pdp11_oeb\[26\]
rlabel metal3 551446 541576 551446 541576 0 pdp11_oeb\[27\]
rlabel metal3 554232 451976 554232 451976 0 pdp11_oeb\[28\]
rlabel metal2 369992 390726 369992 390726 0 pdp11_oeb\[29\]
rlabel metal3 550830 423976 550830 423976 0 pdp11_oeb\[2\]
rlabel metal2 421624 390096 421624 390096 0 pdp11_oeb\[30\]
rlabel metal2 373576 387534 373576 387534 0 pdp11_oeb\[31\]
rlabel metal2 375368 387030 375368 387030 0 pdp11_oeb\[32\]
rlabel metal3 552454 428680 552454 428680 0 pdp11_oeb\[3\]
rlabel metal2 330904 392448 330904 392448 0 pdp11_oeb\[4\]
rlabel metal2 326984 387590 326984 387590 0 pdp11_oeb\[5\]
rlabel metal2 328776 397614 328776 397614 0 pdp11_oeb\[6\]
rlabel metal2 330568 387814 330568 387814 0 pdp11_oeb\[7\]
rlabel metal2 332360 397670 332360 397670 0 pdp11_oeb\[8\]
rlabel metal2 334152 387422 334152 387422 0 pdp11_oeb\[9\]
rlabel metal2 326984 225106 326984 225106 0 qcpu_do\[0\]
rlabel metal2 335944 224266 335944 224266 0 qcpu_do\[10\]
rlabel metal2 336840 255710 336840 255710 0 qcpu_do\[11\]
rlabel metal2 337736 205842 337736 205842 0 qcpu_do\[12\]
rlabel metal2 338632 205786 338632 205786 0 qcpu_do\[13\]
rlabel metal3 434504 187432 434504 187432 0 qcpu_do\[14\]
rlabel metal3 435624 163912 435624 163912 0 qcpu_do\[15\]
rlabel metal3 434000 185640 434000 185640 0 qcpu_do\[16\]
rlabel metal3 437864 168840 437864 168840 0 qcpu_do\[17\]
rlabel metal3 344176 252056 344176 252056 0 qcpu_do\[18\]
rlabel metal3 440104 236824 440104 236824 0 qcpu_do\[19\]
rlabel metal2 327880 219226 327880 219226 0 qcpu_do\[1\]
rlabel metal2 344904 227570 344904 227570 0 qcpu_do\[20\]
rlabel metal2 538888 165270 538888 165270 0 qcpu_do\[21\]
rlabel metal2 540232 153622 540232 153622 0 qcpu_do\[22\]
rlabel metal2 541576 153566 541576 153566 0 qcpu_do\[23\]
rlabel metal2 542920 153510 542920 153510 0 qcpu_do\[24\]
rlabel metal2 544264 172830 544264 172830 0 qcpu_do\[25\]
rlabel metal2 350280 216650 350280 216650 0 qcpu_do\[26\]
rlabel metal2 351176 215810 351176 215810 0 qcpu_do\[27\]
rlabel metal2 352072 214970 352072 214970 0 qcpu_do\[28\]
rlabel metal2 352968 225050 352968 225050 0 qcpu_do\[29\]
rlabel metal2 328776 213346 328776 213346 0 qcpu_do\[2\]
rlabel metal2 353864 224210 353864 224210 0 qcpu_do\[30\]
rlabel metal2 354760 221690 354760 221690 0 qcpu_do\[31\]
rlabel metal3 356328 252056 356328 252056 0 qcpu_do\[32\]
rlabel metal2 329672 207522 329672 207522 0 qcpu_do\[3\]
rlabel metal2 330568 227626 330568 227626 0 qcpu_do\[4\]
rlabel metal2 331464 222530 331464 222530 0 qcpu_do\[5\]
rlabel metal3 332920 252056 332920 252056 0 qcpu_do\[6\]
rlabel metal2 333256 207466 333256 207466 0 qcpu_do\[7\]
rlabel metal3 334656 252056 334656 252056 0 qcpu_do\[8\]
rlabel metal2 335048 207410 335048 207410 0 qcpu_do\[9\]
rlabel metal4 564424 57839 564424 57839 0 qcpu_oeb\[0\]
rlabel metal4 564648 209496 564648 209496 0 qcpu_oeb\[10\]
rlabel metal4 566328 210840 566328 210840 0 qcpu_oeb\[11\]
rlabel metal4 564760 212184 564760 212184 0 qcpu_oeb\[12\]
rlabel metal4 566216 213528 566216 213528 0 qcpu_oeb\[13\]
rlabel metal4 568008 214872 568008 214872 0 qcpu_oeb\[14\]
rlabel metal3 377790 352184 377790 352184 0 qcpu_oeb\[15\]
rlabel metal4 564872 217560 564872 217560 0 qcpu_oeb\[16\]
rlabel metal4 566440 218904 566440 218904 0 qcpu_oeb\[17\]
rlabel metal4 569688 220248 569688 220248 0 qcpu_oeb\[18\]
rlabel metal4 569576 221592 569576 221592 0 qcpu_oeb\[19\]
rlabel metal3 564424 58576 564424 58576 0 qcpu_oeb\[1\]
rlabel metal4 571256 222936 571256 222936 0 qcpu_oeb\[20\]
rlabel metal4 571368 224280 571368 224280 0 qcpu_oeb\[21\]
rlabel metal4 566552 225624 566552 225624 0 qcpu_oeb\[22\]
rlabel metal3 377790 361144 377790 361144 0 qcpu_oeb\[23\]
rlabel metal3 566454 94360 566454 94360 0 qcpu_oeb\[24\]
rlabel metal4 571480 229656 571480 229656 0 qcpu_oeb\[25\]
rlabel metal3 377790 364504 377790 364504 0 qcpu_oeb\[26\]
rlabel metal3 566510 99064 566510 99064 0 qcpu_oeb\[27\]
rlabel metal4 568232 233688 568232 233688 0 qcpu_oeb\[28\]
rlabel metal3 567350 102200 567350 102200 0 qcpu_oeb\[29\]
rlabel metal4 425880 193984 425880 193984 0 qcpu_oeb\[2\]
rlabel metal3 566566 103768 566566 103768 0 qcpu_oeb\[30\]
rlabel metal4 571592 237048 571592 237048 0 qcpu_oeb\[31\]
rlabel metal4 562856 113904 562856 113904 0 qcpu_oeb\[32\]
rlabel metal3 567294 61432 567294 61432 0 qcpu_oeb\[3\]
rlabel metal4 562968 105504 562968 105504 0 qcpu_oeb\[4\]
rlabel metal4 563080 106344 563080 106344 0 qcpu_oeb\[5\]
rlabel metal4 540120 245392 540120 245392 0 qcpu_oeb\[6\]
rlabel metal3 467726 343224 467726 343224 0 qcpu_oeb\[7\]
rlabel metal4 563304 200536 563304 200536 0 qcpu_oeb\[8\]
rlabel metal3 467782 345464 467782 345464 0 qcpu_oeb\[9\]
rlabel metal2 356552 208306 356552 208306 0 qcpu_sram_addr\[0\]
rlabel metal2 357448 209930 357448 209930 0 qcpu_sram_addr\[1\]
rlabel metal2 358344 209090 358344 209090 0 qcpu_sram_addr\[2\]
rlabel metal2 359240 255710 359240 255710 0 qcpu_sram_addr\[3\]
rlabel metal2 360136 208250 360136 208250 0 qcpu_sram_addr\[4\]
rlabel metal2 562856 119392 562856 119392 0 qcpu_sram_addr\[5\]
rlabel metal2 563192 156744 563192 156744 0 qcpu_sram_gwe
rlabel metal2 566216 142520 566216 142520 0 qcpu_sram_in\[0\]
rlabel metal2 562968 144200 562968 144200 0 qcpu_sram_in\[1\]
rlabel metal2 523320 202720 523320 202720 0 qcpu_sram_in\[2\]
rlabel metal2 564648 136472 564648 136472 0 qcpu_sram_in\[3\]
rlabel metal2 376040 213864 376040 213864 0 qcpu_sram_in\[4\]
rlabel metal2 563304 138152 563304 138152 0 qcpu_sram_in\[5\]
rlabel metal2 368200 203266 368200 203266 0 qcpu_sram_in\[6\]
rlabel metal2 548520 201880 548520 201880 0 qcpu_sram_in\[7\]
rlabel metal2 566328 141232 566328 141232 0 qcpu_sram_out\[0\]
rlabel metal2 561288 140728 561288 140728 0 qcpu_sram_out\[1\]
rlabel metal2 564760 142128 564760 142128 0 qcpu_sram_out\[2\]
rlabel metal2 561512 142184 561512 142184 0 qcpu_sram_out\[3\]
rlabel metal2 561176 144424 561176 144424 0 qcpu_sram_out\[4\]
rlabel metal2 467880 289184 467880 289184 0 qcpu_sram_out\[5\]
rlabel metal2 561400 147616 561400 147616 0 qcpu_sram_out\[6\]
rlabel metal2 514878 200088 514878 200088 0 qcpu_sram_out\[7\]
rlabel metal2 376376 382200 376376 382200 0 rst_ay8913
rlabel metal2 235032 301728 235032 301728 0 rst_blinker
rlabel metal2 172872 287910 172872 287910 0 rst_hellorld
rlabel metal3 518070 205016 518070 205016 0 rst_mc14500
rlabel metal3 189714 421736 189714 421736 0 rst_pdp11
rlabel metal4 220024 273448 220024 273448 0 rst_qcpu
rlabel metal2 212296 49322 212296 49322 0 rst_sid
rlabel metal3 358890 84952 358890 84952 0 rst_sn76489
rlabel metal3 217546 371896 217546 371896 0 rst_tbb1143
rlabel metal3 234570 308056 234570 308056 0 sid_do\[0\]
rlabel metal3 234234 319256 234234 319256 0 sid_do\[10\]
rlabel metal4 272440 210560 272440 210560 0 sid_do\[11\]
rlabel metal2 269528 210952 269528 210952 0 sid_do\[12\]
rlabel metal3 271390 186648 271390 186648 0 sid_do\[13\]
rlabel metal3 271166 189560 271166 189560 0 sid_do\[14\]
rlabel metal3 271222 192472 271222 192472 0 sid_do\[15\]
rlabel metal3 232218 325976 232218 325976 0 sid_do\[16\]
rlabel metal3 233002 327096 233002 327096 0 sid_do\[17\]
rlabel metal3 231378 328216 231378 328216 0 sid_do\[18\]
rlabel metal3 235242 329336 235242 329336 0 sid_do\[19\]
rlabel metal3 234626 309176 234626 309176 0 sid_do\[1\]
rlabel metal3 235522 330456 235522 330456 0 sid_do\[20\]
rlabel metal3 234514 310296 234514 310296 0 sid_do\[2\]
rlabel metal3 234402 311416 234402 311416 0 sid_do\[3\]
rlabel metal3 234458 312536 234458 312536 0 sid_do\[4\]
rlabel metal3 234290 313656 234290 313656 0 sid_do\[5\]
rlabel metal3 234346 314776 234346 314776 0 sid_do\[6\]
rlabel metal3 234570 315896 234570 315896 0 sid_do\[7\]
rlabel metal3 234682 317016 234682 317016 0 sid_do\[8\]
rlabel metal3 234626 318136 234626 318136 0 sid_do\[9\]
rlabel metal2 154952 212086 154952 212086 0 sid_oeb
rlabel metal2 304920 192864 304920 192864 0 sn76489_do\[0\]
rlabel metal2 310856 254450 310856 254450 0 sn76489_do\[10\]
rlabel metal2 311752 193970 311752 193970 0 sn76489_do\[11\]
rlabel metal2 312648 254506 312648 254506 0 sn76489_do\[12\]
rlabel metal2 313544 254058 313544 254058 0 sn76489_do\[13\]
rlabel metal2 314440 230090 314440 230090 0 sn76489_do\[14\]
rlabel metal3 354144 138600 354144 138600 0 sn76489_do\[15\]
rlabel metal3 356664 232904 356664 232904 0 sn76489_do\[16\]
rlabel metal2 396984 175518 396984 175518 0 sn76489_do\[17\]
rlabel metal2 399000 122542 399000 122542 0 sn76489_do\[18\]
rlabel metal2 401016 162862 401016 162862 0 sn76489_do\[19\]
rlabel metal2 302792 190722 302792 190722 0 sn76489_do\[1\]
rlabel metal2 403032 174678 403032 174678 0 sn76489_do\[20\]
rlabel metal2 405048 121310 405048 121310 0 sn76489_do\[21\]
rlabel metal2 407064 172158 407064 172158 0 sn76489_do\[22\]
rlabel metal2 407400 179312 407400 179312 0 sn76489_do\[23\]
rlabel metal2 323400 239386 323400 239386 0 sn76489_do\[24\]
rlabel metal3 368704 217672 368704 217672 0 sn76489_do\[25\]
rlabel metal2 326872 242480 326872 242480 0 sn76489_do\[26\]
rlabel metal3 329000 252056 329000 252056 0 sn76489_do\[27\]
rlabel metal2 303688 190666 303688 190666 0 sn76489_do\[2\]
rlabel metal3 307328 252056 307328 252056 0 sn76489_do\[3\]
rlabel metal2 305480 226730 305480 226730 0 sn76489_do\[4\]
rlabel metal2 306376 236922 306376 236922 0 sn76489_do\[5\]
rlabel metal2 307272 191506 307272 191506 0 sn76489_do\[6\]
rlabel metal2 308168 191450 308168 191450 0 sn76489_do\[7\]
rlabel metal2 378840 121310 378840 121310 0 sn76489_do\[8\]
rlabel metal2 380856 121758 380856 121758 0 sn76489_do\[9\]
rlabel metal3 197582 349608 197582 349608 0 tbb1143_do\[0\]
rlabel metal3 197694 352968 197694 352968 0 tbb1143_do\[1\]
rlabel metal3 197638 356328 197638 356328 0 tbb1143_do\[2\]
rlabel metal3 197750 359688 197750 359688 0 tbb1143_do\[3\]
rlabel metal3 217882 377496 217882 377496 0 tbb1143_do\[4\]
rlabel metal3 580160 4200 580160 4200 0 user_irq[0]
rlabel metal2 429240 197064 429240 197064 0 user_irq[1]
rlabel metal3 583744 4200 583744 4200 0 user_irq[2]
rlabel metal2 97384 49378 97384 49378 0 wb_clk_i
rlabel metal2 242984 237384 242984 237384 0 wb_rst_i
rlabel metal3 376166 298424 376166 298424 0 wbs_ack_o
rlabel metal2 22792 112406 22792 112406 0 wbs_adr_i[0]
rlabel metal3 177352 47880 177352 47880 0 wbs_adr_i[10]
rlabel metal2 93240 24206 93240 24206 0 wbs_adr_i[11]
rlabel metal2 98952 22582 98952 22582 0 wbs_adr_i[12]
rlabel metal2 256200 253106 256200 253106 0 wbs_adr_i[13]
rlabel metal2 257096 251034 257096 251034 0 wbs_adr_i[14]
rlabel metal2 116088 20958 116088 20958 0 wbs_adr_i[15]
rlabel metal2 121800 17654 121800 17654 0 wbs_adr_i[16]
rlabel metal4 259784 252947 259784 252947 0 wbs_adr_i[17]
rlabel metal4 260680 252857 260680 252857 0 wbs_adr_i[18]
rlabel metal2 138936 22750 138936 22750 0 wbs_adr_i[19]
rlabel metal2 30408 105630 30408 105630 0 wbs_adr_i[1]
rlabel metal2 144648 15862 144648 15862 0 wbs_adr_i[20]
rlabel metal2 263368 254562 263368 254562 0 wbs_adr_i[21]
rlabel metal2 264264 254674 264264 254674 0 wbs_adr_i[22]
rlabel metal2 161784 19950 161784 19950 0 wbs_adr_i[23]
rlabel metal2 167496 25102 167496 25102 0 wbs_adr_i[24]
rlabel metal2 266952 254058 266952 254058 0 wbs_adr_i[25]
rlabel metal3 228256 48216 228256 48216 0 wbs_adr_i[26]
rlabel metal3 231056 46200 231056 46200 0 wbs_adr_i[27]
rlabel metal2 190568 3262 190568 3262 0 wbs_adr_i[28]
rlabel metal2 196056 12502 196056 12502 0 wbs_adr_i[29]
rlabel metal3 142184 232792 142184 232792 0 wbs_adr_i[2]
rlabel metal2 201768 7462 201768 7462 0 wbs_adr_i[30]
rlabel metal2 279160 148624 279160 148624 0 wbs_adr_i[31]
rlabel metal2 45640 2646 45640 2646 0 wbs_adr_i[3]
rlabel metal2 53256 2366 53256 2366 0 wbs_adr_i[4]
rlabel metal4 52024 117824 52024 117824 0 wbs_adr_i[5]
rlabel metal4 51912 110208 51912 110208 0 wbs_adr_i[6]
rlabel metal2 70392 2310 70392 2310 0 wbs_adr_i[7]
rlabel metal2 76104 18270 76104 18270 0 wbs_adr_i[8]
rlabel metal2 81816 17542 81816 17542 0 wbs_adr_i[9]
rlabel metal3 376278 296184 376278 296184 0 wbs_cyc_i
rlabel metal2 24696 121534 24696 121534 0 wbs_dat_i[0]
rlabel metal2 282184 144466 282184 144466 0 wbs_dat_i[10]
rlabel metal2 95144 9926 95144 9926 0 wbs_dat_i[11]
rlabel metal2 101080 3150 101080 3150 0 wbs_dat_i[12]
rlabel metal2 284872 131810 284872 131810 0 wbs_dat_i[13]
rlabel metal2 285768 131866 285768 131866 0 wbs_dat_i[14]
rlabel metal2 118216 4102 118216 4102 0 wbs_dat_i[15]
rlabel metal2 123704 9086 123704 9086 0 wbs_dat_i[16]
rlabel metal2 288456 136066 288456 136066 0 wbs_dat_i[17]
rlabel metal3 288736 252056 288736 252056 0 wbs_dat_i[18]
rlabel metal2 140840 7406 140840 7406 0 wbs_dat_i[19]
rlabel metal3 153216 234472 153216 234472 0 wbs_dat_i[1]
rlabel metal2 146552 13230 146552 13230 0 wbs_dat_i[20]
rlabel metal2 290024 141736 290024 141736 0 wbs_dat_i[21]
rlabel metal2 158200 3206 158200 3206 0 wbs_dat_i[22]
rlabel metal2 163688 6510 163688 6510 0 wbs_dat_i[23]
rlabel metal2 169400 14966 169400 14966 0 wbs_dat_i[24]
rlabel metal2 284984 147392 284984 147392 0 wbs_dat_i[25]
rlabel metal2 288344 151592 288344 151592 0 wbs_dat_i[26]
rlabel metal2 186536 10710 186536 10710 0 wbs_dat_i[27]
rlabel metal2 192248 19390 192248 19390 0 wbs_dat_i[28]
rlabel metal2 281400 150584 281400 150584 0 wbs_dat_i[29]
rlabel metal3 39256 4200 39256 4200 0 wbs_dat_i[2]
rlabel metal2 283416 147336 283416 147336 0 wbs_dat_i[30]
rlabel metal2 209384 18326 209384 18326 0 wbs_dat_i[31]
rlabel metal2 47544 8190 47544 8190 0 wbs_dat_i[3]
rlabel metal2 55160 9030 55160 9030 0 wbs_dat_i[4]
rlabel metal2 60872 9870 60872 9870 0 wbs_dat_i[5]
rlabel metal2 68936 7000 68936 7000 0 wbs_dat_i[6]
rlabel metal2 72296 12390 72296 12390 0 wbs_dat_i[7]
rlabel metal2 78008 7350 78008 7350 0 wbs_dat_i[8]
rlabel metal2 281288 142730 281288 142730 0 wbs_dat_i[9]
rlabel metal3 376110 259224 376110 259224 0 wbs_dat_o[0]
rlabel metal2 91336 24990 91336 24990 0 wbs_dat_o[10]
rlabel metal2 97048 20846 97048 20846 0 wbs_dat_o[11]
rlabel metal2 102760 16590 102760 16590 0 wbs_dat_o[12]
rlabel metal2 359240 144480 359240 144480 0 wbs_dat_o[13]
rlabel metal2 114408 2310 114408 2310 0 wbs_dat_o[14]
rlabel metal2 119896 19222 119896 19222 0 wbs_dat_o[15]
rlabel metal2 125832 2646 125832 2646 0 wbs_dat_o[16]
rlabel metal2 131544 4830 131544 4830 0 wbs_dat_o[17]
rlabel metal3 377342 279384 377342 279384 0 wbs_dat_o[18]
rlabel metal3 376502 280504 376502 280504 0 wbs_dat_o[19]
rlabel metal3 376446 260344 376446 260344 0 wbs_dat_o[1]
rlabel metal3 376222 281624 376222 281624 0 wbs_dat_o[20]
rlabel metal3 377006 282744 377006 282744 0 wbs_dat_o[21]
rlabel metal4 359016 147187 359016 147187 0 wbs_dat_o[22]
rlabel metal2 165816 2478 165816 2478 0 wbs_dat_o[23]
rlabel metal5 374584 286110 374584 286110 0 wbs_dat_o[24]
rlabel metal3 331800 256088 331800 256088 0 wbs_dat_o[25]
rlabel metal5 374528 288270 374528 288270 0 wbs_dat_o[26]
rlabel metal2 188440 21630 188440 21630 0 wbs_dat_o[27]
rlabel metal3 376390 290584 376390 290584 0 wbs_dat_o[28]
rlabel metal3 377230 291704 377230 291704 0 wbs_dat_o[29]
rlabel metal3 376054 261464 376054 261464 0 wbs_dat_o[2]
rlabel metal3 350504 256032 350504 256032 0 wbs_dat_o[30]
rlabel metal2 211288 17710 211288 17710 0 wbs_dat_o[31]
rlabel metal2 49448 2422 49448 2422 0 wbs_dat_o[3]
rlabel metal3 377454 263704 377454 263704 0 wbs_dat_o[4]
rlabel metal3 377342 264824 377342 264824 0 wbs_dat_o[5]
rlabel metal4 375256 261897 375256 261897 0 wbs_dat_o[6]
rlabel metal3 377286 267064 377286 267064 0 wbs_dat_o[7]
rlabel metal2 355432 137872 355432 137872 0 wbs_dat_o[8]
rlabel metal3 377510 269304 377510 269304 0 wbs_dat_o[9]
rlabel metal3 376558 297304 376558 297304 0 wbs_stb_i
rlabel metal2 20888 108990 20888 108990 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 596040 596040
<< end >>
