magic
tech gf180mcuD
magscale 1 10
timestamp 1702341368
<< nwell >>
rect 1258 44281 46678 44774
rect 1258 44256 25725 44281
rect 1258 43527 6685 43552
rect 1258 42713 46678 43527
rect 1258 42688 16541 42713
rect 1258 41959 6685 41984
rect 1258 41145 46678 41959
rect 1258 41120 10829 41145
rect 1258 40391 6909 40416
rect 1258 39577 46678 40391
rect 1258 39552 2541 39577
rect 1258 38823 6125 38848
rect 1258 38009 46678 38823
rect 1258 37984 21395 38009
rect 1258 37255 3592 37280
rect 1258 36441 46678 37255
rect 1258 36416 7512 36441
rect 1258 35687 2541 35712
rect 1258 34873 46678 35687
rect 1258 34848 8597 34873
rect 1258 34119 23392 34144
rect 1258 33305 46678 34119
rect 1258 33280 2541 33305
rect 1258 32551 13784 32576
rect 1258 31737 46678 32551
rect 1258 31712 2541 31737
rect 1258 30983 12328 31008
rect 1258 30169 46678 30983
rect 1258 30144 3592 30169
rect 1258 29415 4445 29440
rect 1258 28601 46678 29415
rect 1258 28576 3592 28601
rect 1258 27847 14749 27872
rect 1258 27033 46678 27847
rect 1258 27008 2541 27033
rect 1258 26279 6461 26304
rect 1258 25465 46678 26279
rect 1258 25440 3592 25465
rect 1258 24711 11837 24736
rect 1258 23897 46678 24711
rect 1258 23872 10536 23897
rect 1258 23143 2541 23168
rect 1258 22329 46678 23143
rect 1258 22304 8632 22329
rect 1258 21575 2541 21600
rect 1258 20761 46678 21575
rect 1258 20736 6685 20761
rect 1258 20007 21245 20032
rect 1258 19193 46678 20007
rect 1258 19168 2541 19193
rect 1258 18439 2541 18464
rect 1258 17625 46678 18439
rect 1258 17600 10829 17625
rect 1258 16871 2541 16896
rect 1258 16057 46678 16871
rect 1258 16032 24717 16057
rect 1258 15303 2541 15328
rect 1258 14489 46678 15303
rect 1258 14464 7805 14489
rect 1258 13735 2541 13760
rect 1258 12921 46678 13735
rect 1258 12896 17101 12921
rect 1258 12167 2541 12192
rect 1258 11353 46678 12167
rect 1258 11328 7960 11353
rect 1258 10599 2877 10624
rect 1258 9785 46678 10599
rect 1258 9760 2541 9785
rect 1258 9031 18221 9056
rect 1258 8217 46678 9031
rect 1258 8192 6461 8217
rect 1258 7463 3592 7488
rect 1258 6649 46678 7463
rect 1258 6624 8925 6649
rect 1258 5895 2541 5920
rect 1258 5081 46678 5895
rect 1258 5056 10829 5081
rect 1258 4327 6056 4352
rect 1258 3513 46678 4327
rect 1258 3488 10493 3513
<< pwell >>
rect 1258 43552 46678 44256
rect 1258 41984 46678 42688
rect 1258 40416 46678 41120
rect 1258 38848 46678 39552
rect 1258 37280 46678 37984
rect 1258 35712 46678 36416
rect 1258 34144 46678 34848
rect 1258 32576 46678 33280
rect 1258 31008 46678 31712
rect 1258 29440 46678 30144
rect 1258 27872 46678 28576
rect 1258 26304 46678 27008
rect 1258 24736 46678 25440
rect 1258 23168 46678 23872
rect 1258 21600 46678 22304
rect 1258 20032 46678 20736
rect 1258 18464 46678 19168
rect 1258 16896 46678 17600
rect 1258 15328 46678 16032
rect 1258 13760 46678 14464
rect 1258 12192 46678 12896
rect 1258 10624 46678 11328
rect 1258 9056 46678 9760
rect 1258 7488 46678 8192
rect 1258 5920 46678 6624
rect 1258 4352 46678 5056
rect 1258 3050 46678 3488
<< obsm1 >>
rect 1344 3076 46592 44882
<< metal2 >>
rect 6048 47200 6160 48000
rect 17920 47200 18032 48000
rect 29792 47200 29904 48000
rect 41664 47200 41776 48000
rect 2688 0 2800 800
rect 4256 0 4368 800
rect 5824 0 5936 800
rect 7392 0 7504 800
rect 8960 0 9072 800
rect 10528 0 10640 800
rect 12096 0 12208 800
rect 13664 0 13776 800
rect 15232 0 15344 800
rect 16800 0 16912 800
rect 18368 0 18480 800
rect 19936 0 20048 800
rect 21504 0 21616 800
rect 23072 0 23184 800
rect 24640 0 24752 800
rect 26208 0 26320 800
rect 27776 0 27888 800
rect 29344 0 29456 800
rect 30912 0 31024 800
rect 32480 0 32592 800
rect 34048 0 34160 800
rect 35616 0 35728 800
rect 37184 0 37296 800
rect 38752 0 38864 800
rect 40320 0 40432 800
rect 41888 0 42000 800
rect 43456 0 43568 800
rect 45024 0 45136 800
<< obsm2 >>
rect 1708 47140 5988 47200
rect 6220 47140 17860 47200
rect 18092 47140 29732 47200
rect 29964 47140 41604 47200
rect 41836 47140 46900 47200
rect 1708 860 46900 47140
rect 1708 800 2628 860
rect 2860 800 4196 860
rect 4428 800 5764 860
rect 5996 800 7332 860
rect 7564 800 8900 860
rect 9132 800 10468 860
rect 10700 800 12036 860
rect 12268 800 13604 860
rect 13836 800 15172 860
rect 15404 800 16740 860
rect 16972 800 18308 860
rect 18540 800 19876 860
rect 20108 800 21444 860
rect 21676 800 23012 860
rect 23244 800 24580 860
rect 24812 800 26148 860
rect 26380 800 27716 860
rect 27948 800 29284 860
rect 29516 800 30852 860
rect 31084 800 32420 860
rect 32652 800 33988 860
rect 34220 800 35556 860
rect 35788 800 37124 860
rect 37356 800 38692 860
rect 38924 800 40260 860
rect 40492 800 41828 860
rect 42060 800 43396 860
rect 43628 800 44964 860
rect 45196 800 46900 860
<< metal3 >>
rect 47200 45024 48000 45136
rect 47200 40320 48000 40432
rect 47200 35616 48000 35728
rect 47200 30912 48000 31024
rect 47200 26208 48000 26320
rect 47200 21504 48000 21616
rect 47200 16800 48000 16912
rect 47200 12096 48000 12208
rect 47200 7392 48000 7504
rect 47200 2688 48000 2800
<< obsm3 >>
rect 1698 44964 47140 45108
rect 1698 40492 47348 44964
rect 1698 40260 47140 40492
rect 1698 35788 47348 40260
rect 1698 35556 47140 35788
rect 1698 31084 47348 35556
rect 1698 30852 47140 31084
rect 1698 26380 47348 30852
rect 1698 26148 47140 26380
rect 1698 21676 47348 26148
rect 1698 21444 47140 21676
rect 1698 16972 47348 21444
rect 1698 16740 47140 16972
rect 1698 12268 47348 16740
rect 1698 12036 47140 12268
rect 1698 7564 47348 12036
rect 1698 7332 47140 7564
rect 1698 2860 47348 7332
rect 1698 2716 47140 2860
<< metal4 >>
rect 4448 3076 4768 44748
rect 19808 3076 20128 44748
rect 35168 3076 35488 44748
<< obsm4 >>
rect 8428 3602 19748 44334
rect 20188 3602 35108 44334
rect 35548 3602 45892 44334
<< labels >>
rlabel metal3 s 47200 40320 48000 40432 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 47200 45024 48000 45136 6 custom_settings[1]
port 2 nsew signal input
rlabel metal3 s 47200 2688 48000 2800 6 io_in_1[0]
port 3 nsew signal input
rlabel metal3 s 47200 7392 48000 7504 6 io_in_1[1]
port 4 nsew signal input
rlabel metal3 s 47200 12096 48000 12208 6 io_in_1[2]
port 5 nsew signal input
rlabel metal3 s 47200 16800 48000 16912 6 io_in_1[3]
port 6 nsew signal input
rlabel metal3 s 47200 21504 48000 21616 6 io_in_1[4]
port 7 nsew signal input
rlabel metal3 s 47200 26208 48000 26320 6 io_in_1[5]
port 8 nsew signal input
rlabel metal3 s 47200 30912 48000 31024 6 io_in_1[6]
port 9 nsew signal input
rlabel metal3 s 47200 35616 48000 35728 6 io_in_1[7]
port 10 nsew signal input
rlabel metal2 s 29792 47200 29904 48000 6 io_in_2[0]
port 11 nsew signal input
rlabel metal2 s 41664 47200 41776 48000 6 io_in_2[1]
port 12 nsew signal input
rlabel metal2 s 2688 0 2800 800 6 io_out[0]
port 13 nsew signal output
rlabel metal2 s 18368 0 18480 800 6 io_out[10]
port 14 nsew signal output
rlabel metal2 s 19936 0 20048 800 6 io_out[11]
port 15 nsew signal output
rlabel metal2 s 21504 0 21616 800 6 io_out[12]
port 16 nsew signal output
rlabel metal2 s 23072 0 23184 800 6 io_out[13]
port 17 nsew signal output
rlabel metal2 s 24640 0 24752 800 6 io_out[14]
port 18 nsew signal output
rlabel metal2 s 26208 0 26320 800 6 io_out[15]
port 19 nsew signal output
rlabel metal2 s 27776 0 27888 800 6 io_out[16]
port 20 nsew signal output
rlabel metal2 s 29344 0 29456 800 6 io_out[17]
port 21 nsew signal output
rlabel metal2 s 30912 0 31024 800 6 io_out[18]
port 22 nsew signal output
rlabel metal2 s 32480 0 32592 800 6 io_out[19]
port 23 nsew signal output
rlabel metal2 s 4256 0 4368 800 6 io_out[1]
port 24 nsew signal output
rlabel metal2 s 34048 0 34160 800 6 io_out[20]
port 25 nsew signal output
rlabel metal2 s 35616 0 35728 800 6 io_out[21]
port 26 nsew signal output
rlabel metal2 s 37184 0 37296 800 6 io_out[22]
port 27 nsew signal output
rlabel metal2 s 38752 0 38864 800 6 io_out[23]
port 28 nsew signal output
rlabel metal2 s 40320 0 40432 800 6 io_out[24]
port 29 nsew signal output
rlabel metal2 s 41888 0 42000 800 6 io_out[25]
port 30 nsew signal output
rlabel metal2 s 43456 0 43568 800 6 io_out[26]
port 31 nsew signal output
rlabel metal2 s 45024 0 45136 800 6 io_out[27]
port 32 nsew signal output
rlabel metal2 s 5824 0 5936 800 6 io_out[2]
port 33 nsew signal output
rlabel metal2 s 7392 0 7504 800 6 io_out[3]
port 34 nsew signal output
rlabel metal2 s 8960 0 9072 800 6 io_out[4]
port 35 nsew signal output
rlabel metal2 s 10528 0 10640 800 6 io_out[5]
port 36 nsew signal output
rlabel metal2 s 12096 0 12208 800 6 io_out[6]
port 37 nsew signal output
rlabel metal2 s 13664 0 13776 800 6 io_out[7]
port 38 nsew signal output
rlabel metal2 s 15232 0 15344 800 6 io_out[8]
port 39 nsew signal output
rlabel metal2 s 16800 0 16912 800 6 io_out[9]
port 40 nsew signal output
rlabel metal2 s 17920 47200 18032 48000 6 rst_n
port 41 nsew signal input
rlabel metal4 s 4448 3076 4768 44748 6 vdd
port 42 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 44748 6 vdd
port 42 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 44748 6 vss
port 43 nsew ground bidirectional
rlabel metal2 s 6048 47200 6160 48000 6 wb_clk_i
port 44 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 48000 48000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2178192
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1-multi/openlane/wrapped_ay8913/runs/23_12_12_01_33/results/signoff/wrapped_ay8913.magic.gds
string GDS_START 270006
<< end >>

