* NGSPICE file created from wrapped_qcpu.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

.subckt wrapped_qcpu custom_settings[0] custom_settings[10] custom_settings[11] custom_settings[12]
+ custom_settings[13] custom_settings[14] custom_settings[15] custom_settings[16]
+ custom_settings[17] custom_settings[18] custom_settings[19] custom_settings[1] custom_settings[20]
+ custom_settings[21] custom_settings[22] custom_settings[23] custom_settings[24]
+ custom_settings[25] custom_settings[26] custom_settings[27] custom_settings[28]
+ custom_settings[29] custom_settings[2] custom_settings[30] custom_settings[31] custom_settings[3]
+ custom_settings[4] custom_settings[5] custom_settings[6] custom_settings[7] custom_settings[8]
+ custom_settings[9] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[32] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0]
+ io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17]
+ io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0]
+ io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17]
+ io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[24] io_out[25]
+ io_out[27] io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] rst_n sram_addr[0] sram_addr[1]
+ sram_addr[2] sram_addr[3] sram_addr[4] sram_addr[5] sram_gwe sram_in[0] sram_in[1]
+ sram_in[2] sram_in[3] sram_in[4] sram_in[5] sram_in[6] sram_in[7] sram_out[0] sram_out[1]
+ sram_out[2] sram_out[3] sram_out[4] sram_out[5] sram_out[6] sram_out[7] vdd vss
+ wb_clk_i io_oeb[22] io_out[26] io_out[23]
X_05903_ _01371_ _01375_ _01376_ _01377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_94_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09671_ _04671_ _04672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06337__A2 net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06883_ _02336_ _02346_ _02349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08622_ _03753_ _01872_ _03776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05834_ cpu.C _01308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05765_ cpu.uart.busy _01235_ _01239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08553_ _03713_ _03715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09287__A1 _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07504_ _02902_ _02704_ _02903_ _02904_ _01427_ cpu.uart.receive_div_counter\[1\]
+ _02905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_08484_ _03665_ _03666_ _00304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_81_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05696_ _01169_ _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07435_ _01542_ _02612_ _02842_ _02843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05631__I _01104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07366_ cpu.timer_top\[6\] _02781_ _02789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07297_ cpu.timer_capture\[2\] _02712_ _02731_ _02732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09105_ _02557_ _04143_ _04151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06317_ _01786_ _01691_ _01688_ _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__05076__A2 _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09036_ _01135_ _04093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06248_ _01715_ _01718_ _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_79_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06179_ _01648_ _01082_ _01649_ net53 _01432_ _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_13_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05459__S0 _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06025__A1 _01104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09938_ net82 _04894_ _04896_ _04891_ _04897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08389__I _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07293__I _02684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09869_ _04843_ _04844_ _04845_ _00510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_99_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output37_I net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_104_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09013__I _04065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07828__A2 _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10713_ net49 net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10644_ _00516_ clknet_leaf_74_wb_clk_i net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_101_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10575_ _00447_ clknet_leaf_81_wb_clk_i cpu.ROM_addr_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07468__I _00619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06567__A2 _01193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07516__A1 _00664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_60_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_60_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10009_ _02534_ _04763_ _04946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09269__A1 _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05550_ _00601_ _01024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_19_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07819__A2 _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05481_ cpu.base_address\[5\] _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_104_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08762__I _03875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07220_ _01924_ _02661_ _02667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_30_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07151_ _02401_ _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06102_ _01571_ _01572_ _01573_ _01574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_54_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07082_ _02535_ _02543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06270__A4 _01084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06033_ _01342_ _01505_ _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06007__A1 _01473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07755__A1 cpu.regs\[5\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07984_ _03266_ _03267_ _03268_ _03271_ _03272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_09723_ cpu.last_addr\[12\] cpu.last_addr\[11\] _04702_ _04723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06935_ cpu.PC\[4\] _02401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06866_ _02311_ _02330_ _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05369__I0 cpu.regs\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09654_ _04654_ _04630_ _04655_ _04656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_38_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05817_ _01287_ _01288_ _01290_ _01291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08605_ cpu.toggle_ctr\[3\] _03759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06797_ _02260_ _02261_ _02263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09585_ _04585_ _04586_ _04589_ _04590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05748_ net59 _01203_ _01209_ _01220_ _01221_ _01222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_08536_ _03152_ _03703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_38_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06457__I _01328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08467_ _03645_ _03653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05679_ _00005_ _01153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08398_ _03504_ _03598_ _00286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07418_ _02826_ _02827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07349_ _00926_ _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_70_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09432__A1 _02531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06246__A1 _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10042__A2 _04975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10360_ _00233_ clknet_leaf_49_wb_clk_i net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_103_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09019_ _02811_ _04073_ _04076_ _04078_ _00427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_10291_ _00164_ clknet_leaf_3_wb_clk_i cpu.regs\[5\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05964__C _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09499__A1 _02637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06721__A2 _00948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05204__C _00707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06485__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10627_ _00499_ clknet_leaf_70_wb_clk_i cpu.startup_cycle\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06237__A1 _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10558_ _00430_ clknet_leaf_55_wb_clk_i cpu.IO_addr_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10489_ _00362_ clknet_leaf_17_wb_clk_i cpu.pwm_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06720_ _02184_ _02185_ _02186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06651_ cpu.mem_cycle\[1\] _02117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07661__I _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05602_ _01032_ _01015_ _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06582_ cpu.timer_top\[15\] _01169_ _01176_ _02049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09370_ _02403_ _01120_ _04381_ _04382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08321_ _02778_ _03540_ _03541_ _03542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05533_ _01005_ _01006_ _01007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08252_ _02749_ _03487_ _00251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09662__B2 _04340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05464_ _00824_ _00940_ _00852_ _00941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07203_ cpu.PC\[7\] _02653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_7_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08183_ _02794_ _03431_ _00237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05395_ _00874_ _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_43_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07134_ _02586_ _02587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07065_ _02513_ _02527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_76_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05451__A2 _00903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06016_ _01488_ _01093_ _00987_ _01489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05356__I _00835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07967_ _03225_ _03250_ _03255_ _03201_ _03256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__06400__A1 _01337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09706_ cpu.last_addr\[9\] cpu.ROM_addr_buff\[9\] _04705_ _04706_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06918_ _02377_ _02378_ _02382_ _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_07898_ cpu.timer_div\[7\] _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10605__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07900__A1 cpu.timer_div\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09637_ _04362_ _04627_ _04640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06849_ _00763_ _02315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_87_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07900__B2 cpu.timer_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09568_ _00690_ _04441_ _04410_ _04574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08519_ cpu.orig_PC\[6\] _03684_ _03691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09499_ _02637_ _04445_ _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09653__A1 cpu.PC\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10412_ _00285_ clknet_leaf_36_wb_clk_i cpu.uart.receive_div_counter\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10343_ _00216_ clknet_leaf_63_wb_clk_i cpu.spi.data_out_buff\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05293__I2 cpu.regs\[10\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10274_ _00147_ clknet_leaf_4_wb_clk_i cpu.regs\[7\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_49_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10285__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08144__A1 _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08144__B2 _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_14_Left_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06458__A1 _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_104_Right_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_83_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05180_ _00001_ _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_23_Left_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06630__A1 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07656__I _02097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08870_ cpu.timer_capture\[11\] _03959_ _03964_ _03948_ _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_20_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05197__A1 _00003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07821_ cpu.PC\[8\] _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09092__B _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07752_ _03071_ _03076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07683_ _02975_ _03022_ _03028_ _00141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06703_ _02158_ _02168_ _02169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_32_Left_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09422_ _04374_ _04415_ _04432_ _04433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06634_ _01108_ _02100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_35_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09353_ _02848_ _04292_ _04365_ _04078_ _00474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06565_ _02031_ _01197_ _01198_ _02032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_4_5_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08304_ _03524_ _03526_ _03529_ _00261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05516_ _00668_ _00658_ _00990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_47_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09284_ _00983_ _01332_ cpu.base_address\[5\] _00931_ _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_7_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06496_ _01856_ _01960_ _01964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08235_ _03474_ _03475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05447_ _00924_ _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08166_ _03416_ _03417_ _03418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_43_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05378_ _00857_ _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07117_ _00619_ _02573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_41_Left_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08097_ cpu.uart.receive_buff\[2\] _03357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07048_ _02491_ _02500_ _02501_ _02509_ _02510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_100_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08999_ _02109_ _04062_ _04064_ _00421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08126__A1 _02893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07234__C _02666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_117_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_117_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_66_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10326_ _00199_ clknet_leaf_63_wb_clk_i cpu.spi.div_counter\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10257_ _00130_ clknet_leaf_4_wb_clk_i cpu.regs\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10188_ _00065_ clknet_leaf_19_wb_clk_i cpu.timer_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_109_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06983__C _02447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06555__I net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06350_ _01375_ _01815_ _01816_ _01819_ _01635_ _01820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_29_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06281_ cpu.uart.divisor\[12\] _01659_ _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05301_ _00799_ _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08020_ _03299_ _02871_ _03277_ _03300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_71_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06851__A1 _02315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05232_ _00686_ _00734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_114_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05163_ net18 _00611_ _00670_ _00671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09971_ cpu.PORTB_DDR\[4\] _04918_ _04920_ _04916_ _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05094_ _00603_ _00604_ _00605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_73_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05406__A2 _00874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08922_ _02694_ _04004_ _04005_ _04007_ _04008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_0_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08853_ _03943_ _03938_ _03950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08784_ _00613_ _03257_ _03858_ _03890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05996_ cpu.timer_top\[9\] _01170_ _01468_ _01469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07804_ cpu.regs\[3\]\[5\] _03099_ _03108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09156__I0 cpu.regs\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07735_ cpu.regs\[6\]\[3\] _03062_ _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_84_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09405_ _04343_ _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07666_ _03017_ _03019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_48_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07597_ _01735_ _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06617_ _01812_ _02083_ _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09336_ _04297_ _04349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_23_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06548_ _02015_ _02016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09267_ _00875_ _04240_ _04282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_51_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08218_ cpu.uart.div_counter\[4\] _03460_ _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_62_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06479_ _01936_ _01913_ _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_16_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09198_ cpu.last_addr\[7\] _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08149_ cpu.uart.div_counter\[6\] _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_95_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10111_ _03167_ _03278_ _05040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output67_I net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10042_ _04958_ _04975_ _04957_ _04964_ _04976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_101_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07322__A2 _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07858__B1 _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05884__A2 _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_85_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_85_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_53_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05212__C _00003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_14_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_14_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_112_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10309_ _00182_ clknet_leaf_15_wb_clk_i cpu.regs\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05495__S1 _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05850_ _01319_ _01175_ _01033_ _01323_ _01324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_89_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07561__A2 _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07520_ _00676_ _02920_ _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05781_ _01173_ _01254_ _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_99_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08765__I _02771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07451_ _00742_ _02857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06402_ cpu.toggle_top\[13\] _01871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07382_ _02795_ _02802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09121_ cpu.ROM_addr_buff\[3\] _04162_ _04155_ _04163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06333_ _01801_ _01802_ _01803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09052_ _02722_ _04105_ _04107_ _04108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06264_ _01734_ _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08003_ cpu.spi.div_counter\[2\] _03286_ _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_114_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06195_ cpu.uart.dout\[3\] _01192_ _01665_ _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05215_ _00718_ net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_25_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05146_ cpu.TIE cpu.needs_timer_interrupt cpu.needs_interrupt cpu.IE _00655_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_40_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09954_ _04906_ _04908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05077_ cpu.base_address\[0\] _00588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08905_ _02722_ _03987_ _03988_ _03993_ _03994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09885_ cpu.pwm_top\[5\] cpu.pwm_counter\[5\] _04857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08836_ cpu.timer_capture\[6\] _03930_ _03935_ _03924_ _03936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05979_ _01238_ _01448_ _01451_ _01452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08767_ cpu.timer_top\[9\] _03877_ _03880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_56_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08698_ cpu.pwm_counter\[4\] _03830_ _03832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_0_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07718_ _02015_ _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07649_ _02975_ _03004_ _03010_ _00125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_94_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10660_ _00532_ clknet_leaf_59_wb_clk_i net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_36_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07068__A1 _00609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09319_ _04329_ _04331_ _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10591_ _00463_ clknet_leaf_79_wb_clk_i cpu.last_addr\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_97_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08568__A1 _02695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput42 net42 io_oeb[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput64 net64 io_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput75 net75 io_out[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07240__A1 _02679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput53 net53 io_oeb[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput97 net97 sram_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput86 net86 sram_addr[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10025_ _04733_ _04960_ _04961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_106_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06806__A1 _00772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08559__A1 cpu.toggle_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06951_ _02122_ _02417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05902_ cpu.C _01357_ _01376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10090__I _05019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09670_ cpu.PC\[13\] _04670_ _04671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08621_ _03758_ _03774_ _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06882_ _02346_ _02347_ _02348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05184__I _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05833_ _01152_ _01166_ _01305_ _01306_ _01307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_EDGE_ROW_6_Left_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05764_ _00606_ _01179_ _01238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08552_ _03713_ _03714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07503_ cpu.uart.receive_div_counter\[6\] _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08483_ cpu.IO_addr_buff\[7\] _03659_ _03663_ _03666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05695_ _01075_ _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07434_ _02612_ _02841_ _02823_ _02842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07365_ _02787_ _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_73_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07296_ _02728_ _02715_ _02716_ _02730_ _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06316_ _01689_ _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09104_ _04150_ _00440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05076__A3 _00583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09035_ _02713_ _04086_ _04091_ _04092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06247_ _01716_ _01717_ _01718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06178_ _01215_ _01216_ _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_92_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07222__A1 _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05459__S1 _00935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06025__A2 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05129_ cpu.instr_buff\[15\] _00636_ cpu.base_address\[5\] _00637_ _00638_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_09937_ _02775_ _04895_ _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_5_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07574__I _02951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10109__A1 _01359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09868_ cpu.ROM_spi_cycle\[1\] _04840_ _04845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09799_ _04786_ _04784_ _04787_ _00498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08819_ _03231_ _03920_ _03921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05387__I1 cpu.regs\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07289__A1 _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10712_ net49 net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_83_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10643_ _00515_ clknet_leaf_19_wb_clk_i net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10574_ _00446_ clknet_leaf_85_wb_clk_i cpu.ROM_addr_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09450__A2 _01112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08801__C _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_79_Left_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10008_ _03432_ _04945_ _00549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08248__C _03479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09269__A2 _02705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05480_ _00956_ net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07150_ _02602_ _02603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_112_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06101_ cpu.timer_top\[2\] _01459_ _01264_ _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09441__A2 _04448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07081_ _02540_ _02542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05302__I1 _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06032_ _01364_ _01502_ _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08952__A1 _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07983_ cpu.spi.div_counter\[2\] _03269_ cpu.spi.div_counter\[4\] _03270_ _03271_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_09722_ _04704_ _04706_ _04707_ _04721_ _04722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_10_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06934_ cpu.PC\[6\] _02400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06865_ _02311_ _02330_ _02331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__05369__I1 _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09653_ cpu.PC\[11\] _00878_ _04655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_38_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05816_ _00646_ _01289_ _01290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08604_ cpu.toggle_ctr\[4\] _03756_ _03757_ cpu.toggle_ctr\[3\] _03758_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09584_ _04587_ _04562_ _04588_ _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_118_Right_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08535_ _03701_ _03693_ _03702_ _03695_ _00319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_54_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06796_ _02260_ _02261_ _02262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05747_ _00999_ _01221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08466_ cpu.orig_IO_addr_buff\[4\] _03648_ _03652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05678_ _01146_ _01052_ _01151_ _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_49_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09680__A2 _04671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08397_ _02904_ _03576_ _03597_ _03571_ _03598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_92_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07417_ _02631_ _02822_ _02826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_73_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07348_ _02773_ _02765_ _02774_ _02772_ _00060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_18_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06246__A2 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07279_ _02711_ _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09018_ _04077_ _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_60_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10290_ _00163_ clknet_leaf_3_wb_clk_i cpu.regs\[5\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09196__A1 cpu.ROM_addr_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08943__A1 cpu.spi.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05757__A1 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09024__I _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10626_ _00498_ clknet_leaf_70_wb_clk_i cpu.startup_cycle\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_70_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10557_ _00429_ clknet_leaf_31_wb_clk_i cpu.uart.divisor\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_114_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10488_ _00361_ clknet_leaf_17_wb_clk_i cpu.pwm_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_87_Left_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08103__I _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05748__A1 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_12_0_wb_clk_i clknet_0_wb_clk_i clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_75_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05890__C _01309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06558__I net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06650_ _02115_ _02116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_78_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05601_ _01040_ _01043_ _01048_ _01075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__05220__I0 cpu.regs\[4\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06581_ _02043_ _02045_ _02047_ _02048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_96_Left_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08320_ cpu.uart.data_buff\[6\] _03539_ _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05532_ cpu.IO_addr_buff\[4\] _00600_ _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08773__I _03875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08251_ _03399_ _03456_ _03486_ _03444_ _03487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05463_ cpu.regs\[4\]\[4\] cpu.regs\[5\]\[4\] cpu.regs\[6\]\[4\] cpu.regs\[7\]\[4\]
+ _00932_ _00935_ _00940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_07202_ _02593_ _02364_ _02651_ _02652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08182_ _03161_ _03418_ _03430_ _03417_ _03431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_70_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05394_ _00873_ _00874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07133_ _02107_ _02584_ _02585_ _02126_ _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__07425__A1 _01406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07064_ _02500_ _02522_ _02525_ _02526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06015_ _01487_ _01488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06242__B _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07728__A2 _03060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07966_ _03205_ _03254_ _03255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input29_I sram_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09705_ cpu.last_addr\[8\] _04700_ _04705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06917_ _02377_ _02378_ _02382_ _02383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07897_ cpu.timer_div_counter\[5\] _03186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09636_ _04626_ _04638_ _04436_ _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06468__I _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06164__B2 _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05372__I _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06848_ _02267_ _02313_ _02314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_87_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09567_ _04408_ _04315_ _04556_ _04573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06779_ _02214_ _02240_ _02243_ _02244_ _02245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_08518_ _03688_ _03690_ _00314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09498_ _04506_ _00478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09102__A1 _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08449_ _00623_ _00659_ _03638_ _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09653__A2 _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07299__I _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10411_ _00284_ clknet_leaf_35_wb_clk_i cpu.uart.receive_div_counter\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10342_ _00215_ clknet_leaf_61_wb_clk_i cpu.spi.data_out_buff\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output97_I net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05978__A1 cpu.spi.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05293__I3 cpu.regs\[11\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07719__A2 _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10273_ _00146_ clknet_leaf_2_wb_clk_i cpu.regs\[7\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_39_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_39_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_49_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06155__A1 _01132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06155__B2 _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05902__A1 cpu.C vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07655__A1 _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09638__B _04413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10609_ _00481_ clknet_leaf_96_wb_clk_i cpu.PC\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07820_ _03120_ _03121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__07672__I _03020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06394__A1 _01622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07751_ _03034_ _03073_ _03075_ _00162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06702_ _02165_ _02167_ _02168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07682_ cpu.regs\[8\]\[3\] _03025_ _03028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07894__A1 cpu.timer_div\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09421_ cpu.orig_PC\[3\] _04237_ _04432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06633_ _02019_ _02098_ _02099_ _00020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06564_ cpu.uart.divisor\[7\] _02031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09352_ _00625_ _04364_ _04321_ _04365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08303_ cpu.uart.data_buff\[0\] _03528_ _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07646__A1 cpu.regs\[10\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05515_ _00988_ _00989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_47_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09283_ _01331_ _01332_ _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06495_ _01865_ _01961_ _01948_ _01963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_7_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08234_ _03390_ _03469_ _03474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_51_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05446_ _00916_ _00923_ _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_28_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08165_ _03332_ _03417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05377_ _00856_ _00857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07116_ _00989_ _02568_ _02572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07847__I cpu.PC\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08096_ _03355_ _03352_ _03356_ _00226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_101_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07047_ _02111_ _02490_ _02508_ _00626_ _02509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_100_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09571__A1 _03696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08998_ _04063_ _04062_ _04064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07949_ cpu.timer_top\[3\] _03236_ _03237_ cpu.timer_top\[2\] _03238_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_46_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09619_ _03701_ _04554_ _04622_ _00483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_108_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10325_ _00198_ clknet_leaf_53_wb_clk_i cpu.needs_timer_interrupt vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10256_ _00129_ clknet_leaf_111_wb_clk_i cpu.regs\[10\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10187_ _00064_ clknet_leaf_20_wb_clk_i cpu.timer_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_89_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07628__A1 cpu.regs\[11\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06280_ _01749_ _01428_ _01659_ _01750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05300_ _00798_ _00799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05231_ _00711_ _00733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06851__A2 _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05162_ _00669_ _00670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09970_ _02778_ _04919_ _04920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05093_ cpu.IO_addr_buff\[2\] _00604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_73_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07800__A1 cpu.regs\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05257__I3 cpu.regs\[11\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05187__I _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08921_ cpu.timer\[12\] _04006_ _04007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08852_ _03949_ _00389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07803_ _01826_ _03101_ _03107_ _00182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08783_ _02815_ _03883_ _03889_ _03886_ _00380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05995_ _01177_ _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09156__I1 _02414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09305__A1 _04293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07734_ _03045_ _03059_ _03064_ _00156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07867__A1 _02531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07665_ _01736_ _03018_ _00133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09404_ _02860_ _04414_ _04415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06616_ _00818_ _01952_ _02083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_84_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07596_ _02973_ _02968_ _02974_ _00108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05650__I _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09335_ _04343_ _04331_ _04346_ _04347_ _04348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_23_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06547_ _01924_ _01926_ _01970_ _02014_ _02015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_09266_ cpu.orig_flags\[1\] _04272_ _04280_ _04281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_51_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06478_ net96 _01945_ _01946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08217_ _03457_ _03454_ _03460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05429_ _00906_ _00907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09197_ _04215_ _04219_ _04221_ _00462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_50_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08044__A1 _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08148_ _01661_ _03399_ _03400_ _02883_ _03401_ _03402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08079_ cpu.spi.data_in_buff\[4\] _03340_ _03342_ cpu.spi.data_in_buff\[5\] _03344_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08595__A2 _01413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05097__I _00607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10110_ _05039_ _00557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10041_ _04973_ _04974_ _04975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09544__A1 _04454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_6_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08092__B _00679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05192__S1 _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_54_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_54_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10308_ _00181_ clknet_leaf_14_wb_clk_i cpu.regs\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__06597__A1 _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_60_Left_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09535__A1 _04529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06349__A1 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10239_ _00112_ clknet_leaf_113_wb_clk_i cpu.regs\[12\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05780_ _01174_ _01180_ _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_88_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07450_ _02845_ _02854_ _02856_ _00080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07381_ _02795_ _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06401_ net31 _01096_ _01869_ _01403_ _01870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__08274__A1 _01423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09120_ _00743_ _02861_ _04153_ _04162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_57_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06332_ net93 _00924_ _01802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09051_ cpu.orig_IO_addr_buff\[1\] _04106_ _04107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10081__A1 _01359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08002_ cpu.spi.div_counter\[2\] _03286_ _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06263_ _01686_ _01732_ _01733_ _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06194_ _01664_ _01665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05214_ _00717_ _00718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05145_ _00625_ _00653_ _00654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09953_ _04906_ _04907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05076_ _00572_ _00576_ _00583_ _00586_ _00587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_110_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08904_ cpu.timer\[9\] _03989_ _03993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09884_ cpu.pwm_top\[0\] _03826_ cpu.pwm_counter\[1\] _04854_ _04855_ _04856_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08835_ _03227_ _03918_ _03894_ _03934_ _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08766_ _02671_ _03876_ _03878_ _03879_ _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_input11_I io_in[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05978_ cpu.spi.divisor\[1\] _01238_ _01450_ _01451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_56_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07717_ _03051_ _03040_ _03052_ _00151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_67_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08697_ _03830_ _03831_ _00352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_0_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06512__A1 cpu.uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07648_ cpu.regs\[10\]\[3\] _03007_ _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07579_ cpu.regs\[13\]\[6\] _02959_ _02962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_36_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09318_ _04330_ _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10590_ _00462_ clknet_leaf_80_wb_clk_i cpu.last_addr\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_97_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05618__A3 _01074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09249_ _04259_ _04262_ _04263_ _04264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_106_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput43 net43 io_oeb[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_31_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput54 net54 io_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput76 net76 io_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput65 net65 io_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_101_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09517__A1 _04413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput87 net87 sram_addr[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10024_ _02581_ _02112_ _02487_ _04960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_106_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_101_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_101_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_86_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07945__I cpu.timer_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06950_ _02125_ _02415_ _02416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input3_I io_in[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05901_ _01374_ _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06881_ _02321_ _00857_ _02347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05832_ _01052_ _01055_ _01151_ _01306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_08620_ _03767_ _03773_ _03761_ _03774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08776__I _02771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05763_ _01192_ _01233_ _01235_ _01236_ _01237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_08551_ _01415_ _03712_ _03713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07502_ cpu.uart.divisor\[6\] _02903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_77_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08482_ cpu.orig_IO_addr_buff\[7\] _03655_ _03665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05694_ _01009_ _01168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05414__B _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07433_ _02838_ _02429_ _02615_ _02840_ _02841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_33_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07364_ _01915_ _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_84_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09103_ _00881_ _04142_ _04149_ _04145_ _04150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_45_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07295_ _02729_ _02718_ _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06315_ _01783_ _01784_ _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_5_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05076__A4 _00586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09034_ cpu.orig_IO_addr_buff\[0\] _04090_ _04091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06246_ _01600_ net92 _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_107_Left_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_103_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06177_ net82 _01648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07222__A2 _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05128_ cpu.base_address\[4\] _00637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_110_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09936_ _04886_ _04895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_86_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05059_ cpu.br_rel_dest\[7\] _00570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_5_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09867_ cpu.ROM_spi_cycle\[1\] _04840_ _04844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09798_ _04786_ _04784_ _03912_ _04787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_116_Left_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08818_ _03236_ _03914_ _03920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__05387__I2 cpu.regs\[2\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08749_ _03863_ _03866_ _03867_ _00368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_95_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08486__A1 _01310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_95_Right_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10642_ _00514_ clknet_leaf_63_wb_clk_i net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_101_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10573_ _00445_ clknet_leaf_81_wb_clk_i cpu.ROM_addr_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_63_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06972__A1 _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10007_ cpu.ROM_spi_mode _04944_ _04945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09910__A1 _03849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08545__B _03709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10036__A1 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09977__A1 cpu.PORTB_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06100_ cpu.timer_capture\[10\] _01460_ _01464_ _01572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07080_ _02540_ _02541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05302__I2 cpu.regs\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06031_ _01503_ _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_23_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07452__A2 _01732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07982_ cpu.spi.divisor\[4\] _03270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_09721_ _04708_ _04709_ _04718_ _04720_ _04721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__06963__A1 cpu.PC\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06933_ cpu.PC\[8\] _02399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05518__A2 cpu.br_rel_dest\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09652_ cpu.PC\[11\] _00878_ _04654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06864_ _02318_ _02328_ _02329_ _02330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_38_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05815_ _01062_ _01289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08603_ cpu.toggle_top\[3\] _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06795_ _02230_ _02228_ _02261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09583_ cpu.PC\[8\] _00821_ _04588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05746_ _01212_ _01214_ _01218_ _01219_ net39 _01220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_77_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08534_ cpu.orig_PC\[10\] _03641_ _03702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08468__A1 _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08465_ _03641_ _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05677_ _01147_ _01150_ _01151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08396_ _02904_ _03596_ _03597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_107_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07691__A2 _03032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07416_ _02821_ _02824_ _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07347_ cpu.timer_top\[2\] _02766_ _02774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09017_ _02531_ _04077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07278_ _02714_ _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06229_ _01687_ _01699_ _01700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05757__A2 _01229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09919_ _02698_ _04879_ _04883_ _04882_ _00522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_output42_I net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06182__A2 _01203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10625_ _00497_ clknet_leaf_70_wb_clk_i cpu.startup_cycle\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09959__A1 cpu.PORTB_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10556_ _00428_ clknet_leaf_31_wb_clk_i cpu.uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_114_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10487_ _00360_ clknet_leaf_18_wb_clk_i cpu.pwm_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05748__A2 _01203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06945__A1 cpu.PC\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08147__B1 _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05600_ _00606_ _01073_ _01074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_59_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06173__A2 _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05220__I1 cpu.regs\[5\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06580_ _02046_ _01258_ _01075_ _02047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_24_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05920__A2 _01380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05531_ _00603_ _00604_ _01005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_74_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07122__A1 _01591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08250_ _03399_ _03485_ _03486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08870__A1 cpu.timer_capture\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05462_ _00913_ _00938_ _00939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08181_ _03161_ _03429_ _03430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10009__A1 _02534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06507__C _01225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer1_I _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07201_ _02331_ _02362_ _02363_ _02651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_9_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_9_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_55_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05393_ _00872_ _00873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07132_ _01109_ _02103_ _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_113_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07063_ cpu.ROM_addr_buff\[3\] _02523_ _02524_ cpu.ROM_addr_buff\[7\] _02498_ _02525_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__07976__A3 _01424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05918__I _01380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06014_ cpu.br_rel_dest\[1\] _01487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_07965_ _03214_ _03253_ _03254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09704_ cpu.ROM_addr_buff\[11\] _04703_ _04704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06916_ _02379_ _02381_ _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07896_ cpu.timer_div_counter\[1\] _03185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_69_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09350__A2 _04362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09635_ _04633_ _04637_ _04341_ _04638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07361__A1 cpu.timer_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10211__D _00084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06847_ _00689_ _00900_ _02313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09566_ _04368_ _04556_ _04571_ _04400_ _04572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06778_ _00761_ net116 _02244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05729_ _01202_ _01203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08517_ _02622_ _03686_ _03689_ _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09497_ _02622_ _04445_ _04505_ _04476_ _04506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07113__A1 _01105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08448_ _03637_ _00628_ _03638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08861__A1 _03259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10410_ _00283_ clknet_leaf_36_wb_clk_i cpu.uart.receive_div_counter\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08379_ _02877_ _03581_ _03582_ _03583_ _03584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_92_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10341_ _00214_ clknet_leaf_62_wb_clk_i cpu.spi.data_out_buff\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08204__I _02809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10272_ _00145_ clknet_leaf_110_wb_clk_i cpu.regs\[8\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_79_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_79_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_79_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07352__A1 _02776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08095__B _00679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10608_ _00480_ clknet_leaf_91_wb_clk_i cpu.PC\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10539_ _00412_ clknet_leaf_48_wb_clk_i cpu.spi.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05418__A1 _00825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07750_ cpu.regs\[5\]\[0\] _03074_ _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06701_ _02136_ _02166_ _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07681_ _02973_ _03022_ _03027_ _00140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09420_ _04421_ _04424_ _04430_ _04394_ _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06632_ cpu.regs\[9\]\[7\] _02019_ _02099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06563_ _02027_ _02028_ _02029_ _02030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09351_ _04324_ _04360_ _04363_ _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08302_ _03527_ _03528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05514_ cpu.br_rel_dest\[1\] _00988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09282_ _04295_ _04296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08233_ _03403_ _03470_ _03468_ _03473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08843__A1 cpu.timer_capture\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06494_ _01865_ _01959_ _01961_ _01962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_35_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05445_ _00920_ _00922_ _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08164_ _03262_ _03415_ _03416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_7_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05376_ _00855_ _00856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08095_ cpu.uart.dout\[1\] _03353_ _00679_ _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07115_ _02549_ _02571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_15_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08071__A2 _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07046_ _02503_ _02507_ _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__06082__A1 _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_113_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09020__A1 cpu.uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09571__A2 _04554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08997_ _03637_ _04063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07582__A1 _02098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07948_ _02729_ _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07879_ cpu.spi.dout\[3\] _03165_ _03169_ cpu.spi.data_in_buff\[3\] _03173_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07334__A1 _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09618_ _04367_ _04618_ _04621_ _04622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09549_ _03122_ _04531_ _04555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07103__I _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08598__B1 _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10324_ _00197_ clknet_leaf_44_wb_clk_i cpu.spi.dout\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09011__A1 _02690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10255_ _00128_ clknet_leaf_117_wb_clk_i cpu.regs\[10\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10186_ _00063_ clknet_leaf_20_wb_clk_i cpu.timer_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_109_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09078__A1 _02745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05230_ _00694_ _00732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05161_ _00668_ _00669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09250__A1 _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05092_ cpu.IO_addr_buff\[3\] _00603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_40_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08920_ _01254_ _04006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08851_ cpu.timer_capture\[8\] _03930_ _03946_ _03948_ _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07802_ cpu.regs\[3\]\[4\] _03103_ _03107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06367__A2 _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05994_ _01458_ _01462_ _01466_ _01467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08782_ cpu.timer_top\[15\] _03884_ _03889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07733_ cpu.regs\[6\]\[2\] _03062_ _03064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_79_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07664_ _01644_ _03018_ _00132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_84_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09403_ _02403_ _02837_ _02829_ _04414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_1_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06615_ _00818_ _02081_ _02082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07595_ cpu.regs\[12\]\[2\] _02969_ _02974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06546_ _01314_ _01587_ _02011_ _02013_ _02014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_09334_ _04296_ _04347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_23_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09265_ _04275_ _04277_ _04278_ _04279_ _04280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_7_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06477_ net95 _01850_ _01945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08216_ _02749_ _03459_ _00243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09196_ cpu.ROM_addr_buff\[6\] _04220_ _04221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05428_ _00905_ _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_105_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08147_ _03390_ _02704_ _01658_ cpu.uart.div_counter\[3\] _03401_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__07079__B _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05359_ _00826_ _00838_ _00839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_113_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08078_ _03343_ _00221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05489__S0 _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07029_ _02486_ _02490_ _02491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__05802__A1 _01275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10040_ cpu.ROM_addr_buff\[2\] _02494_ _02523_ cpu.ROM_addr_buff\[6\] _02495_ _04974_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__06358__A2 _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06937__I cpu.PC\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05413__S0 _00829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07858__A2 _02412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09188__C _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09983__I _04928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09232__A1 _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07794__A1 _01406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06597__A2 _01164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10307_ _00180_ clknet_leaf_13_wb_clk_i cpu.regs\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xclkbuf_leaf_94_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_94_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10238_ _00111_ clknet_leaf_113_wb_clk_i cpu.regs\[12\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10169_ _00046_ clknet_leaf_22_wb_clk_i cpu.uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xclkbuf_leaf_23_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_23_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05237__B _00707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06400_ _01337_ _01833_ _01849_ _01868_ _01869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_07380_ _02768_ _02800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06331_ _01704_ _01712_ _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09050_ _04089_ _04106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09471__A1 _02401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06262_ net29 _01334_ _01733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08001_ _03279_ _03287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05213_ _00708_ _00716_ _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_06193_ _01234_ _01243_ _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10037__C _03421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05144_ _00629_ _00652_ _00653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09952_ _01741_ _04036_ _04906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05075_ _00584_ _00585_ _00586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08730__C _03853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08903_ _03992_ _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10053__B _04731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09883_ cpu.pwm_top\[4\] cpu.pwm_counter\[4\] _04855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_0_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08834_ _03932_ _03933_ _03934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08765_ _02771_ _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05977_ _01449_ _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_56_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07716_ cpu.regs\[7\]\[5\] _03038_ _03052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08696_ cpu.pwm_counter\[3\] _03829_ _03709_ _03831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_0_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07647_ _02973_ _03004_ _03009_ _00124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_94_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07578_ _01922_ _02958_ _02961_ _00103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_36_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06529_ _01994_ _01995_ _01996_ _01997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09317_ _02837_ _02829_ _04330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_118_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06276__A1 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07588__I _02967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09248_ _01638_ _01518_ _02124_ _04263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09179_ cpu.last_addr\[2\] _04199_ _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput66 net66 io_out[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput55 net55 io_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_output72_I net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput44 net44 io_oeb[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05836__I _01309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput77 net77 io_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_101_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08212__I _03440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput88 net88 sram_addr[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09517__A2 _04315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10023_ cpu.ROM_addr_buff\[0\] _02494_ _02495_ _04959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_106_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06019__A1 _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09508__A2 _01119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05900_ _01372_ _01373_ _01374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06880_ _02345_ _00871_ _02346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05831_ _01292_ _01298_ _01304_ _01305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_118_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05762_ cpu.uart.dout\[0\] _01192_ _01236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08550_ _02673_ _03712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07501_ cpu.uart.receive_div_counter\[7\] _02902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08481_ _03661_ _03664_ _00303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05693_ cpu.toggle_top\[0\] _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_49_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07432_ _02596_ _02348_ _02839_ _02840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_85_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07363_ _02784_ _02780_ _02785_ _02786_ _00063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_61_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09102_ _02552_ _04143_ _04149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07294_ cpu.timer\[2\] _02729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06314_ _00768_ _00961_ _01784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09033_ _04089_ _04090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06245_ _01617_ _01620_ _01716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06176_ _01421_ _01647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05127_ cpu.instr_buff\[14\] _00636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_92_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09935_ _04886_ _04894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05058_ _00567_ _00568_ _00569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_5_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09866_ _03181_ _04842_ _04843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08183__A1 _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08817_ _03890_ _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09797_ cpu.startup_cycle\[5\] _04786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_99_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05387__I3 cpu.regs\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08748_ cpu.timer_div_counter\[3\] _03864_ _03867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_67_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08679_ _03795_ _03818_ _03819_ _00346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_95_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10641_ _00513_ clknet_leaf_65_wb_clk_i cpu.ROM_spi_cycle\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_101_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06249__A1 _01132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10572_ _00444_ clknet_leaf_81_wb_clk_i cpu.ROM_addr_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07111__I _02567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06249__B2 _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05566__I _01039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08174__A1 _03421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10006_ _04793_ _00582_ _04943_ _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_86_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08477__A2 _03655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06488__A1 _01622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09426__A1 _04362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_30_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05302__I3 cpu.regs\[3\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06030_ _01364_ _01502_ _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06660__A1 _02123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07452__A3 _01733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07981_ cpu.spi.divisor\[2\] _03269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_09720_ cpu.last_addr\[6\] cpu.ROM_addr_buff\[6\] _04719_ _04720_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_06932_ cpu.PC\[12\] _02398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09901__A2 _03712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07912__A1 cpu.timer_top\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09651_ _04498_ _04649_ _04652_ _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06863_ _02326_ _02327_ _02329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_38_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05814_ _01283_ _01288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08602_ cpu.toggle_top\[4\] _03756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06794_ _02252_ _02258_ _02259_ _02260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__05369__I3 cpu.regs\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09582_ cpu.PC\[8\] _00588_ _04587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05745_ _01030_ _01032_ _01042_ _01215_ _01219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_08533_ _03700_ _03701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_65_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05676_ _00618_ _01149_ _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08464_ _00603_ _03642_ _03650_ _03646_ _00300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_08395_ _02881_ _03590_ _03596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07415_ _02823_ _02824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07346_ _02685_ _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10209__D _00082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09016_ cpu.uart.divisor\[13\] _04074_ _04076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07277_ _01181_ _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06228_ _01692_ _01698_ _01347_ _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06159_ _01509_ _01613_ _01630_ _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_09918_ net64 _04880_ _04883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_69_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09849_ cpu.ROM_spi_dat_out\[4\] _04831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07903__A1 cpu.timer_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06706__A2 _00973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06167__B1 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07903__B2 cpu.timer_div\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output35_I net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09408__A1 cpu.PC\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10624_ _00496_ clknet_leaf_68_wb_clk_i cpu.startup_cycle\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10555_ _00427_ clknet_leaf_31_wb_clk_i cpu.uart.divisor\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10486_ _00359_ clknet_leaf_18_wb_clk_i cpu.pwm_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_114_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_14_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05530_ _01003_ _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_47_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07122__A2 _02567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06855__I _00689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05461_ cpu.regs\[0\]\[4\] cpu.regs\[1\]\[4\] cpu.regs\[2\]\[4\] cpu.regs\[3\]\[4\]
+ _00932_ _00935_ _00938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_117_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08180_ _03425_ _03428_ _03429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_55_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05392_ _00871_ _00872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07200_ _02630_ _02649_ _02650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07131_ _02109_ _02583_ _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_54_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08622__A2 _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07062_ _02501_ _02524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06013_ _01484_ _01312_ _01485_ _01486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_103_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07964_ _03221_ _03252_ _03211_ _03253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05934__I _01141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09703_ cpu.last_addr\[11\] _04702_ _04703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07895_ cpu.timer_div\[3\] cpu.timer_div_counter\[3\] _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06915_ _02376_ _02380_ _02381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09634_ _01126_ _04388_ _04636_ _04394_ _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06846_ _00741_ _00870_ _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09565_ _04373_ _04559_ _04570_ _04397_ _04571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06777_ _02242_ _02241_ _02243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05728_ _01038_ _01201_ _01202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08516_ _03662_ _03689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09496_ _04478_ _04482_ _04484_ _04453_ _04504_ _04505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08447_ _00584_ _03637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05659_ cpu.instr_buff\[14\] _01133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_93_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08980__I _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06872__A1 _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08378_ _03570_ _03583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07329_ cpu.timer_capture\[7\] _02738_ _02758_ _02759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08613__A2 cpu.toggle_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10340_ _00213_ clknet_leaf_65_wb_clk_i cpu.spi.data_out_buff\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10271_ _00144_ clknet_leaf_117_wb_clk_i cpu.regs\[8\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09316__I _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_48_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_48_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_83_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05210__S1 _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10607_ _00479_ clknet_leaf_91_wb_clk_i cpu.PC\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10538_ _00411_ clknet_leaf_48_wb_clk_i cpu.spi.divisor\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10469_ _00342_ clknet_leaf_5_wb_clk_i cpu.toggle_ctr\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_48_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06700_ _00805_ _00950_ _02166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08540__A1 _02414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07680_ cpu.regs\[8\]\[2\] _03025_ _03027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06631_ _02097_ _02098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_35_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06562_ net14 _01072_ _01196_ _02029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_86_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09350_ _04324_ _04362_ _04331_ _04363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08301_ _03408_ _03413_ _03520_ _03527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09281_ _01332_ _04294_ _04295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05513_ _00986_ _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_117_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08232_ _03471_ _03472_ _00246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06493_ _01960_ _01961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05444_ _00913_ _00921_ _00852_ _00922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_28_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08163_ _00623_ _01424_ _03310_ _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_43_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05375_ _00839_ _00848_ _00850_ _00854_ _00855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_27_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08094_ cpu.uart.receive_buff\[1\] _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07114_ _02560_ _02569_ _02570_ _02533_ _00030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07045_ _02504_ _02506_ _02479_ _02507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_3_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08359__A1 _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08996_ _04061_ _04062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_89_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09159__I0 cpu.regs\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07947_ cpu.timer\[3\] _03236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07878_ _03172_ _00192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_97_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09617_ _04402_ _04605_ _04620_ _04439_ _02624_ _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_06829_ _02268_ _02292_ _02293_ _02294_ _02295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_09548_ _03181_ _04243_ _04554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_65_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09479_ _04486_ _04487_ _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_65_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10323_ _00196_ clknet_leaf_42_wb_clk_i cpu.spi.dout\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06073__A2 _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10254_ _00127_ clknet_leaf_118_wb_clk_i cpu.regs\[10\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10185_ _00062_ clknet_leaf_20_wb_clk_i cpu.timer_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08770__A1 _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07089__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05160_ net71 _00668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05091_ _00598_ _00601_ _00602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08850_ _03947_ _03948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08761__A1 _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07801_ _01735_ _03100_ _03106_ _00181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05993_ _01463_ _01464_ _01465_ _01466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08781_ _02788_ _03883_ _03888_ _03886_ _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_79_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08513__A1 _02605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07732_ _03042_ _03059_ _03063_ _00155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08728__C _03853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07663_ _01543_ _03018_ _00131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09402_ _04407_ _04413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06614_ net95 _00804_ _01850_ _02081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09333_ _04342_ _04345_ _04346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07594_ _01643_ _02973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06545_ _02012_ _01152_ _02013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_23_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06476_ _01834_ _01942_ _01943_ _01944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__05186__S0 _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09264_ _01316_ _02820_ _02345_ _01488_ _04279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_118_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09195_ _04202_ _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08215_ cpu.uart.div_counter\[3\] _03456_ _03458_ _03444_ _03459_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_63_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05427_ cpu.base_address\[3\] _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08146_ cpu.uart.div_counter\[9\] _03400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05358_ cpu.regs\[12\]\[0\] cpu.regs\[13\]\[0\] cpu.regs\[14\]\[0\] cpu.regs\[15\]\[0\]
+ _00832_ _00837_ _00838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_31_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08077_ cpu.spi.data_in_buff\[3\] _03340_ _03342_ cpu.spi.data_in_buff\[4\] _03343_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_101_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05489__S1 _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05289_ _00774_ _00788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07028_ _02487_ _02489_ _02490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__05802__A2 _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07555__A2 _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05394__I _00873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08979_ _03180_ _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_98_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05318__A1 _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05413__S1 _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07858__A3 _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07243__A1 _02685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06046__A2 _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10306_ _00179_ clknet_leaf_14_wb_clk_i cpu.regs\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_72_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10237_ _00110_ clknet_leaf_113_wb_clk_i cpu.regs\[12\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10168_ _00045_ clknet_leaf_40_wb_clk_i cpu.uart.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10099_ _00817_ _02081_ _05029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_63_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_63_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_88_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06330_ _01387_ _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_29_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06261_ _00982_ _01731_ _01732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08000_ _03280_ _03285_ _03286_ _00200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_72_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05212_ _00699_ _00713_ _00715_ _00003_ _00716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_06192_ _01657_ _01660_ _01662_ _01663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07234__A1 _02671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05143_ cpu.uart.busy cpu.spi.busy _00651_ _00652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_13_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09951_ _04905_ _00532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05074_ cpu.instr_cycle\[2\] _00585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08902_ cpu.timer_capture\[8\] _03986_ _03991_ _03979_ _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_57_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09882_ cpu.pwm_top\[1\] _04854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09842__C _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08833_ _02751_ _03931_ _03890_ _03933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05976_ _00606_ _01174_ _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08764_ cpu.timer_top\[8\] _03877_ _03878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_56_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07715_ _01920_ _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08695_ cpu.pwm_counter\[3\] _03829_ _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07646_ cpu.regs\[10\]\[2\] _03007_ _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07577_ cpu.regs\[13\]\[5\] _02959_ _02961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_36_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06528_ cpu.pwm_top\[6\] _01268_ _01270_ _01996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09316_ _04327_ _04329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06276__A2 _01221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09247_ _01529_ _04255_ _04261_ _04262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_97_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06459_ _01904_ _01906_ _01909_ _01911_ _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_105_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09178_ _04193_ _04205_ _04207_ _00457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_90_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08129_ cpu.uart.div_counter\[0\] _03383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08973__A1 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput34 net34 io_oeb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_31_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput67 net67 io_out[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput56 net56 io_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput45 net45 io_oeb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput78 net78 io_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_output65_I net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput89 net89 sram_gwe vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08725__A1 _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10022_ _04763_ _04958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06200__A2 _01669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06948__I _02398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_113_Right_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07700__A2 _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09994__I _04928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_110_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_110_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_117_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06019__A2 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_9_0_wb_clk_i clknet_0_wb_clk_i clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07519__A2 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08192__A2 _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05830_ _01300_ _01303_ _01304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09234__I _03503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07500_ _02885_ cpu.uart.receive_div_counter\[15\] _02899_ cpu.uart.divisor\[3\]
+ _02900_ _02901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05761_ _01234_ _01235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09141__A1 _03696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08480_ cpu.IO_addr_buff\[6\] _03659_ _03663_ _03664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05692_ _01165_ _01166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07431_ _02345_ _00979_ _00875_ _02820_ _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_91_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07362_ _02771_ _02786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_33_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06313_ _01782_ _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09101_ _04148_ _00439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_84_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07293_ _02684_ _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_45_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09032_ _04088_ _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_60_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06244_ _01695_ _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06175_ _01113_ _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06542__B _02009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05126_ _00633_ _00634_ _00635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_92_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05769__A1 _01186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09934_ _02773_ _04887_ _04893_ _00527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05057_ cpu.IO_addr_buff\[0\] _00568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09865_ cpu.ROM_spi_cycle\[4\] _00578_ _04840_ _04842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_clkbuf_leaf_59_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08816_ _03907_ _03918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09796_ _04779_ _04780_ _04784_ _04785_ _00497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05959_ _01003_ _01210_ _01432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08747_ cpu.timer_div_counter\[3\] _03864_ _03866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_95_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08678_ cpu.toggle_ctr\[13\] _03816_ _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_67_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07629_ _02977_ _02991_ _02997_ _00118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10640_ _00512_ clknet_leaf_65_wb_clk_i cpu.ROM_spi_cycle\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10571_ _00443_ clknet_leaf_80_wb_clk_i cpu.ROM_addr_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_98_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08946__A1 _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_2_Left_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_39_Left_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_112_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10005_ _02480_ _04786_ _02475_ _04943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_99_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_48_Left_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09674__A2 _04671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07685__A1 _02977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09426__A2 _04415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07988__A2 cpu.spi.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_57_Left_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05999__A1 _01413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07980_ cpu.spi.div_counter\[0\] cpu.spi.divisor\[0\] _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06931_ _02135_ _02395_ _02396_ _02397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09650_ cpu.orig_PC\[12\] _04088_ _04652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_66_Left_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08601_ _03753_ cpu.toggle_top\[5\] cpu.toggle_top\[4\] _03754_ _03755_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06862_ _02326_ _02327_ _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05813_ _00984_ _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06793_ _02254_ _02255_ _02257_ _02259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_09581_ cpu.PC\[9\] _00882_ _04586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_38_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05744_ _01215_ _01217_ cpu.PORTA_DDR\[0\] _01218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08532_ cpu.PC\[10\] _03700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08463_ cpu.orig_IO_addr_buff\[3\] _03648_ _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06479__A2 _01913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07676__A1 _02964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05675_ _00585_ _01148_ _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07414_ _02126_ _02585_ _02822_ _02823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08394_ _02881_ _03590_ _03595_ _03585_ _00285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_107_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07345_ _02769_ _02765_ _02770_ _02772_ _00059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07428__A1 _02340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_75_Left_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_72_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06100__A1 cpu.timer_capture\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07276_ _02669_ _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_61_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09015_ _04047_ _04073_ _04075_ _04070_ _00426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_61_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06227_ _01695_ _01697_ _01698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_115_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07087__C _02547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06158_ net91 _01513_ _01630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06089_ _01440_ _01558_ _01559_ _01560_ _01561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05109_ _00618_ _00619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09917_ _04047_ _04879_ _04881_ _04882_ _00521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09353__A1 _02848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09848_ _04830_ _00504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06167__B2 _01638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09779_ _02513_ _04770_ _04771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__09105__A1 _02557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10623_ _00495_ clknet_leaf_68_wb_clk_i cpu.startup_cycle\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08616__B1 _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10554_ _00426_ clknet_leaf_31_wb_clk_i cpu.uart.divisor\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05577__I _00991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10485_ _00358_ clknet_leaf_102_wb_clk_i cpu.pwm_top\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_114_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09592__A1 _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06158__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05460_ _00841_ _00936_ _00846_ _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_15_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08607__B1 cpu.toggle_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05391_ _00870_ _00871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07130_ _02116_ _02580_ _02582_ _02583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_82_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07061_ _02491_ _02523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06633__A2 _02098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06012_ _01313_ _01485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07963_ _03223_ _03251_ _03220_ _03252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09702_ _04228_ _04701_ _04702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07894_ cpu.timer_div\[4\] cpu.timer_div_counter\[4\] _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06914_ _00800_ _01929_ _02380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09633_ _03152_ _04634_ _04425_ _04635_ _04636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06845_ _02305_ _02306_ _02301_ _02311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_09564_ _04566_ _04569_ _04570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08515_ cpu.orig_PC\[5\] _03684_ _03688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06776_ _00724_ _00943_ _02242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05727_ _01032_ _01015_ _01201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09495_ _04454_ _04503_ _04504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08446_ _02873_ _00616_ _03636_ _00296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05658_ _01131_ _01132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_37_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08377_ _02877_ cpu.uart.receive_div_counter\[1\] cpu.uart.receive_div_counter\[0\]
+ _03582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XPHY_EDGE_ROW_83_Left_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07328_ _02739_ _02755_ _02740_ _02757_ _02758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05589_ _01061_ _01062_ _01063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_61_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07259_ _02698_ _02691_ _02699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05397__I _00876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10270_ _00143_ clknet_leaf_118_wb_clk_i cpu.regs\[8\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_92_Left_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06388__A1 _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07117__I _00619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06312__A1 _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_88_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_88_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10606_ _00478_ clknet_leaf_91_wb_clk_i cpu.PC\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10537_ _00410_ clknet_leaf_47_wb_clk_i cpu.spi.divisor\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_17_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_17_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_101_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10468_ _00341_ clknet_leaf_6_wb_clk_i cpu.toggle_ctr\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_75_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10399_ _00272_ clknet_leaf_44_wb_clk_i cpu.uart.receive_buff\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08411__I _03503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06630_ net33 _00985_ _02062_ _02096_ _02097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_35_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05770__I _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06551__A1 _01408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06561_ net5 _01436_ _01745_ _02028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08286__C _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08300_ _03525_ _03526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09280_ _01095_ _00957_ _04294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06492_ _01833_ _00976_ _01960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05512_ _00982_ _00985_ _00986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_08231_ _03403_ _03468_ _03464_ _03472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05443_ cpu.regs\[0\]\[3\] cpu.regs\[1\]\[3\] cpu.regs\[2\]\[3\] cpu.regs\[3\]\[3\]
+ _00828_ _00910_ _00921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_83_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08162_ _03373_ _03409_ _00239_ _03414_ _00233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_43_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05374_ _00826_ _00851_ _00853_ _00854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08093_ _03347_ _03352_ _03354_ _00225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07803__A1 _01826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07113_ _01105_ _02568_ _02570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07044_ _02505_ _02506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09556__A1 _04529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05945__I _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05417__I0 cpu.regs\[4\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08995_ _04060_ _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09159__I1 _03708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07946_ _03233_ _02734_ cpu.timer\[4\] _03234_ _03235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input27_I sram_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07877_ cpu.spi.dout\[2\] _03165_ _03169_ cpu.spi.data_in_buff\[2\] _03172_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09616_ _00727_ _04450_ _04619_ _04620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06828_ _00710_ _00949_ _00944_ _00688_ _02294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09547_ _04553_ _00480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06759_ _02222_ _02224_ _02225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_26_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09478_ cpu.PC\[4\] cpu.br_rel_dest\[4\] _04461_ _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08429_ _03609_ _03623_ _00292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_108_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_11_0_wb_clk_i clknet_0_wb_clk_i clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_19_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10322_ _00195_ clknet_leaf_47_wb_clk_i cpu.spi.dout\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output95_I net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09755__C _00666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05281__A1 _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10253_ _00126_ clknet_leaf_119_wb_clk_i cpu.regs\[10\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10184_ _00061_ clknet_leaf_20_wb_clk_i cpu.timer_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_70_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06533__A1 _00663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09997__I _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07089__A2 _02543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10093__A1 _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05195__S1 _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08406__I cpu.uart.receive_div_counter\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08038__A1 _02760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09786__A1 _04771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05090_ _00599_ _00600_ _00601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09538__A1 _04529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08780_ cpu.timer_top\[14\] _03884_ _03888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07800_ cpu.regs\[3\]\[3\] _03103_ _03106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05992_ _01169_ _01465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07731_ cpu.regs\[6\]\[1\] _03062_ _03063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07662_ _01407_ _03018_ _00130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09401_ _04366_ _04412_ _00475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06613_ _02076_ _02079_ _02080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07593_ _02971_ _02968_ _02972_ _00107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_75_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06544_ _01773_ _02012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09332_ _02847_ _01488_ _04344_ _04345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_48_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06475_ _01848_ _01941_ _01943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09263_ _01600_ _02855_ _00742_ _01806_ _04278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_08214_ _03457_ _03454_ _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09194_ cpu.last_addr\[6\] _04216_ _04219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05426_ _00904_ net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08145_ cpu.uart.div_counter\[11\] _03399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05357_ _00836_ _00837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08076_ _03335_ _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09529__A1 _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05288_ _00750_ _00787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07027_ _02488_ _02118_ _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_30_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07095__C _02547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08978_ _04047_ _04040_ _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_59_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07929_ cpu.timer_top\[11\] _03217_ _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08504__A2 _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Left_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10305_ _00178_ clknet_leaf_105_wb_clk_i cpu.regs\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_72_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10236_ _00109_ clknet_leaf_121_wb_clk_i cpu.regs\[12\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09940__A1 net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10167_ _00044_ clknet_leaf_22_wb_clk_i cpu.uart.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08896__I _03985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10098_ _02092_ _05021_ _01629_ _05028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07305__I _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_32_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_32_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_72_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06260_ _01703_ _01721_ _01730_ net93 _01491_ _01731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_32_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05211_ _00002_ _00714_ _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06191_ _01661_ _01194_ _01191_ _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05142_ _00632_ _00644_ _00650_ _00651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_4_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09950_ net58 _04894_ _04903_ _04904_ _04905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05073_ net71 _00584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_40_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_49_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08901_ _02713_ _03987_ _03988_ _03990_ _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09931__A1 net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09881_ net73 _04853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08832_ _02751_ _03931_ _03932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05975_ _01423_ _01446_ _01447_ _01448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08763_ _03875_ _03877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_56_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07714_ _03049_ _03040_ _03050_ _00150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_95_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08694_ _03305_ _03825_ _03829_ _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_0_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07645_ _02971_ _03004_ _03008_ _00123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_0_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07576_ _01827_ _02958_ _02960_ _00102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_36_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09998__A1 _04047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09315_ _04327_ _04328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06527_ cpu.timer_top\[14\] _01465_ _01468_ _01995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09246_ _01852_ _01959_ _02086_ _04260_ _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_8_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06458_ _01925_ _01094_ _01333_ _01926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_106_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05409_ cpu.regs\[12\]\[2\] cpu.regs\[13\]\[2\] cpu.regs\[14\]\[2\] cpu.regs\[15\]\[2\]
+ _00830_ _00835_ _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_105_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09177_ cpu.ROM_addr_buff\[1\] _04206_ _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_88_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06389_ _01131_ _01840_ _01855_ _01857_ _01858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08128_ cpu.uart.div_counter\[5\] _03382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_43_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08059_ cpu.spi.data_out_buff\[6\] _03322_ _03320_ cpu.spi.data_out_buff\[7\] _03330_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput57 net57 io_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_113_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput46 net46 io_oeb[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput35 net35 io_oeb[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06984__A1 cpu.regs\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput68 net68 io_out[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput79 net79 io_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10021_ _04956_ _04957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09922__A1 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output58_I net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_106_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07161__A1 _01920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09989__A1 _04039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10219_ _00092_ clknet_leaf_0_wb_clk_i cpu.regs\[14\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05760_ _01186_ _01070_ _01234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_89_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05691_ _01164_ _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_76_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07430_ _02837_ _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06874__I _00710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07361_ cpu.timer_top\[5\] _02781_ _02785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09100_ _00884_ _04142_ _04147_ _04145_ _04148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_06312_ _00767_ _00960_ _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_33_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07292_ _00621_ _02727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09031_ _04087_ _04088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06243_ _01705_ _01712_ _01713_ _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06174_ _01143_ _01644_ _01645_ _00015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_5_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05218__A1 _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05125_ cpu.base_address\[0\] _00634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_111_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10064__C _02818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09933_ net81 _04888_ _02682_ _04893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05056_ cpu.IO_addr_buff\[1\] _00567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_110_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09864_ _04840_ _04841_ _00509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09904__A1 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08815_ _03896_ _03916_ _03917_ _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09795_ _04778_ _04782_ _00666_ _04785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05958_ cpu.PORTA_DDR\[1\] _01081_ _01429_ _01430_ _01431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_08746_ _03863_ _03864_ _03865_ _00367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_95_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08677_ cpu.toggle_ctr\[13\] _03816_ _03818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05889_ _01362_ _01352_ _01363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07628_ cpu.regs\[11\]\[4\] _02993_ _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07559_ _02017_ _02945_ _02949_ _00096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_101_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10570_ _00442_ clknet_leaf_81_wb_clk_i cpu.ROM_addr_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09229_ _00614_ _04245_ _04246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08932__C _04015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_112_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10004_ _02706_ _04936_ _04942_ _04939_ _00548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06185__A2 _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_103_Left_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09123__A2 _02129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08882__A1 _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09070__I _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_82_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08634__A1 _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_112_Left_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_91_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06930_ _02212_ _02372_ _02394_ _02396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__05620__A1 _01051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I io_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08600_ cpu.toggle_ctr\[4\] _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06861_ _02302_ _02304_ _02327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_89_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05812_ net75 _01279_ _01285_ _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06792_ _02256_ _02257_ _02258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09580_ _03135_ _00882_ _04585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_38_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05743_ _01216_ _01217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09114__A2 _03130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08531_ _03698_ _03699_ _00318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07125__A1 _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05674_ _00668_ _00610_ _01148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08462_ _00996_ _03642_ _03649_ _03646_ _00299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07413_ _02106_ _02566_ _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_65_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08393_ cpu.uart.receive_div_counter\[5\] _03581_ _03594_ _03566_ _03595_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07344_ _02771_ _02772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07275_ _02711_ _02712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09014_ _02893_ _04074_ _04075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_85_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06226_ _01601_ _01605_ _01696_ _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_26_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06939__A1 _02401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06157_ _01375_ _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06088_ _00607_ _01560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05108_ _00572_ _00618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09916_ _04077_ _04882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05611__A1 _01084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09847_ cpu.ROM_spi_dat_out\[3\] _04806_ _04828_ _04829_ _04830_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09778_ _02477_ cpu.startup_cycle\[0\] _04770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_96_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08729_ cpu.pwm_top\[5\] _03842_ _03854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07116__A1 _00989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05632__B _01097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07667__A2 _03019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10622_ _00494_ clknet_leaf_69_wb_clk_i cpu.startup_cycle\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10553_ _00425_ clknet_leaf_31_wb_clk_i cpu.uart.divisor\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10484_ _00357_ clknet_leaf_18_wb_clk_i cpu.pwm_top\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_114_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05461__S0 _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07313__I _02012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07658__A2 _03015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05133__A3 _00641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05390_ _00869_ _00870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_54_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07060_ _02519_ _02490_ _02520_ _02521_ _02522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_82_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06011_ cpu.Z _01484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_112_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05841__A1 _01310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09583__A2 _00821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09701_ cpu.last_addr\[9\] cpu.last_addr\[8\] _04700_ _04701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07962_ _03199_ _03208_ _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07893_ _03181_ _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09335__A2 _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06913_ _00807_ _00975_ _02379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09632_ _04634_ _04624_ _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06844_ _02291_ _02309_ _02310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09563_ _00978_ _04425_ _04568_ _04423_ _04569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09099__A1 _02549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08514_ _03685_ _03687_ _00313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06775_ cpu.regs\[1\]\[3\] _00948_ _02241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05726_ _01199_ _01200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_78_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09494_ _04455_ _04482_ _04501_ _04502_ _04503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08445_ cpu.had_int _03635_ cpu.needs_interrupt _03636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05657_ _01128_ _01130_ _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_08376_ _03574_ _03581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05588_ _01053_ _01054_ _01062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07327_ _02756_ _02741_ _02757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07258_ _02012_ _02698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_61_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09023__A1 _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06209_ cpu.toggle_top\[11\] _01274_ _01679_ _01580_ _01680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_07189_ _02332_ _02361_ _02640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_103_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07893__I _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09326__A2 _00651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05899__A1 _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05443__S0 _00828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output40_I net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06312__A2 _00960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10605_ _00477_ clknet_4_8_0_wb_clk_i cpu.PC\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_40_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10536_ _00409_ clknet_leaf_48_wb_clk_i cpu.spi.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_108_Right_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09014__A1 _02893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08899__I _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10467_ _00340_ clknet_leaf_8_wb_clk_i cpu.toggle_ctr\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10398_ _00271_ clknet_leaf_37_wb_clk_i cpu.uart.receiving vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_57_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_57_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_19_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06000__A1 _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07471__C _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06560_ _02023_ _02024_ _02026_ _02027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_86_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05511_ _00983_ cpu.instr_buff\[14\] _00984_ _00985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_06491_ _01948_ _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08230_ _03403_ _03456_ _03469_ _03470_ _03471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05442_ _00909_ _00919_ _00920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_117_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08161_ cpu.uart.data_buff\[0\] _03409_ _03414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09253__A1 _01585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05498__I _00973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05373_ _00852_ _00853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06067__A1 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08092_ cpu.uart.dout\[0\] _03353_ _00679_ _03354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07112_ _02568_ _02569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07043_ cpu.startup_cycle\[2\] _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08359__A3 _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08602__I cpu.toggle_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05417__I1 cpu.regs\[5\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08994_ _00618_ _02534_ _02537_ _04059_ _04060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__07218__I _02574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07945_ cpu.timer_top\[4\] _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07876_ _03171_ _00191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09615_ _04328_ _04605_ _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06827_ _00725_ _00899_ _02293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_66_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09546_ _04529_ _04445_ _04552_ _04476_ _04553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06758_ _02223_ _02215_ _02224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05709_ cpu.timer_div\[0\] _01183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09477_ _02401_ _00648_ _04486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08428_ cpu.uart.receive_div_counter\[12\] _03613_ _03622_ _03611_ _03623_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06689_ _02149_ _02153_ _02155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08359_ _02872_ _02931_ _03566_ _03349_ _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__09244__A1 _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10321_ _00194_ clknet_leaf_45_wb_clk_i cpu.spi.dout\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output88_I net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10252_ _00125_ clknet_leaf_119_wb_clk_i cpu.regs\[10\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10183_ _00060_ clknet_leaf_53_wb_clk_i cpu.timer_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06781__A2 _00869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05804__C _01277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_104_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_104_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_96_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05111__I _00620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10519_ _00392_ clknet_leaf_9_wb_clk_i cpu.timer\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07797__A1 _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_39_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08761__A3 _02763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05991_ _01258_ _01464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07730_ _03057_ _03062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_88_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09710__A2 cpu.ROM_addr_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07661_ _03017_ _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09400_ _04367_ _04401_ _04409_ _04411_ _04412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06612_ _02077_ _02078_ _02079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07592_ cpu.regs\[12\]\[1\] _02969_ _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06543_ _02006_ _02010_ _01479_ _02011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09331_ cpu.PC\[0\] cpu.br_rel_dest\[0\] _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06474_ _01848_ _01941_ _01942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09262_ _01113_ _02857_ _04276_ _04277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08213_ cpu.uart.div_counter\[3\] _03457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09193_ _04215_ _04217_ _04218_ _00461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_clkbuf_leaf_78_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05425_ _00881_ _00887_ _00903_ _00904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_16_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08144_ _02909_ _03396_ cpu.uart.div_counter\[3\] _01658_ _03397_ _03398_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_7_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05356_ _00835_ _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07788__A1 _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08075_ _03341_ _00220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_113_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05287_ _00786_ net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_07026_ _02117_ _02488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_101_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06212__A1 _00903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08977_ _00962_ _04047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_2_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_2_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07928_ cpu.timer\[11\] _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05691__I _01164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07859_ net20 _03114_ _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_3_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09529_ _02436_ _04449_ _04535_ _04536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_109_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09465__B2 _04453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09465__A1 _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05640__B _01097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09217__A1 cpu.ROM_addr_buff\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10304_ _00177_ clknet_leaf_107_wb_clk_i cpu.regs\[4\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10235_ _00108_ clknet_leaf_121_wb_clk_i cpu.regs\[12\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10166_ _00043_ clknet_leaf_41_wb_clk_i cpu.uart.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10097_ _01349_ _05025_ _05026_ _02073_ _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_16_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_112_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06190_ cpu.uart.divisor\[11\] _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05210_ cpu.regs\[4\]\[1\] cpu.regs\[5\]\[1\] cpu.regs\[6\]\[1\] cpu.regs\[7\]\[1\]
+ _00695_ _00696_ _00714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_106_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05141_ _00647_ _00649_ _00650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05072_ _00578_ _00579_ _00580_ _00582_ _00583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_09880_ _02533_ _04852_ _00514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_110_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_94_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08900_ _03943_ _03989_ _03990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08831_ _03228_ _03230_ _03920_ _03931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__05725__B _01198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05974_ _01011_ _01425_ _01447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08762_ _03875_ _03876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08498__A2 _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08693_ _03826_ _03827_ _03828_ _03829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_07713_ cpu.regs\[7\]\[4\] _03043_ _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07644_ cpu.regs\[10\]\[1\] _03007_ _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07575_ cpu.regs\[13\]\[4\] _02959_ _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_36_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07231__I _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06526_ _01989_ _01991_ _01993_ _01994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09314_ _01637_ _01343_ _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_90_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09245_ _01356_ _01596_ _01705_ _01785_ _04260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_06457_ _01328_ _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_8_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05408_ _00860_ _00885_ _00886_ _00887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09176_ _04202_ _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06388_ _01530_ _01856_ _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08127_ _02889_ _03378_ _03379_ _02679_ _03380_ _03381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05339_ _00819_ net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08058_ _02788_ _03308_ _03328_ _03329_ _00215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xoutput58 net58 io_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_07009_ net54 _02471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput47 net47 io_oeb[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06984__A2 _02128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput36 net36 io_oeb[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_31_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput69 net69 io_out[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10020_ _04955_ _02511_ _04956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09686__A1 _00773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06727__A2 _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10218_ _00091_ clknet_leaf_0_wb_clk_i cpu.regs\[14\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10149_ _00026_ clknet_4_10_0_wb_clk_i cpu.base_address\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08856__B _03912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05690_ _01158_ _01163_ _01164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__05163__A1 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07360_ _02783_ _02784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_9_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06311_ _00768_ _01781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_33_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07291_ _02710_ _02726_ _00051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09030_ _00632_ _01281_ _04087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_60_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06242_ _01705_ _01712_ _01530_ _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06173_ cpu.regs\[9\]\[2\] _01544_ _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_111_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05124_ cpu.base_address\[1\] _00633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09932_ _04892_ _00526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_111_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08168__A1 _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09863_ _02515_ _04803_ _04290_ _04841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_5_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09794_ _04761_ _04783_ _04784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_99_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08814_ cpu.timer_capture\[3\] _03899_ _03912_ _03917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08745_ cpu.timer_div_counter\[0\] cpu.timer_div_counter\[1\] cpu.timer_div_counter\[2\]
+ _03865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05957_ net80 _01003_ _01029_ _01080_ _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__09668__A1 _03708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08676_ _03795_ _03816_ _03817_ _00345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05888_ _00905_ _01361_ _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_67_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07627_ _02975_ _02990_ _02996_ _00117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_76_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07558_ cpu.regs\[14\]\[6\] _02946_ _02949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06509_ net13 _01226_ _01555_ _01977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_36_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07489_ cpu.uart.receive_div_counter\[14\] _02890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_101_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09228_ _04242_ _04244_ _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09159_ cpu.regs\[3\]\[5\] _03708_ _00669_ _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_31_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06406__A1 cpu.PORTB_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output70_I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10003_ cpu.PORTA_DDR\[7\] _04937_ _04942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07906__A1 cpu.timer_div\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06040__I _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07136__I _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08634__A2 _03786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08430__I _03503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05620__A2 _00593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06860_ _02325_ _02326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05811_ _01284_ _01285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08570__A1 _02811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06791_ _02222_ _02224_ _02257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_38_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05742_ _01024_ _01083_ _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08530_ _03136_ _03686_ _03689_ _03699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08322__B2 _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08461_ cpu.orig_IO_addr_buff\[2\] _03648_ _03649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05673_ _00595_ _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07125__A2 _02567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07412_ _02820_ _02821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_18_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08392_ cpu.uart.receive_div_counter\[5\] _03588_ _03589_ _03594_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_46_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07343_ _00665_ _02771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07274_ _01070_ _01242_ _01036_ _02673_ _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_103_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09013_ _04065_ _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06225_ _01602_ _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10075__C _03421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06156_ _01612_ _01616_ _01627_ _01628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06087_ cpu.uart.divisor\[10\] _01440_ _01559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05107_ _00614_ cpu.needs_timer_interrupt _00616_ _00617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09915_ net63 _04880_ _04881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07384__C _02697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09846_ _04049_ _04829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08561__A1 cpu.toggle_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09777_ _04768_ _04769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08496__B _03663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06989_ _02386_ _02439_ _02453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08728_ _02695_ _03844_ _03852_ _03853_ _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_08659_ cpu.toggle_ctr\[7\] _03803_ _03806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05632__C _00821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06875__A1 _02340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10621_ _00493_ clknet_leaf_69_wb_clk_i cpu.startup_cycle\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_91_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08616__A2 _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10552_ _00424_ clknet_leaf_40_wb_clk_i cpu.uart.divisor\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06627__A1 _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10483_ _00356_ clknet_leaf_19_wb_clk_i cpu.pwm_counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05461__S1 _00935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10111__A1 _03167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08607__A2 cpu.toggle_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06618__A1 _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07291__A1 _02710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06010_ _01480_ _01482_ _01306_ _01483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_23_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07961_ _03226_ _03249_ _03250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09700_ _04222_ _04699_ _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06912_ _02201_ _02202_ _02378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07892_ _03180_ _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09631_ _04298_ _04634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06843_ _02301_ _02307_ _02308_ _02309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_65_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09562_ _04390_ _04555_ _04567_ _04350_ _04568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06774_ _00725_ _00948_ _02240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05725_ cpu.uart.divisor\[0\] _01197_ _01198_ _01199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08513_ _02605_ _03686_ _03677_ _03687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_81_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09493_ _04399_ _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08444_ net17 _03635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05656_ _01129_ _01130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08375_ _02878_ _03569_ _03580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05587_ _01060_ _01061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07326_ cpu.timer\[7\] _02756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07257_ _02695_ _02676_ _02696_ _02697_ _00046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_5_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07188_ _01064_ _01311_ _02002_ _02639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06208_ _01676_ _01677_ _01678_ _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06139_ _01594_ _01611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08782__A1 cpu.timer_top\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05694__I _01009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09829_ _04807_ _04811_ _04814_ _04815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_69_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05443__S1 _00910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05520__A1 _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10604_ _00476_ clknet_leaf_91_wb_clk_i cpu.PC\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_40_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10535_ _00408_ clknet_leaf_47_wb_clk_i cpu.spi.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10466_ _00339_ clknet_leaf_8_wb_clk_i cpu.toggle_ctr\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_29_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10397_ _00270_ clknet_leaf_49_wb_clk_i cpu.uart.data_buff\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_97_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_97_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09804__I _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_26_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_26_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07328__A2 _02755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08525__A1 _02654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05510_ net98 _00984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06490_ _01957_ _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_28_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05511__A1 _00983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05441_ cpu.regs\[4\]\[3\] cpu.regs\[5\]\[3\] cpu.regs\[6\]\[3\] cpu.regs\[7\]\[3\]
+ _00918_ _00834_ _00919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA_clkbuf_leaf_68_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08160_ _03413_ _00239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09253__A2 _02684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07111_ _02567_ _02568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05372_ _00007_ _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08091_ _03350_ _03353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07042_ cpu.startup_cycle\[3\] _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_42_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08993_ _00615_ _04058_ _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07944_ cpu.timer_top\[3\] _03233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07875_ cpu.spi.dout\[1\] _03165_ _03169_ cpu.spi.data_in_buff\[1\] _03171_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09614_ _04368_ _04605_ _04617_ _04400_ _04618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06826_ _00689_ _00950_ _02292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09545_ _04478_ _04534_ _04536_ _04453_ _04551_ _04552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_06757_ cpu.regs\[1\]\[5\] _00898_ _02223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05708_ _01178_ _01181_ _01182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09476_ _02621_ _00647_ _04485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06688_ _02149_ _02153_ _02154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08427_ _02894_ _03621_ _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05639_ _01112_ _01113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08358_ _02919_ _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09244__A2 _02095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08289_ _03410_ _03516_ _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07255__A1 cpu.uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07309_ cpu.timer\[4\] _02741_ _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10320_ _00193_ clknet_leaf_44_wb_clk_i cpu.spi.dout\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10251_ _00124_ clknet_leaf_120_wb_clk_i cpu.regs\[10\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07007__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07558__A2 _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10182_ _00059_ clknet_leaf_21_wb_clk_i cpu.timer_top\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09624__I _04624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09180__A1 cpu.ROM_addr_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_102_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07494__A1 _02893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10518_ _00391_ clknet_leaf_26_wb_clk_i cpu.timer\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10449_ _00322_ clknet_leaf_81_wb_clk_i cpu.orig_PC\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07319__I _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05990_ cpu.timer_top\[1\] _01463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_88_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07660_ _02103_ _02965_ _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06611_ _01937_ _02021_ _02078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07591_ _01541_ _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_48_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06542_ _01474_ _01285_ _02009_ _02010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09330_ _04342_ _04343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09261_ _02436_ _02315_ _02297_ _02433_ _04276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_08212_ _03440_ _03456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06473_ _01349_ _01933_ _01940_ _01941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09192_ cpu.ROM_addr_buff\[5\] _04206_ _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05424_ _00902_ _00903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_7_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08143_ cpu.uart.div_counter\[2\] cpu.uart.divisor\[2\] _03397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05355_ _00834_ _00835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_113_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08074_ cpu.spi.data_in_buff\[2\] _03340_ _03336_ cpu.spi.data_in_buff\[3\] _03341_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_70_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07025_ cpu.mem_cycle\[5\] cpu.mem_cycle\[4\] _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_70_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05286_ _00785_ _00786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_30_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07229__I _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input32_I sram_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08976_ _04033_ _04046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06289__B _01758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07927_ _03206_ cpu.timer\[8\] _03208_ _03215_ _03216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_97_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07858_ _02591_ _02412_ _03153_ _03155_ _02626_ _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XTAP_TAPCELL_ROW_3_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06809_ _02271_ _02274_ _02275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07789_ _02601_ _02987_ _03098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09528_ _04404_ _04534_ _04535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_66_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09465__A2 _04448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09459_ _01778_ _04465_ _04468_ _04355_ _04469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05640__C _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10303_ _00176_ clknet_leaf_107_wb_clk_i cpu.regs\[4\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05368__B _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07139__I _02123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06451__A2 _01870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08728__A1 _02695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10234_ _00107_ clknet_leaf_1_wb_clk_i cpu.regs\[12\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10165_ _00042_ clknet_leaf_22_wb_clk_i cpu.uart.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07400__A1 _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05962__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09153__A1 _03703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10096_ _00907_ net96 net97 _01934_ _05026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_58_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07602__I _02967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05140_ _00648_ _00649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_12_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05071_ _00581_ _00582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_110_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_41_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_41_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_0_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08830_ _03894_ _03930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05973_ _01426_ _01441_ _01443_ _01445_ _01446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_08761_ _01179_ _01262_ _02763_ _03875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08692_ cpu.pwm_counter\[2\] _03828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07712_ _01825_ _03049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07643_ _03002_ _03007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09313_ _04325_ _04326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09447__A2 _04448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07574_ _02951_ _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06525_ _01992_ _01464_ _01169_ _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_36_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06130__A1 _01120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09244_ _01968_ _02095_ _04258_ _04259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_35_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06456_ _01119_ _01924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_113_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09175_ cpu.last_addr\[1\] _04199_ _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05407_ _00884_ _00874_ _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08958__A1 _02791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06572__B _01421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05967__I _01198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08126_ _02893_ cpu.uart.div_counter\[12\] _03380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06387_ _01838_ _01854_ _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07387__C _02697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10094__B _01638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05338_ cpu.ROM_OEB cpu.ROM_spi_mode _00819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08057_ cpu.spi.data_out_buff\[5\] _03322_ _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05269_ _00757_ _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_113_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput48 net48 io_oeb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_12_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07008_ _02462_ _02423_ _02463_ _02470_ _00024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xoutput37 net37 io_oeb[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput59 net59 io_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09383__A1 _01591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08959_ _01028_ _02674_ _04033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09902__I _04871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07449__A1 _02855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09349__I _04361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09610__A2 _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10217_ _00090_ clknet_leaf_0_wb_clk_i cpu.regs\[14\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10148_ _00025_ clknet_leaf_69_wb_clk_i net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05935__A1 cpu.regs\[9\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10079_ _02124_ _01517_ _02761_ _05009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05117__I _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07688__A1 cpu.regs\[8\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09429__A2 _04315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07290_ cpu.timer_capture\[1\] _02712_ _02725_ _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_33_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06310_ _01779_ _01137_ _01780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_61_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09687__C _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06241_ _00722_ _00730_ _00902_ _01613_ _01623_ _01712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_115_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06172_ _01643_ _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06415__A2 _01193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05123_ _00631_ _00632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07612__A1 cpu.regs\[12\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09931_ net80 _04887_ _04890_ _04891_ _04892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_41_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09862_ _02515_ _04803_ _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06179__B2 net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09793_ _04778_ _04782_ _04783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08813_ _02734_ _03910_ _03915_ _03891_ _03916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05956_ _01211_ _01429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08744_ cpu.timer_div_counter\[0\] cpu.timer_div_counter\[1\] cpu.timer_div_counter\[2\]
+ _03864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06567__B _00607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08675_ cpu.toggle_ctr\[12\] _03814_ _03817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07679__A1 _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05887_ _00877_ _01343_ _01361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__07242__I _02684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07626_ cpu.regs\[11\]\[3\] _02993_ _02996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07557_ _01922_ _02945_ _02948_ _00095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06508_ net4 _01436_ _01745_ _01976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_101_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07488_ cpu.uart.divisor\[14\] _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_91_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05697__I _00598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09227_ _04243_ _04244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06439_ cpu.regs\[4\]\[6\] cpu.regs\[5\]\[6\] cpu.regs\[6\]\[6\] cpu.regs\[7\]\[6\]
+ _01902_ _00935_ _01908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__07851__A1 _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09158_ _04190_ _00454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08109_ cpu.uart.receive_buff\[5\] _03366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06406__A2 _01039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09089_ _01111_ _04123_ _04138_ _04084_ _04139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_102_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05090__A1 _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output63_I net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08022__B net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10002_ _02701_ _04936_ _04941_ _04939_ _00547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_86_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_17_Left_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_30_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10018__I net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05400__I _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_26_Left_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05620__A3 _00641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05908__A1 _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05810_ _00984_ _01280_ _01283_ _01284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_38_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06790_ _02254_ _02255_ _02256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05741_ _01206_ _01215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08460_ _03640_ _03648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05672_ _01145_ _01146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08391_ _03591_ _03593_ _00284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07411_ _02321_ _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_35_Left_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_70_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07342_ cpu.timer_top\[1\] _02766_ _02770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07273_ _02574_ _02710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06636__A2 _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09012_ _04065_ _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06224_ _01693_ _01694_ _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_1_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06155_ _01132_ _01599_ _01621_ _01525_ _01626_ _01627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_13_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05106_ _00611_ _00615_ _00616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XPHY_EDGE_ROW_44_Left_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06086_ cpu.uart.divisor\[2\] _01230_ _01554_ _01557_ _01558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_09914_ _04871_ _04880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09845_ _04805_ _04811_ _04827_ _04828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07237__I _00664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09776_ cpu.startup_cycle\[2\] _04768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06988_ _02431_ _02443_ _02451_ _02452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08727_ _03724_ _03853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05939_ _01411_ _01412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_53_Left_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08658_ _03789_ _03805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_8_0_wb_clk_i clknet_0_wb_clk_i clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07609_ cpu.regs\[12\]\[6\] _02979_ _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08589_ cpu.toggle_ctr\[14\] _03743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06875__A2 _01477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10620_ _00492_ clknet_leaf_76_wb_clk_i cpu.mem_cycle\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10551_ _00423_ clknet_leaf_40_wb_clk_i cpu.uart.divisor\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10482_ _00355_ clknet_leaf_19_wb_clk_i cpu.pwm_counter\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_62_Left_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_19_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09577__A1 cpu.regs\[2\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06260__B1 net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09329__A1 _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08687__B _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06563__A1 _02027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_71_Left_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09362__I _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_58_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09568__A1 _00690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07960_ _03232_ _03248_ _03229_ _03249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06911_ _02161_ _02376_ _02377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07891_ _00664_ _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09630_ _04416_ _04627_ _04632_ _04386_ _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06842_ _02305_ _02306_ _02308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09561_ _03122_ _04427_ _04567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06773_ _02218_ _02232_ _02233_ _02239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA_clkbuf_leaf_97_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05724_ _01171_ _01017_ _01198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08512_ _03657_ _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09492_ _04471_ _04497_ _04500_ _04335_ _04501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__06306__A1 _00952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05305__I _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08443_ cpu.uart.receive_div_counter\[15\] _03631_ _03634_ _03585_ _00295_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_77_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05655_ _00820_ _00634_ _01129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08374_ _02877_ _03579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_92_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05586_ _00991_ _00642_ _01060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07325_ _02705_ _02755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_45_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07806__A1 cpu.regs\[3\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07256_ _02574_ _02697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_45_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06207_ cpu.toggle_top\[3\] _01416_ _01411_ _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06580__B _01075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07187_ _02637_ _02620_ _02638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06138_ _01504_ _01608_ _01609_ _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06069_ _01541_ _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09828_ _04812_ _04797_ _04813_ _04814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08534__A2 _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06545__A1 _02012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09759_ _02480_ _04753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_96_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10603_ _00475_ clknet_leaf_89_wb_clk_i cpu.PC\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_40_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10534_ _00407_ clknet_leaf_47_wb_clk_i cpu.spi.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10465_ _00338_ clknet_leaf_8_wb_clk_i cpu.toggle_ctr\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_20_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05885__I cpu.C vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10396_ _00269_ clknet_leaf_52_wb_clk_i cpu.uart.data_buff\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09970__A1 _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07605__I _01920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_66_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_66_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_86_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05440_ _00917_ _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__07340__I _01585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05371_ cpu.regs\[4\]\[0\] cpu.regs\[5\]\[0\] cpu.regs\[6\]\[0\] cpu.regs\[7\]\[0\]
+ _00832_ _00837_ _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_28_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07110_ _02535_ _02565_ _02566_ _02539_ _02567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__08880__B _03894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08090_ _03351_ _03352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_82_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07041_ _02484_ _02502_ _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_23_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09961__A1 _02685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08992_ _00586_ _00644_ _01055_ _01281_ _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XANTENNA__06775__A1 cpu.regs\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07943_ cpu.timer_top\[5\] _03228_ _03231_ cpu.timer_top\[4\] _03232_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07874_ _03170_ _00190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05744__B cpu.PORTA_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06527__A1 cpu.timer_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09613_ _04373_ _04607_ _04616_ _04397_ _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06825_ _02277_ _02286_ _02291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_97_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09544_ _04454_ _04550_ _04551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06756_ _02220_ _02221_ _02222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05707_ _01179_ _01180_ _01181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09475_ _02297_ _04449_ _04483_ _04484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06687_ _02151_ _02152_ _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_109_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08426_ _03617_ _03618_ _03621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05638_ cpu.br_rel_dest\[3\] _01112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08357_ _03565_ _00278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05569_ _01042_ _01043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08288_ _03507_ cpu.uart.counter\[1\] cpu.uart.counter\[2\] _03516_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07308_ _02714_ _02741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06058__A3 _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07239_ _02682_ _02683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_6_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10250_ _00123_ clknet_leaf_120_wb_clk_i cpu.regs\[10\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10181_ _00058_ clknet_leaf_53_wb_clk_i cpu.timer_top\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10116__I _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08507__A2 _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08965__B _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10078__A1 _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08994__A2 _02534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10517_ _00390_ clknet_leaf_26_wb_clk_i cpu.timer\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_113_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_113_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_110_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10002__A1 _02701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10448_ _00321_ clknet_leaf_83_wb_clk_i cpu.orig_PC\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09943__A1 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10379_ _00252_ clknet_leaf_29_wb_clk_i cpu.uart.div_counter\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06757__A1 cpu.regs\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07182__A1 _02297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05732__A2 _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_9_Left_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06610_ _01948_ _01964_ _02077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07590_ _02964_ _02968_ _02970_ _00106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_87_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06541_ _02008_ _02009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08131__B1 cpu.uart.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09260_ _01105_ _02821_ _04273_ _04274_ _04275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06472_ _01348_ _01939_ _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08211_ _03451_ _03452_ _03455_ _03450_ _00242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__07070__I _02531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05496__A1 _00825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05423_ _00901_ _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_117_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09191_ cpu.last_addr\[5\] _04216_ _04217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_99_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08142_ _03392_ _03396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05354_ _00833_ _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08073_ _03333_ _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05285_ _00769_ _00778_ _00784_ _00785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_15_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07024_ _02111_ _02113_ _02486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05799__A2 _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09934__A1 _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06748__A1 cpu.regs\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08975_ _04045_ _00416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07926_ _03211_ _03214_ _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input25_I rst_n vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07857_ _03154_ _02371_ _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07173__A1 _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06808_ _00770_ _00870_ _02274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07788_ _02985_ _03092_ _03097_ _00177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09527_ _04533_ _04534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06739_ _02204_ _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_109_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09458_ _04093_ _04447_ _04466_ _04467_ _04468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_19_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08409_ _03605_ _03575_ _03607_ _03566_ _03608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09389_ _04368_ _04371_ _04398_ _04400_ _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_50_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output93_I net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10302_ _00175_ clknet_leaf_106_wb_clk_i cpu.regs\[4\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10233_ _00106_ clknet_leaf_1_wb_clk_i cpu.regs\[12\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10164_ _00041_ clknet_leaf_102_wb_clk_i cpu.br_rel_dest\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05384__B _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10095_ _02065_ _02069_ _02064_ _05025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_58_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05070_ cpu.startup_cycle\[3\] cpu.startup_cycle\[2\] cpu.startup_cycle\[1\] cpu.startup_cycle\[0\]
+ _00581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_40_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_6_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_10_0_wb_clk_i clknet_0_wb_clk_i clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__05294__B _00707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05972_ _01444_ _01426_ _01445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08760_ _03861_ _03874_ _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_81_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_81_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_73_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08691_ cpu.pwm_counter\[1\] _03827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07711_ _03047_ _03039_ _03048_ _00149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07642_ _02964_ _03004_ _03006_ _00122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_0_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09312_ _04293_ _04325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07573_ _02951_ _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06524_ cpu.timer_top\[6\] _01992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06455_ _01408_ _01922_ _01923_ _00018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06130__A2 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09243_ _01822_ _01869_ _04257_ _04258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09174_ _04193_ _04200_ _04204_ _00456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_44_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06386_ _01852_ _01854_ _01855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05406_ _00884_ _00874_ _00885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08125_ cpu.uart.div_counter\[1\] _03379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05337_ cpu.PORTB_DDR\[0\] net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_44_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06969__A1 _02433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08056_ cpu.spi.data_out_buff\[6\] _03320_ _03328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05268_ _00768_ net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XANTENNA__09907__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput49 net49 io_oeb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_05199_ _00703_ net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_07007_ net20 _02132_ _02419_ _02469_ _02470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xoutput38 net38 io_oeb[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07394__A1 _02695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08958_ _02791_ _04027_ _04032_ _00412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07909_ cpu.timer\[9\] _03198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08889_ _03980_ _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_106_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05632__A1 _01105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10216_ _00089_ clknet_leaf_37_wb_clk_i cpu.uart.receive_counter\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05935__A2 _01408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10147_ _00024_ clknet_leaf_99_wb_clk_i cpu.regs\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10078_ _03305_ _05007_ _05008_ _00556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__05491__S0 _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07137__A1 _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_99_Left_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06240_ _01523_ _01698_ _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10202__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06171_ _01642_ _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_111_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05122_ cpu.br_rel_dest\[7\] _00630_ _00631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09930_ _04111_ _04891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_68_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09275__I _00678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09861_ _04839_ _00508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06179__A2 _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09792_ _04781_ _04770_ _04782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08812_ _02734_ _03914_ _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05955_ _01196_ _01428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08743_ _03860_ _03863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08674_ cpu.toggle_ctr\[12\] _03814_ _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05886_ _01349_ _01353_ _01358_ _01359_ _01360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_95_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07625_ _02973_ _02990_ _02995_ _00116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07556_ cpu.regs\[14\]\[5\] _02946_ _02948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06507_ net66 _01078_ _01208_ _01974_ _01225_ _01975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_76_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07487_ cpu.uart.divisor\[14\] _02886_ cpu.uart.receive_div_counter\[13\] _02880_
+ _02887_ _02888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_91_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09226_ _00660_ _01148_ _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06583__B _01009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06438_ _01904_ _01906_ _01907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09157_ cpu.ROM_addr_buff\[12\] _04189_ _04181_ _04190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06369_ _01836_ _01837_ _01838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_31_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08108_ _03364_ _03361_ _03365_ _00229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08800__A1 _03259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09088_ _02755_ _04086_ _04137_ _04138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08039_ cpu.spi.data_out_buff\[1\] _03314_ _03316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07367__A1 _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10001_ cpu.PORTA_DDR\[6\] _04937_ _04941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_output56_I net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09913__I _04871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_67_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_48_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05853__A1 _01186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07101__C _02547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05605__A1 _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07608__I _02016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07358__A1 _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_87_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05740_ net79 _01172_ _01213_ _01084_ _01214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_77_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07343__I _00665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05671_ _01144_ _01118_ _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05216__S0 _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08390_ _03588_ _03589_ _03592_ _03593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07410_ _02578_ _02817_ _02579_ _02819_ _00077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_18_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07341_ _02768_ _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_73_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07272_ _02709_ _00049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09011_ _02690_ _04066_ _04072_ _04070_ _00425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09035__A1 _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05844__A1 _01229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06223_ _01112_ _00749_ _01694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06154_ _01622_ _01606_ _01624_ _01625_ _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XPHY_EDGE_ROW_103_Right_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05105_ _00584_ net18 _00615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_41_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06085_ _01556_ _01557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09913_ _04871_ _04879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09844_ cpu.ROM_spi_dat_out\[2\] _02527_ _04827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09775_ _02533_ _04767_ _00494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06987_ _02392_ _02441_ _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05938_ _01178_ _01012_ _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__07253__I _00962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08726_ cpu.pwm_top\[4\] _03847_ _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08657_ _03796_ _03803_ _03804_ _00339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05869_ _00633_ _00588_ _01343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07608_ _02016_ _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08588_ cpu.toggle_ctr\[15\] _03742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_63_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07539_ _01138_ _02936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_107_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10550_ _00422_ clknet_leaf_41_wb_clk_i cpu.uart.divisor\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09209_ _04228_ _04203_ _04229_ _03421_ _00466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_10481_ _00354_ clknet_leaf_102_wb_clk_i cpu.pwm_counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06260__B2 _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_121_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_4_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06000__C _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08068__A2 _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06079__A1 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10679_ _00551_ clknet_leaf_69_wb_clk_i net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06251__A1 _00722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05685__S0 _00917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06910_ _00772_ _02009_ _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07890_ _03179_ _00197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_65_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06841_ _02305_ _02306_ _02307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08169__I _00665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09560_ _04386_ _04564_ _04565_ _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06772_ _02213_ _02237_ _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05723_ _01196_ _01197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08511_ cpu.orig_PC\[4\] _03684_ _03685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09491_ _04498_ _04482_ _04499_ _04500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08442_ _02890_ _03632_ cpu.uart.receive_div_counter\[15\] _03634_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_93_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05654_ _01126_ _01127_ _01128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08373_ _03504_ _03578_ _00281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05585_ _01040_ _01058_ _01059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07324_ _02749_ _02754_ _00056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_34_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09008__A1 _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07255_ cpu.uart.divisor\[4\] _02677_ _02696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05817__A1 _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06206_ cpu.pwm_top\[3\] _01268_ _01270_ _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07186_ _02636_ _02637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06137_ _01504_ _01608_ _01361_ _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07248__I _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06068_ _01490_ _01540_ _01541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_111_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05991__I _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09827_ _04766_ _04751_ _04813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09758_ _04751_ _04752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_68_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08709_ _03624_ _03839_ _00356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_69_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09689_ _04669_ _04689_ _04251_ _00486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09495__A1 _04454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10602_ _00474_ clknet_leaf_89_wb_clk_i cpu.PC\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_40_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10533_ _00406_ clknet_leaf_48_wb_clk_i cpu.spi.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05231__I _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10464_ _00337_ clknet_leaf_8_wb_clk_i cpu.toggle_ctr\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_20_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10395_ _00268_ clknet_leaf_52_wb_clk_i cpu.uart.data_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_75_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07621__I _02988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10096__A2 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05511__A3 _00984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05370_ _00843_ _00849_ _00850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_28_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_35_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_35_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_43_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07040_ cpu.startup_cycle\[5\] _02474_ _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08452__I _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08991_ _04057_ _00420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07972__A1 _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06775__A2 _00948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07942_ _03230_ _03231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07873_ cpu.spi.dout\[0\] _03165_ _03169_ cpu.spi.data_in_buff\[0\] _03170_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09713__A2 cpu.ROM_addr_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09612_ _04612_ _04615_ _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06824_ _02266_ _02289_ _02290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09543_ _04455_ _04534_ _04549_ _04502_ _04550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05750__A3 _01005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09477__A1 _02401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06755_ _02144_ _02173_ _02172_ _02221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_78_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05706_ _01027_ _01180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09474_ _04450_ _04482_ _04483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06686_ _00762_ _00974_ _02152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08425_ _03609_ _03620_ _00291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05637_ _01110_ _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_19_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08356_ cpu.uart.receive_buff\[6\] _03554_ _03562_ cpu.uart.receive_buff\[7\] _03565_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_93_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05568_ _01021_ _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07307_ _02711_ _02740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08287_ _03515_ _00258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05986__I _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05499_ _00974_ _00975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07238_ _02681_ _02682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07169_ cpu.PC\[5\] _02621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06215__A1 _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09952__A2 _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10180_ _00057_ clknet_leaf_30_wb_clk_i cpu.timer_capture\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07706__I _01642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08965__C _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08140__A1 _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09640__A1 _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08272__I _00620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10516_ _00389_ clknet_leaf_26_wb_clk_i cpu.timer\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10447_ _00320_ clknet_leaf_82_wb_clk_i cpu.orig_PC\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10378_ _00251_ clknet_leaf_29_wb_clk_i cpu.uart.div_counter\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06757__A2 _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07616__I _02988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09459__A1 _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06540_ _02007_ _02008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06471_ _01935_ _01938_ _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08210_ cpu.uart.div_counter\[2\] _03453_ _03454_ _03448_ _03455_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06693__A1 _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05422_ _00900_ _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_28_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09190_ _04197_ _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_99_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08141_ _03390_ _02704_ _02906_ _03391_ _03394_ _03395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_56_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05353_ _00005_ _00833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08072_ _03339_ _00219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_113_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05284_ _00757_ _00781_ _00783_ _00784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_113_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07023_ _02484_ _02481_ _00582_ _02485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_3_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08974_ cpu.timer_div\[3\] _04035_ _04044_ _04015_ _04045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_11_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_89_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07925_ _03212_ cpu.timer\[14\] cpu.timer\[13\] _03213_ _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07856_ _02238_ _02370_ _03154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input18_I io_in[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06807_ _00799_ _00855_ _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07787_ cpu.regs\[4\]\[7\] _03093_ _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_66_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09526_ _04531_ _04532_ _04533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06738_ _02199_ _02203_ _02204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08122__B2 _02891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09457_ _04349_ _04467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08408_ _03605_ _03601_ _03607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_98_Right_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06669_ _02134_ _02135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_108_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09388_ _04399_ _04400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_50_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08339_ _02922_ _03349_ _03554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_74_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10127__I _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10301_ _00174_ clknet_leaf_106_wb_clk_i cpu.regs\[4\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10232_ _00105_ clknet_leaf_111_wb_clk_i cpu.regs\[13\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10163_ _00040_ clknet_leaf_102_wb_clk_i cpu.br_rel_dest\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10094_ _00820_ _05019_ _01638_ _05024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_107_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_83_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06675__A1 _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06427__A1 cpu.timer_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07346__I _02685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05971_ cpu.uart.dout\[1\] _01444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07710_ cpu.regs\[7\]\[3\] _03043_ _03048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08690_ cpu.pwm_counter\[0\] _03826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07641_ cpu.regs\[10\]\[0\] _03005_ _03006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_76_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07572_ _01736_ _02952_ _02957_ _00101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_50_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_50_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_87_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06523_ _01260_ _01990_ _01991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09311_ _02555_ _04324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07081__I _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06454_ cpu.regs\[9\]\[5\] _01142_ _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09242_ _01639_ _01731_ _04256_ _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_29_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09173_ cpu.ROM_addr_buff\[0\] _04203_ _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06385_ _01785_ _01803_ _01853_ _01854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05405_ _00883_ _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08124_ cpu.uart.div_counter\[14\] _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05336_ cpu.PORTA_DDR\[0\] net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_71_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09080__A2 _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06969__A2 _02009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08055_ _02784_ _03309_ _03327_ _00214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05267_ _00767_ _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05198_ _00682_ _00693_ _00702_ _00703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_07006_ _02417_ _02427_ _02468_ _02469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xoutput39 net39 io_oeb[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07256__I _02574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08957_ cpu.spi.divisor\[7\] _04028_ _04032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07908_ _03196_ _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08888_ cpu.timer_capture\[14\] _03959_ _03978_ _03979_ _03980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_55_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07839_ net12 _03121_ _03134_ _03138_ _03139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_TAPCELL_ROW_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_38_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05504__I _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09509_ _04383_ _04509_ _04517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_117_Right_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06409__A1 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05880__A2 _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08550__I _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05632__A2 _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10215_ _00088_ clknet_leaf_36_wb_clk_i cpu.uart.receive_counter\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06070__I _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10146_ _00023_ clknet_leaf_98_wb_clk_i cpu.regs\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_89_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_77_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10077_ _02713_ _01058_ _04036_ _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__05491__S1 _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08334__B2 _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07137__A2 _02133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06170_ _01593_ _01641_ _01642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_68_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05121_ cpu.br_rel_dest\[6\] _00630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09860_ cpu.ROM_spi_dat_out\[7\] _04807_ _04838_ _04829_ _04839_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_68_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09791_ _02476_ _04768_ _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08811_ cpu.timer\[0\] cpu.timer\[1\] cpu.timer\[2\] _03914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05954_ cpu.uart.divisor\[1\] _01427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08742_ _03861_ _03862_ _00366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08325__A1 _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08673_ _03795_ _03814_ _03815_ _00344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07624_ cpu.regs\[11\]\[2\] _02993_ _02995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05885_ cpu.C _01359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07555_ _01827_ _02945_ _02947_ _00094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_118_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07486_ cpu.uart.receive_div_counter\[4\] cpu.uart.divisor\[4\] _02887_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06506_ _01429_ _01971_ _01972_ _01973_ _01974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_75_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09225_ _00625_ _04241_ _04242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06437_ _00824_ _01905_ _00846_ _01906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_33_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09156_ cpu.regs\[3\]\[4\] _02414_ _04167_ _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06368_ _00786_ _00976_ _01837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08107_ cpu.uart.dout\[4\] _03358_ _03362_ _03365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09087_ cpu.orig_IO_addr_buff\[7\] _04090_ _04137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06299_ _01738_ _01412_ _01768_ _01277_ _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_05319_ _00816_ _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08038_ _02760_ _03309_ _03315_ _00209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_111_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10000_ _02698_ _04936_ _04940_ _04939_ _00546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_101_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09989_ _04039_ _04929_ _04933_ _04932_ _00542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_99_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10123__A1 _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05225__S1 _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08619__A2 _01413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10129_ _01826_ _05050_ _05052_ _00563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_89_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08858__A2 cpu.timer\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05670_ _00570_ _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09807__A1 _04098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07340_ _01585_ _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_58_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07271_ _02704_ _02689_ _02707_ _02708_ _02709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_100_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09010_ cpu.uart.divisor\[11\] _04067_ _04072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06222_ _01112_ _00749_ _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_26_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06153_ _01530_ _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08404__B _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05104_ _00613_ _00614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_111_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06084_ net8 _01226_ _01555_ _01556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09912_ _02690_ _04872_ _04878_ _04875_ _00520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__05319__I _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09843_ _04826_ _00503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09235__B _04251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09774_ _04766_ _04762_ _04767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06986_ _02417_ _02427_ _02450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05780__A1 _01174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08725_ _02806_ _03843_ _03851_ _03846_ _00360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05937_ cpu.toggle_top\[9\] _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08656_ _03765_ _03801_ _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05868_ _01340_ _01341_ _01342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08587_ _03735_ _03736_ _03737_ _03740_ _03741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_07607_ _02981_ _02978_ _02982_ _00111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05799_ _01261_ _01011_ _01008_ _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_49_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07538_ _01102_ _01108_ _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07469_ _02871_ _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07285__A1 _02710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09208_ cpu.ROM_addr_buff\[10\] _04202_ _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10480_ _00353_ clknet_leaf_102_wb_clk_i cpu.pwm_counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09139_ _04176_ _00449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07709__I _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_107_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_107_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_94_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_43_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10678_ _00550_ clknet_leaf_73_wb_clk_i cpu.ROM_OEB vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_35_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07579__A2 _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06251__A2 _00730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08528__A1 _03696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05139__I cpu.br_rel_dest\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06840_ _02281_ _02282_ _02306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07354__I _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06771_ _02218_ _02235_ _02236_ _02237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05722_ _01195_ _01057_ _01196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08510_ _03654_ _03684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09490_ cpu.orig_PC\[5\] _04236_ _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08441_ _03631_ _03633_ _00294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_81_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05653_ _00640_ _01127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08372_ _02878_ _03576_ _03577_ _03571_ _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_105_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05584_ _01006_ _01057_ _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_85_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07323_ cpu.timer_capture\[6\] _02738_ _02753_ _02754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07254_ _02694_ _02695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06205_ cpu.timer_top\[11\] _01465_ _01177_ _01675_ _01676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_54_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07185_ _02400_ _02636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06136_ _01346_ _01599_ _01607_ _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06067_ net27 _01334_ _01539_ _01403_ _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_09826_ _04808_ _04812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09757_ cpu.startup_cycle\[0\] _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_100_Left_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05753__A1 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06969_ _02433_ _02009_ _02434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07742__A2 _03060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_5_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_5_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08708_ cpu.pwm_counter\[7\] _03838_ _03839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_96_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09688_ _04413_ _04685_ _04688_ _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05505__A1 _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08639_ _03711_ _03751_ cpu.toggle_ctr\[1\] _03792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_83_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10601_ _00473_ clknet_leaf_89_wb_clk_i cpu.PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10532_ _00405_ clknet_leaf_48_wb_clk_i cpu.spi.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10463_ _00336_ clknet_leaf_8_wb_clk_i cpu.toggle_ctr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06481__A2 _01914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10394_ _00267_ clknet_leaf_52_wb_clk_i cpu.uart.data_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_75_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09183__A1 cpu.ROM_addr_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07497__A1 _02893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10096__A3 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07349__I _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09410__A2 _04420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08990_ cpu.timer_div\[7\] _04046_ _04056_ _04050_ _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07972__A2 _00616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07941_ cpu.timer\[4\] _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07872_ _03168_ _03169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06202__B _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09611_ _00881_ _04388_ _04614_ _04423_ _04615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06823_ _02277_ _02286_ _02288_ _02289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09542_ _04372_ _04538_ _04548_ _04471_ _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06754_ _02144_ _02219_ _02220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05705_ _01043_ _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09473_ _04481_ _04482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06685_ _02143_ _02150_ _02151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08424_ _03617_ _03613_ _03619_ _03611_ _03620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05332__I cpu.PORTB_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05636_ _01053_ _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08355_ _03564_ _00277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05567_ _01018_ _01034_ _01037_ _01040_ _01041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_19_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07306_ _02714_ _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08286_ cpu.uart.counter\[1\] _03513_ _03514_ _02708_ _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05498_ _00973_ _00974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07237_ _00664_ _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_104_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07168_ _02406_ _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06119_ _01120_ _01591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07099_ net20 _02543_ _02557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__05974__A1 _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09809_ _02503_ _04754_ _04795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_70_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08553__I _03713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10515_ _00388_ clknet_leaf_27_wb_clk_i cpu.timer\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07651__A1 _02977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06454__A2 _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10446_ _00319_ clknet_leaf_82_wb_clk_i cpu.orig_PC\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07403__A1 _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10377_ _00250_ clknet_leaf_32_wb_clk_i cpu.uart.div_counter\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05965__A1 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05732__A4 _01205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06470_ _01937_ _01842_ _01938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05421_ _00899_ _00900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08140_ _02909_ _03392_ _03393_ _03394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05352_ _00831_ _00832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_08071_ cpu.spi.data_in_buff\[1\] _03334_ _03336_ cpu.spi.data_in_buff\[2\] _03339_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_70_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07642__A1 _02964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05283_ _00750_ _00782_ _00783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07022_ _02480_ _02484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_3_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08973_ _02775_ _04040_ _04044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07924_ cpu.timer_top\[13\] _03213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07855_ _03152_ _02410_ _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_108_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06806_ _00772_ _00872_ _02271_ _02272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__07542__I _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07786_ _03053_ _03092_ _03096_ _00176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_94_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_28_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09525_ _02654_ _04530_ _04532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06737_ _02201_ _02202_ _02203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_66_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09456_ _02604_ _04389_ _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06668_ _01287_ _02133_ _02134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08407_ _03605_ _03606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05619_ _01092_ _01093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09387_ _00983_ _03310_ _04399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06599_ _02065_ _02066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_22_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08338_ _02921_ _03352_ _00271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09622__A2 _04624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08269_ _03498_ _03501_ _00254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07633__A1 _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10300_ _00173_ clknet_leaf_13_wb_clk_i cpu.regs\[4\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10231_ _00104_ clknet_leaf_111_wb_clk_i cpu.regs\[13\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output79_I net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10162_ _00039_ clknet_leaf_101_wb_clk_i cpu.br_rel_dest\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_67_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10093_ _01518_ _05022_ _05023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06372__A1 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09310__A1 _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10429_ _00302_ clknet_leaf_54_wb_clk_i cpu.orig_IO_addr_buff\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07927__A2 cpu.timer\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05970_ _01442_ _01194_ _01443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_57_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05166__A2 cpu.needs_timer_interrupt vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07362__I _02771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07640_ _03002_ _03005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07571_ cpu.regs\[13\]\[3\] _02953_ _02957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09310_ _03624_ _04323_ _00473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06522_ cpu.timer_capture\[14\] _01256_ _01990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06453_ _01921_ _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09241_ _01402_ _01539_ _04255_ _04256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_28_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_103_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09172_ _04202_ _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_90_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_90_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_56_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06384_ _01781_ _00945_ _01853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05404_ _00882_ _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08123_ _03374_ cpu.uart.divisor\[6\] _01881_ cpu.uart.div_counter\[5\] _03376_ _03377_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05335_ cpu.PORTA_DDR\[7\] net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_08054_ cpu.spi.data_out_buff\[4\] _03322_ _03320_ cpu.spi.data_out_buff\[5\] _03327_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_98_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_101_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07005_ _02452_ _02464_ _02466_ _02455_ _02467_ _02468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05266_ _00756_ _00760_ _00766_ _00757_ _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA__09368__A1 cpu.PC\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05197_ _00003_ _00698_ _00701_ _00702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__08591__A2 _01275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input30_I sram_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08956_ _02788_ _04027_ _04031_ _00411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06441__I2 cpu.regs\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07907_ _03183_ _03184_ _03192_ _03195_ _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_08887_ _03947_ _03979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09540__A1 _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07838_ _02409_ _03137_ _03120_ _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_55_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09508_ _02400_ _01119_ _04515_ _04516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_07769_ _03085_ _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09439_ _04329_ _04449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_35_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06409__A2 _01221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10214_ _00087_ clknet_leaf_37_wb_clk_i cpu.uart.receive_counter\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08582__A2 _01738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10145_ _00022_ clknet_leaf_99_wb_clk_i cpu.regs\[2\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06593__A1 _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10076_ _01058_ _04036_ net75 _05007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05148__A2 _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_10_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09598__A1 _03136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05120_ _00628_ _00629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08022__A1 _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08810_ _03896_ _03911_ _03913_ _00383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09790_ _04764_ _04758_ _04780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05953_ _01002_ _01425_ _01426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_84_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08741_ _03188_ cpu.timer_div_counter\[1\] _03862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08672_ cpu.toggle_ctr\[11\] _03812_ _03815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05884_ _01357_ _01349_ _01358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07623_ _02971_ _02990_ _02994_ _00115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_105_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06887__A2 _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07554_ cpu.regs\[14\]\[4\] _02946_ _02947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07485_ cpu.uart.receive_div_counter\[14\] _02886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06505_ cpu.PORTB_DDR\[6\] _01003_ _01741_ _01973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09224_ _04238_ _04240_ _04082_ _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06436_ cpu.regs\[12\]\[6\] cpu.regs\[13\]\[6\] cpu.regs\[14\]\[6\] cpu.regs\[15\]\[6\]
+ _01902_ _01153_ _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_8_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09155_ _04188_ _00453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06367_ _01832_ _01772_ _01836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08106_ cpu.uart.receive_buff\[4\] _03364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09086_ _04122_ _04135_ _04136_ _00436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06298_ cpu.toggle_top\[4\] _01417_ _01412_ _01767_ _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_05318_ _00769_ _00810_ _00815_ _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_08037_ cpu.spi.data_out_buff\[0\] _03314_ _03315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05496__B _00853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05249_ _00732_ _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_101_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06171__I _01642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09988_ cpu.PORTA_DDR\[1\] _04930_ _04933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06575__A1 cpu.timer_capture\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05217__I3 cpu.regs\[15\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08939_ _04020_ _04021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09513__A1 _01924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10694_ _00566_ clknet_leaf_112_wb_clk_i cpu.regs\[15\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05250__I _00733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05853__A3 _01203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09392__I _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10128_ cpu.regs\[15\]\[4\] _05051_ _05052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10059_ _04808_ _04991_ _04992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09504__A1 _04238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_29_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_29_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_89_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07640__I _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07270_ _02546_ _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05160__I net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08491__A1 _00672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06221_ _01690_ _01691_ _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06152_ _01596_ _01623_ _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06083_ _01196_ _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09991__A1 _03849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05103_ cpu.TIE _00613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09911_ net62 _04873_ _04878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_111_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09842_ cpu.ROM_spi_dat_out\[2\] _04806_ _04825_ _04736_ _04826_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06557__A1 net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_13_Left_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_111_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09773_ _04755_ _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08724_ cpu.pwm_top\[3\] _03847_ _03851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06985_ _02015_ _02423_ _02449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05936_ _01143_ _01407_ _01409_ _00013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08655_ cpu.toggle_ctr\[6\] _03801_ _03803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05867_ _00883_ _00634_ _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08586_ _03738_ cpu.toggle_top\[13\] cpu.toggle_top\[12\] _03739_ _03740_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07606_ cpu.regs\[12\]\[5\] _02979_ _02982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09259__B1 _02855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07537_ _02934_ _00089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05798_ _01167_ _01168_ _01267_ _01271_ _01272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XPHY_EDGE_ROW_22_Left_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07468_ _00619_ _02871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06419_ _01885_ _01886_ _01887_ _01888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09207_ cpu.last_addr\[10\] _04228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07399_ cpu.toggle_top\[14\] _02797_ _02814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09138_ cpu.ROM_addr_buff\[7\] _04175_ _04169_ _04176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09069_ _02624_ _04122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_31_Left_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08537__A2 _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output61_I net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06076__I net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10677_ _00549_ clknet_leaf_73_wb_clk_i cpu.ROM_spi_mode vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_82_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09973__A1 _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06251__A3 _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09725__A1 cpu.ROM_addr_buff\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05211__A1 _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06770_ _02232_ _02234_ _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05721_ _01038_ _01029_ _01195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08440_ _02890_ _03632_ _03592_ _03633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05652_ _00639_ _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_58_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08371_ _02878_ _03569_ _03577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_105_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05583_ _01013_ _01042_ _01057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_58_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07322_ _02739_ _02750_ _02740_ _02752_ _02753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07253_ _00962_ _02694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_61_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06204_ _01672_ _01673_ _01674_ _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07184_ _02015_ _02612_ _02635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__10023__A1 cpu.ROM_addr_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09964__A1 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06135_ _01346_ _01606_ _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06066_ _01492_ _01538_ _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_10_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09825_ _04808_ _04810_ _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09756_ _04747_ _04744_ _04750_ _00492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05753__A2 _01225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06968_ _00800_ _02433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_96_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09687_ _04402_ _04672_ _04687_ _04439_ _02761_ _04688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08707_ _03836_ _03834_ _03838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05919_ _01381_ _01384_ _01388_ _01370_ _01391_ _01392_ _01393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08638_ cpu.toggle_clkdiv cpu.toggle_ctr\[1\] cpu.toggle_ctr\[0\] _03791_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06899_ _02266_ _02289_ _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05505__A2 _00979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08569_ _01872_ _03722_ _03726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_92_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10600_ _00472_ clknet_leaf_89_wb_clk_i cpu.Z vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_12_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10531_ _00404_ clknet_leaf_25_wb_clk_i cpu.timer_capture\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_40_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10462_ _00335_ clknet_leaf_7_wb_clk_i cpu.toggle_ctr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10393_ _00266_ clknet_leaf_52_wb_clk_i cpu.uart.data_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_20_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08930__A2 _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08694__A1 _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08446__A1 _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09946__A1 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_7_0_wb_clk_i clknet_0_wb_clk_i clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07940_ cpu.timer_top\[6\] _03227_ _03228_ cpu.timer_top\[5\] _03229_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xclkbuf_leaf_44_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_44_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07365__I _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07871_ _00620_ _03167_ _03168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09610_ _04094_ _04604_ _04613_ _04392_ _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06822_ _02287_ _02285_ _02288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09541_ _04544_ _04547_ _04548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06753_ cpu.regs\[1\]\[0\] _00973_ _02219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05704_ _01173_ _01178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09472_ _02621_ _04480_ _04481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06684_ _00740_ _01927_ _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08423_ _03617_ _03618_ _03619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05635_ _01102_ _01108_ _01109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08354_ cpu.uart.receive_buff\[5\] _03554_ _03562_ cpu.uart.receive_buff\[6\] _03564_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_86_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05566_ _01039_ _01040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07305_ _02711_ _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08285_ _03508_ cpu.uart.counter\[1\] _03499_ _03514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05497_ _00966_ _00968_ _00970_ _00972_ _00973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_07236_ _00875_ _02677_ _02680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09937__A1 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07167_ _02615_ _02618_ _02619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06118_ _00672_ _01589_ _01093_ _01590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_100_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07098_ _02555_ _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_57_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07275__I _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06049_ _01130_ _01366_ _01522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09808_ _02512_ _04793_ _04794_ _00500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_70_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09739_ _04737_ _00488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_4_15_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10514_ _00387_ clknet_leaf_30_wb_clk_i cpu.timer\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_96_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09928__A1 _02760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10445_ _00318_ clknet_leaf_83_wb_clk_i cpu.orig_PC\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05662__A1 _01000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10376_ _00249_ clknet_leaf_33_wb_clk_i cpu.uart.div_counter\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05965__A2 _01000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06914__A1 _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05420_ _00898_ _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_56_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05351_ _00830_ _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_99_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08070_ _03338_ _00218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05282_ cpu.regs\[12\]\[5\] cpu.regs\[13\]\[5\] cpu.regs\[14\]\[5\] cpu.regs\[15\]\[5\]
+ _00752_ _00754_ _00782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_3_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06264__I _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07021_ _02475_ _02476_ _02479_ _02482_ _02483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__09919__A1 _02698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08972_ _01546_ _04035_ _04043_ _04038_ _00415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07923_ cpu.timer_top\[14\] _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07854_ cpu.PC\[11\] _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08919__I _03985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06805_ _02242_ _02267_ _02269_ _02270_ _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_79_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07785_ cpu.regs\[4\]\[6\] _03093_ _03096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_108_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09524_ _02653_ _04530_ _04531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06736_ _00799_ _00975_ _02202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05343__I _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09455_ _04349_ _04465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06667_ _00593_ _01637_ _01130_ _02133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_38_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08406_ cpu.uart.receive_div_counter\[8\] _03605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05618_ _01000_ _01068_ _01074_ _01091_ _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_19_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09386_ _04373_ _04376_ _04396_ _04397_ _04398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06598_ _00816_ _01164_ _02065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_19_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08337_ _03553_ _00270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05549_ _01022_ _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09083__A1 _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08268_ _03378_ _03500_ _03464_ _03501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_34_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07219_ _02571_ _02663_ _02665_ _02666_ _00039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_15_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08199_ _03445_ _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10230_ _00103_ clknet_leaf_114_wb_clk_i cpu.regs\[13\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07397__A1 _02811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Left_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10161_ _00038_ clknet_leaf_102_wb_clk_i cpu.br_rel_dest\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10092_ _02086_ _02079_ _05021_ _05022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_58_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05253__I _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08564__I _03713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09395__I _04293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10428_ _00301_ clknet_leaf_90_wb_clk_i cpu.orig_IO_addr_buff\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10359_ _00232_ clknet_leaf_39_wb_clk_i cpu.uart.dout\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06060__A1 _01309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08888__A1 cpu.timer_capture\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07643__I _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_69_Left_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07570_ _01644_ _02952_ _02956_ _00100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_76_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06521_ _01460_ _01987_ _01988_ _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_118_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09240_ _01491_ _01385_ _04255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06452_ _01920_ _01921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_103_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09171_ _04201_ _04202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09065__A1 _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06383_ _01838_ _01852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05403_ cpu.base_address\[1\] _00882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08122_ _02883_ cpu.uart.div_counter\[9\] _03375_ _02891_ _03376_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_05334_ cpu.PORTB_DDR\[7\] net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_71_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08053_ _03324_ _03326_ _00213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_78_Left_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07004_ _02453_ _02459_ _02467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05265_ _00764_ _00765_ _00732_ _00766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07379__A1 _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05196_ _00699_ _00700_ _00701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08955_ cpu.spi.divisor\[6\] _04028_ _04031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07906_ cpu.timer_div\[6\] _03193_ cpu.timer_div_counter\[7\] _03187_ _03194_ _03195_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__06441__I3 cpu.regs\[3\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input23_I io_in[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08886_ _03204_ _03918_ _03901_ _03977_ _03978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07553__I _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06354__A2 _01823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07837_ _03136_ _02408_ _02626_ _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_55_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07768_ _02966_ _03036_ _03085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_94_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05073__I net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09507_ _04513_ _04488_ _04514_ _04515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06719_ _02155_ _02156_ _02185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07699_ _03037_ _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_109_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09438_ _04447_ _04448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_35_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07221__C _02666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09369_ _04379_ _04344_ _04380_ _04381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05617__A1 _01075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output91_I net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10213_ _00086_ clknet_leaf_38_wb_clk_i cpu.uart.receive_counter\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06042__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10144_ _00021_ clknet_leaf_98_wb_clk_i cpu.regs\[2\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_100_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06593__A2 _02021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05396__A3 _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10075_ _04998_ _05004_ _05006_ _03421_ _00555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_89_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09531__A2 _04534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_qcpu_110 io_out[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_97_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09598__A2 _04443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07638__I _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05084__A2 _00593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08022__A2 _03167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05158__I _00665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07373__I _02793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05952_ _01320_ _01424_ _01207_ _01425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_08740_ cpu.timer_div_counter\[0\] _03861_ _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08671_ cpu.toggle_ctr\[11\] _03812_ _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05883_ _01354_ _01356_ _01357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_23_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07622_ cpu.regs\[11\]\[1\] _02993_ _02994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_105_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07553_ _02938_ _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07484_ _02033_ _02885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06504_ net57 _01171_ _01213_ _01083_ _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_64_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09223_ _04239_ _04240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09038__A1 _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06435_ _00841_ _01903_ _01904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_17_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_86_Left_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09154_ _02521_ _04187_ _04181_ _04188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_60_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08105_ _03360_ _03361_ _03363_ _00228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06366_ _01701_ _01793_ _01835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09085_ cpu.IO_addr_buff\[6\] _03446_ _04127_ _04136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06297_ _01764_ _01765_ _01766_ _01767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_44_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05317_ _00769_ _00812_ _00814_ _00815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__09249__B _04263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08036_ _03313_ _03314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06272__A1 cpu.PORTB_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05248_ _00749_ net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_4_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06452__I _01920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05179_ _00683_ _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_95_Left_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09987_ _03840_ _04929_ _04931_ _04932_ _00541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_08938_ _02871_ _01023_ _03638_ _03415_ _04020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XTAP_TAPCELL_ROW_4_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08869_ _03909_ _03963_ _03904_ _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10693_ _00565_ clknet_leaf_112_wb_clk_i cpu.regs\[15\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10127_ _05043_ _05051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10058_ _04946_ _04986_ _04988_ _04990_ _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_89_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_69_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_69_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05829__A1 _00874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06220_ _01595_ _01598_ _01611_ _01691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_38_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06151_ _00718_ _01513_ _01529_ _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_26_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06082_ _01552_ _01553_ _01554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07368__I _02705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05102_ cpu.instr_cycle\[3\] _00611_ _00612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09910_ _03849_ _04872_ _04877_ _04875_ _00519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_95_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09841_ _04777_ _04823_ _04824_ _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09772_ _04762_ _04765_ _02683_ _00493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_111_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08199__I _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06984_ cpu.regs\[2\]\[6\] _02128_ _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08723_ _03849_ _03843_ _03850_ _03846_ _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05935_ cpu.regs\[9\]\[0\] _01408_ _01409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07506__B2 _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08654_ _03796_ _03801_ _03802_ _00338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05866_ _01127_ _01340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05797_ cpu.pwm_top\[0\] _01269_ _01270_ _01271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08585_ cpu.toggle_ctr\[12\] _03739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07605_ _01920_ _02981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09259__B2 _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07536_ _02930_ _02933_ _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07052__B _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05351__I _00830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09206_ _04215_ _04226_ _04227_ _00465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08482__A2 _03655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07467_ _02571_ _02870_ _02665_ _02819_ _00083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_106_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06418_ cpu.spi.divisor\[5\] _01244_ _01887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07398_ _02750_ _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_8_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09137_ _02654_ _04063_ _04174_ _04175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06349_ net94 _01818_ _01819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09982__A2 _03712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09068_ _04081_ _04120_ _04121_ _00433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09431__B2 _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08019_ cpu.spi.counter\[0\] _03299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07745__A1 _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output54_I net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06357__I _01826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09670__A1 cpu.PC\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10676_ _00548_ clknet_leaf_59_wb_clk_i cpu.PORTA_DDR\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05720_ _01193_ _01194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_81_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05651_ _01051_ _01125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08370_ _03575_ _03576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_86_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05171__I _00677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07321_ _02751_ _02741_ _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05582_ _01051_ _00643_ _01052_ _01055_ _01056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07252_ _02693_ _00045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06203_ cpu.timer_top\[3\] _01260_ _01263_ _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07183_ _02613_ _02629_ _02634_ _00035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_53_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06134_ _01603_ _01605_ _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06065_ _01504_ _01506_ _01510_ _01537_ _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA_clkbuf_leaf_47_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09716__A2 cpu.ROM_addr_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09824_ _04809_ _04801_ _04810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05346__I _00825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09755_ _04747_ _04744_ _04748_ _04749_ _00666_ _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06967_ _02383_ _02386_ _02432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09686_ _00773_ _04450_ _04686_ _04687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08706_ _03836_ _03834_ _03837_ _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06898_ _02331_ _02362_ _02363_ _02364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05918_ _01380_ _01392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05849_ _01043_ _01180_ _01008_ _01045_ _01322_ _01323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_68_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08637_ _03789_ _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06177__I net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08568_ _02695_ _03721_ _03723_ _03725_ _00329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07519_ _02918_ net15 _02920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08499_ _03662_ _03677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09652__A1 cpu.PC\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10530_ _00403_ clknet_leaf_25_wb_clk_i cpu.timer_capture\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_40_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_86_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10461_ _00334_ clknet_4_1_0_wb_clk_i cpu.toggle_ctr\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08207__A2 _03391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06218__A1 _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10392_ _00265_ clknet_leaf_51_wb_clk_i cpu.uart.data_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_20_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05965__B _01229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08567__I _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08446__A2 _00616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09643__A1 _03703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09398__I _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10659_ _00531_ clknet_leaf_60_wb_clk_i net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__06209__A1 cpu.toggle_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05968__B1 _01438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07870_ _03166_ _03167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06821_ _02284_ _02287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_84_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_84_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_50_Left_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09540_ _01111_ _04465_ _04546_ _04355_ _04547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06752_ _00806_ _00871_ _02217_ _02218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_05703_ _01176_ _01177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07381__I _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09471_ _02401_ _04479_ _04480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_13_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_13_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08422_ _02910_ _03614_ _03618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08685__A2 _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06683_ _02143_ _02144_ _02147_ _02148_ _02149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_116_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_120_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05634_ _01103_ _00986_ _01107_ _01108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_08353_ _03563_ _00276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05565_ _01038_ _01039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09634__A1 _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08284_ _03507_ _03499_ _03512_ _03509_ _03513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07304_ _02727_ _02737_ _00053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06448__A1 _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07235_ _01427_ _02679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05496_ _00825_ _00971_ _00853_ _00972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_81_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07166_ _02616_ _02617_ _02618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05785__B _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07097_ _00983_ _02555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06117_ _01056_ _01589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06620__A1 _01396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06048_ _01516_ _01520_ _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07999_ cpu.spi.div_counter\[1\] _03282_ _03286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09807_ _04098_ _02516_ _04794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09738_ _02117_ _04692_ _04735_ _04736_ _04737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_96_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09669_ _02398_ _02412_ _04479_ _04670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_65_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09625__A1 _03701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_53_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10513_ _00386_ clknet_leaf_23_wb_clk_i cpu.timer\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07100__A2 _02557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10444_ _00317_ clknet_leaf_82_wb_clk_i cpu.orig_PC\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10375_ _00248_ clknet_leaf_33_wb_clk_i cpu.uart.div_counter\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06678__A1 cpu.regs\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09616__A1 _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05350_ _00829_ _00830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_28_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_112_Right_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05281_ _00779_ _00780_ _00781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07020_ _02480_ _02481_ _02482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_12_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07376__I _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08971_ _00903_ _04040_ _04043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07922_ cpu.timer_top\[13\] _03209_ _03210_ cpu.timer_top\[12\] _03211_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07853_ _03142_ _03151_ _00188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06804_ _00740_ _00899_ _02270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__05264__S1 _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07784_ _03051_ _03092_ _03095_ _00175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05624__I _01097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09523_ _02400_ _02828_ _02406_ _04530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06735_ _02198_ _02200_ _02201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_78_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09454_ _04458_ _04462_ _04463_ _04347_ _04464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06666_ _02122_ _02132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08405_ _03603_ _03604_ _00287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09385_ _04340_ _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05617_ _01075_ _01078_ _01090_ _01091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_47_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08336_ cpu.uart.data_buff\[9\] _03520_ _03525_ _03553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_52_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06597_ _00816_ _01164_ _02064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_22_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05548_ _00994_ _01021_ _01022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_50_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08267_ _03494_ _03499_ _03436_ _03490_ _03500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_61_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05479_ _00947_ _00955_ _00956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_34_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08198_ _00677_ _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07218_ _02574_ _02666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07149_ _02600_ _02601_ _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06404__B cpu.PORTA_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07286__I _01585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07219__C _02666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10160_ _00037_ clknet_leaf_99_wb_clk_i cpu.regs\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10091_ net97 _01165_ _05021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09006__I _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_106_Left_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08845__I cpu.timer\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_85_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08580__I cpu.toggle_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06832__A1 _00762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05635__A2 _01108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10427_ _00300_ clknet_leaf_55_wb_clk_i cpu.orig_IO_addr_buff\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_115_Left_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05709__I cpu.timer_div\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10358_ _00231_ clknet_leaf_42_wb_clk_i cpu.uart.dout\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10289_ _00162_ clknet_leaf_3_wb_clk_i cpu.regs\[5\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_94_Right_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07924__I cpu.timer_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07560__A2 _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06520_ cpu.timer_capture\[6\] _01420_ _01988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_87_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06451_ _01831_ _01870_ _01919_ _01920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_118_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05402_ _00880_ _00881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09170_ _04194_ _00627_ _04195_ _04201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06382_ _01833_ _01850_ _01851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08121_ cpu.uart.div_counter\[8\] _03375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05333_ cpu.PORTA_DDR\[6\] net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__07076__A1 _00627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08052_ cpu.spi.data_out_buff\[3\] _03301_ _03325_ _03326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_98_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05264_ cpu.regs\[4\]\[4\] cpu.regs\[5\]\[4\] cpu.regs\[6\]\[4\] cpu.regs\[7\]\[4\]
+ _00751_ _00753_ _00765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_31_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07003_ _02380_ _02465_ _02466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05182__S0 _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05619__I _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05195_ cpu.regs\[8\]\[0\] cpu.regs\[9\]\[0\] cpu.regs\[10\]\[0\] cpu.regs\[11\]\[0\]
+ _00695_ _00696_ _00700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08954_ _02784_ _04027_ _04030_ _00410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07905_ _01546_ cpu.timer_div_counter\[2\] _03193_ cpu.timer_div\[6\] _03194_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08885_ _03919_ _03976_ _03977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10135__A1 _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07000__A1 cpu.regs\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09128__I0 _00773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07836_ _03135_ _03136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input16_I io_in[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07767_ _02462_ _03083_ _03084_ _00169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09506_ cpu.PC\[5\] _00645_ _04514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06718_ _02177_ _02183_ _02184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08500__A1 _02831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07698_ _03038_ _03039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06649_ cpu.mem_cycle\[5\] _02114_ _02115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_82_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09437_ _02604_ _04446_ _04447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__05314__A1 _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05303__B _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09368_ cpu.PC\[1\] _00988_ _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08319_ _01321_ _03311_ _03539_ _03540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_09299_ _04311_ _04312_ _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05617__A2 _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05529__I _00993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10212_ _00085_ clknet_leaf_13_wb_clk_i _00003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_30_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10143_ _00020_ clknet_leaf_110_wb_clk_i cpu.regs\[9\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06042__A2 _00873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10074_ _04998_ _05005_ net77 _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08575__I cpu.toggle_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_qcpu_100 io_oeb[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_qcpu_111 io_out[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_69_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09047__A2 _04098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10062__B1 _00627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08558__A1 _02800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07230__A1 _01005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input8_I io_in[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05951_ _00605_ _01424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_84_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05882_ _01355_ _01356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08670_ _03805_ _03812_ _03813_ _00343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08730__A1 _02811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07621_ _02988_ _02993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_105_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07552_ _02938_ _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06503_ _01215_ _01217_ cpu.PORTA_DDR\[6\] _01971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_75_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07483_ _02880_ cpu.uart.receive_div_counter\[13\] _02881_ cpu.uart.divisor\[5\]
+ _02882_ _02883_ _02884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_76_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09222_ _00650_ _01055_ _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06434_ cpu.regs\[8\]\[6\] cpu.regs\[9\]\[6\] cpu.regs\[10\]\[6\] cpu.regs\[11\]\[6\]
+ _01902_ _01153_ _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_17_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09153_ _03703_ _04173_ _04186_ _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_60_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06365_ _01361_ _01834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08104_ cpu.uart.dout\[3\] _03358_ _03362_ _03363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05316_ _00787_ _00813_ _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09084_ _01924_ _04123_ _04134_ _04084_ _04135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06296_ cpu.pwm_top\[4\] _01269_ _01168_ _01766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08035_ _03312_ _03300_ _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06272__A2 _01039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05247_ _00748_ _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05349__I _00828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05178_ _00000_ _00683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_101_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09986_ _04077_ _04932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07564__I _02951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08937_ _04019_ _00404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10108__A1 _04453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08868_ _03960_ _03962_ _03963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07819_ _02107_ _03113_ _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_98_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08799_ _03898_ _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10692_ _00564_ clknet_leaf_112_wb_clk_i cpu.regs\[15\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06129__B _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05310__I1 _00807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07460__A1 _02135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06263__A2 _01732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09201__A2 _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07212__A1 _02534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10126_ _05043_ _05050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07407__C _02818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10057_ _04753_ _04989_ _04756_ _00580_ _04990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_89_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10035__B1 _04969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08779__A1 _02784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_38_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_38_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06150_ _01522_ _01622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_110_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06081_ net23 _01436_ _01228_ _01553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05101_ _00610_ _00611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_37_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05169__I _00663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09840_ cpu.ROM_spi_dat_out\[1\] _04790_ _04824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09771_ _04751_ _04764_ _04765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05765__A1 cpu.uart.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06983_ _01921_ _02423_ _02424_ _02447_ _00022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_111_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08722_ cpu.pwm_top\[2\] _03847_ _03850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05934_ _01141_ _01408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_28_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08653_ cpu.toggle_ctr\[5\] _03799_ _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05865_ _01338_ _01339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_89_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05796_ _01009_ _01270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08584_ cpu.toggle_ctr\[13\] _03738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07604_ _02977_ _02978_ _02980_ _00110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09259__A2 _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07535_ _00620_ _02875_ _02931_ _02932_ _02933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__09104__I _04150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07466_ _02560_ _02870_ _02664_ _02819_ _00082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_06417_ cpu.uart.dout\[5\] _01560_ _01665_ _01886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09205_ cpu.ROM_addr_buff\[9\] _04220_ _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_76_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07397_ _02811_ _02796_ _02812_ _02810_ _00071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09136_ _04173_ cpu.regs\[2\]\[7\] _04174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09431__A2 _04422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06348_ _01817_ _01807_ _01818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06279_ cpu.uart.divisor\[4\] _01749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09067_ _01019_ _04112_ _04103_ _04121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_32_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08018_ _03280_ _03298_ _00206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08942__A1 _02760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09969_ _04906_ _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_99_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output47_I net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05508__A1 net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10675_ _00547_ clknet_leaf_86_wb_clk_i cpu.PORTA_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09422__A2 _04415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07433__A1 _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09617__C _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05717__I _00607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10109_ _01359_ _05009_ _05038_ _04098_ _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_65_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05650_ _01123_ _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06548__I _02015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05581_ _01053_ _01054_ _01055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_clkbuf_leaf_110_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07320_ cpu.timer\[6\] _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_85_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08763__I _03875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07251_ cpu.uart.divisor\[3\] _02689_ _02692_ _02687_ _02693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_45_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06202_ cpu.timer_capture\[11\] _01256_ _01258_ _01673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_60_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07182_ _02297_ _02633_ _02634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_103_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09413__A2 _04422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06133_ _01498_ _01499_ _01604_ _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_26_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07424__A1 _02831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06064_ _01521_ _01532_ _01536_ _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09177__A1 cpu.ROM_addr_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09823_ _02479_ _04776_ _04782_ _04809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09754_ _04694_ _04749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06966_ _02430_ _02395_ _02431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_09685_ _04328_ _04672_ _04686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08705_ _03836_ _03834_ _03371_ _03837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06897_ _02309_ _02291_ _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05917_ _01390_ _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_96_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05848_ _01321_ _01026_ _01023_ _01019_ _01322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_08636_ _03180_ _03786_ _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05779_ _01182_ _01247_ _01249_ _01252_ _01253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_76_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08567_ _03724_ _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07518_ _02918_ _02916_ _02919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08498_ cpu.orig_PC\[0\] _03672_ _03676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09652__A2 _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07663__A1 _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07449_ _02855_ _02827_ _02856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10460_ _00333_ clknet_leaf_8_wb_clk_i cpu.toggle_ctr\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09119_ _04161_ _00444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06218__A2 _00951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10391_ _00264_ clknet_leaf_51_wb_clk_i cpu.uart.data_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08915__A1 cpu.timer_capture\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08143__A2 cpu.uart.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09340__A1 _02848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06154__A1 _01622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06154__B2 _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09643__A2 _04554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07654__A1 cpu.regs\[10\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10658_ _00530_ clknet_leaf_60_wb_clk_i net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_82_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10589_ _00461_ clknet_leaf_80_wb_clk_i cpu.last_addr\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05968__A1 _01427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06831__I _00772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08906__A1 cpu.timer_capture\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05447__I _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06393__B2 _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06820_ _02284_ _02285_ _02286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06751_ _02187_ _02214_ _02216_ _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05702_ _01173_ _01175_ _01176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09331__A1 cpu.PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06682_ _00740_ _00974_ _02148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09470_ _04446_ _04479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08421_ cpu.uart.receive_div_counter\[11\] _03617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05633_ _01106_ _01107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08352_ cpu.uart.receive_buff\[4\] _03554_ _03562_ cpu.uart.receive_buff\[5\] _03563_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05564_ _00993_ _01038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_86_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_53_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_53_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08493__I _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08283_ cpu.uart.counter\[3\] cpu.uart.counter\[2\] _03439_ _03512_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_74_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07303_ cpu.timer_capture\[3\] _02712_ _02736_ _02737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06448__A2 _01901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07645__A1 _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05495_ cpu.regs\[4\]\[5\] cpu.regs\[5\]\[5\] cpu.regs\[6\]\[5\] cpu.regs\[7\]\[5\]
+ _00918_ _00834_ _00971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_07234_ _02671_ _02676_ _02678_ _02666_ _00042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_61_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07165_ _02596_ _02361_ _02617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05959__A1 _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06116_ _01583_ _01586_ _01587_ _01588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07096_ _02554_ _00028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06047_ _01387_ _01497_ _01519_ _01507_ _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_100_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07998_ cpu.spi.div_counter\[1\] _03282_ _03285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09806_ _04759_ _04793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09273__B _04263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09737_ _04049_ _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06949_ _02414_ _02412_ _02415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06188__I _01198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09668_ _03708_ _04292_ _04669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08619_ _03748_ _01413_ _03752_ _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09599_ _04603_ _00482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_25_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07240__C _02683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07636__A1 _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10512_ _00385_ clknet_leaf_23_wb_clk_i cpu.timer\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10443_ _00316_ clknet_leaf_82_wb_clk_i cpu.orig_PC\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05662__A3 _01074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10374_ _00247_ clknet_leaf_33_wb_clk_i cpu.uart.div_counter\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06611__A2 _02021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05267__I _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09561__A1 _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05280_ cpu.regs\[8\]\[5\] cpu.regs\[9\]\[5\] cpu.regs\[10\]\[5\] cpu.regs\[11\]\[5\]
+ _00752_ _00754_ _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_15_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06602__A2 _01914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08970_ _04042_ _00414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05177__I _00003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_100_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_100_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09805__C _04792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07921_ cpu.timer\[12\] _03210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07852_ _01593_ _01641_ _02105_ _03150_ _03151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xinput1 io_in[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06803_ _02240_ _02268_ _02269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_78_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09304__A1 _04293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09522_ cpu.PC\[7\] _04529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07783_ cpu.regs\[4\]\[5\] _03093_ _03095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_108_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06118__A1 _00672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06734_ _00770_ _01928_ _02200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09453_ _04377_ _04447_ _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06665_ net1 _02131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08404_ cpu.uart.receive_div_counter\[7\] _03600_ _03592_ _03604_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05616_ _01082_ _01086_ _01089_ _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09384_ _04387_ _04395_ _04396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08335_ _03552_ _00269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09607__A2 _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06596_ _00817_ _01935_ _02063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_22_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05547_ _01020_ cpu.IO_addr_buff\[0\] _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08266_ _03407_ _03499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05478_ _00953_ _00929_ _00954_ _00955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07094__A2 _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08197_ _03443_ _03444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07217_ _01830_ _02662_ _02665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07148_ _01116_ _01124_ _01138_ _02601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_112_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07079_ _02535_ _02120_ _02121_ _02539_ _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_72_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10090_ _05019_ _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_58_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06109__A1 cpu.toggle_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10426_ _00299_ clknet_leaf_55_wb_clk_i cpu.orig_IO_addr_buff\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09782__A1 _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10357_ _00230_ clknet_leaf_43_wb_clk_i cpu.uart.dout\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10288_ _00161_ clknet_leaf_108_wb_clk_i cpu.regs\[6\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07848__A1 _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08257__B _03464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06450_ _00946_ _01584_ _01485_ _01918_ _01919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_118_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06520__A1 cpu.timer_capture\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05401_ _00879_ _00880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06381_ _01781_ _01817_ _01807_ _01850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08120_ cpu.uart.div_counter\[6\] _03374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05332_ cpu.PORTB_DDR\[6\] net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08051_ _02778_ _03307_ _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05263_ cpu.regs\[0\]\[4\] _00763_ cpu.regs\[2\]\[4\] cpu.regs\[3\]\[4\] _00751_
+ _00753_ _00764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_113_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07002_ _02458_ _02465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05194_ _00692_ _00699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06587__A1 _02053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08953_ cpu.spi.divisor\[5\] _04028_ _04030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07904_ cpu.timer_div_counter\[6\] _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__09525__A1 _02654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08884_ _03203_ _03975_ _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07000__A2 _02128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07835_ cpu.PC\[9\] _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09128__I1 _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07766_ cpu.regs\[5\]\[7\] _03083_ _03084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_69_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09505_ cpu.PC\[5\] _00596_ _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06717_ _02178_ _02182_ _02183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07839__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07697_ _03037_ _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09436_ _02828_ _02404_ _04446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06648_ cpu.mem_cycle\[4\] _02114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_93_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06579_ cpu.timer_top\[7\] _02046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09367_ cpu.PC\[1\] _00988_ _04379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08318_ _03407_ _03411_ _03539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_74_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09298_ _00652_ _02762_ _04312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08249_ _03396_ _03480_ _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06578__A1 _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10211_ _00084_ clknet_leaf_13_wb_clk_i _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output77_I net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10142_ _00019_ clknet_leaf_112_wb_clk_i cpu.regs\[9\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10073_ _04795_ _04796_ _05002_ _04801_ _05005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08319__A2 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09017__I _02531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_qcpu_101 io_oeb[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_84_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_qcpu_112 io_oeb[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_65_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05459__I3 cpu.regs\[11\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10409_ _00282_ clknet_leaf_34_wb_clk_i cpu.uart.receive_div_counter\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05950_ cpu.uart.has_byte _01423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05881_ _01338_ _00857_ _01355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07620_ _02964_ _02990_ _02992_ _00114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_23_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07551_ _01736_ _02939_ _02944_ _00093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06502_ _00982_ _01968_ _01969_ _01970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_07482_ _01442_ _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_76_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_66_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09221_ _04237_ _04238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_17_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06433_ _00827_ _01902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_29_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09152_ _03637_ cpu.regs\[3\]\[3\] _04186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_60_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06364_ _01832_ _01833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08103_ _02681_ _03362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05315_ cpu.regs\[12\]\[7\] cpu.regs\[13\]\[7\] cpu.regs\[14\]\[7\] cpu.regs\[15\]\[7\]
+ _00794_ _00795_ _00813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09083_ _02750_ _04086_ _04133_ _04134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06295_ cpu.timer_top\[12\] _01170_ _01468_ _01765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08034_ _02871_ _03262_ _03311_ _03312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05246_ _00736_ _00739_ _00745_ _00747_ _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_31_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08549__A2 _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05177_ _00003_ _00682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_12_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09985_ cpu.PORTA_DDR\[0\] _04930_ _04931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08936_ cpu.timer_capture\[15\] _04003_ _04018_ _04015_ _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_4_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05365__I _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08867_ _03907_ _03961_ _03962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07818_ _03115_ _03119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08798_ _02723_ _03892_ _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_8_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_8_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06732__A1 _00762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07749_ _03071_ _03074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_80_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09419_ _01646_ _04425_ _04429_ _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10691_ _00563_ clknet_leaf_113_wb_clk_i cpu.regs\[15\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09985__A1 cpu.PORTA_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06263__A3 _01733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05310__I2 cpu.regs\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05275__I _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10125_ _01735_ _05044_ _05049_ _00562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10056_ _02502_ _04781_ _04989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_100_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09976__A1 _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06080_ net61 _01434_ _01550_ _01551_ _01224_ _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_05100_ _00608_ _00609_ _00610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_111_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_78_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_78_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09770_ _02473_ _04763_ _04764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_107_Right_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06982_ net12 _02132_ _02419_ _02446_ _02447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_111_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08721_ _02685_ _03849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05933_ _01406_ _01407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08652_ cpu.toggle_ctr\[5\] _03799_ _03801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05517__A2 _00608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07603_ cpu.regs\[12\]\[4\] _02979_ _02980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05864_ _00703_ _01338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_37_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05795_ _01268_ _01269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08583_ cpu.toggle_ctr\[10\] _03730_ _01410_ cpu.toggle_ctr\[9\] _03737_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07534_ cpu.uart.receive_counter\[3\] _02932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_66_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07465_ _02662_ _02870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_8_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06416_ _01880_ _01882_ _01884_ _01885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08445__B cpu.needs_interrupt vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09204_ cpu.last_addr\[9\] _04216_ _04226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07396_ cpu.toggle_top\[13\] _02797_ _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09135_ _03637_ _04173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06347_ _01715_ _01727_ _01817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06278_ _01744_ _01746_ _01747_ _01748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09066_ _01646_ _04096_ _04119_ _04109_ _04120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07442__A2 _02848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08017_ cpu.spi.div_counter\[7\] _03297_ _03298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05229_ _00731_ net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_102_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09968_ _04906_ _04918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08919_ _03985_ _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09899_ net89 _04869_ _00656_ _04829_ _04870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06705__A1 _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10017__A1 _03432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10674_ _00546_ clknet_leaf_86_wb_clk_i cpu.PORTA_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09958__A1 _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10109__C _04098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06944__A1 cpu.PC\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10108_ _04453_ _05020_ _05037_ _05009_ _05038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_10039_ cpu.ROM_addr_buff\[10\] _02524_ _04973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05580_ cpu.br_rel_dest\[6\] _01054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_105_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07250_ _02690_ _02691_ _02692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10008__A1 _03432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06201_ cpu.timer_capture\[3\] _01569_ _01252_ _01671_ _01672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_42_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07181_ _02632_ _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06132_ _00988_ _00718_ _01604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_113_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07395__I _02745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06063_ _01367_ _01534_ _01535_ _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_10_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09822_ _04759_ _04808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09753_ _04196_ _04693_ _04748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08704_ cpu.pwm_counter\[6\] _03836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06965_ _02373_ _02393_ _02430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09684_ _04362_ _04672_ _04684_ _04436_ _04685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05916_ _01389_ _01390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06896_ _02332_ _02361_ _02362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05643__I _01116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05847_ _01001_ _01320_ _01321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08635_ _03788_ _00333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08566_ _02573_ _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10201__D _00074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07517_ cpu.uart.receiving _02918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05778_ _01251_ _01252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08497_ _03673_ _03675_ _00308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07448_ _00726_ _02855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_91_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07379_ _02794_ _02799_ _00066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09118_ cpu.ROM_addr_buff\[2\] _04160_ _04155_ _04161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10390_ _00263_ clknet_leaf_51_wb_clk_i cpu.uart.data_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09049_ _04085_ _04105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_102_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09340__A2 _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08864__I _03898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08851__A1 cpu.timer_capture\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10657_ _00529_ clknet_leaf_60_wb_clk_i net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_82_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10588_ _00460_ clknet_leaf_79_wb_clk_i cpu.last_addr\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07590__A1 _02964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06750_ _00771_ _00900_ _02215_ _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_116_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05701_ _01174_ _01048_ _01175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06681_ _02146_ _02145_ _02147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08420_ _03609_ _03616_ _00290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05632_ _01105_ _01092_ _01097_ _00821_ _01106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08774__I _03875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08351_ _03556_ _03562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05563_ _01014_ _01036_ _01037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09095__A1 _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08282_ _03510_ _03511_ _00257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07302_ _02733_ _02715_ _02716_ _02735_ _02736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05494_ _00842_ _00969_ _00970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07233_ cpu.uart.divisor\[0\] _02677_ _02678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_93_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_93_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_6_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05200__S0 _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_22_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_22_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_42_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07164_ _02333_ _02360_ _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06115_ _01306_ _01587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07095_ _01133_ _02541_ _02553_ _02547_ _02554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_2_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06081__A1 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06046_ _01517_ _01518_ _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09805_ _02484_ _04788_ _04789_ _04791_ _04792_ _00499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_07997_ _03280_ _03282_ _03284_ _00199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_66_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06384__A2 _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09736_ _04693_ _04734_ _04694_ _04735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06948_ _02398_ _02414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09667_ _04668_ _00485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_96_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07333__A1 _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08618_ _03749_ _03752_ _03762_ _03771_ _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_06879_ _00710_ _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_84_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09598_ _03136_ _04443_ _04602_ _04476_ _04603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08549_ _03711_ _00622_ _00324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05895__A1 _01310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07636__A2 _03000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10511_ _00384_ clknet_leaf_23_wb_clk_i cpu.timer\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05647__A1 _01120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10442_ _00315_ clknet_leaf_84_wb_clk_i cpu.orig_PC\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10373_ _00246_ clknet_leaf_32_wb_clk_i cpu.uart.div_counter\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05186__I0 cpu.regs\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05886__A1 _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05886__C _01359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07920_ cpu.timer\[13\] _03209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__05810__A1 _00984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09552__A2 _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07851_ _03132_ _03149_ _03115_ _03150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput2 io_in[10] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06802_ _00709_ _00943_ _02268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07782_ _03049_ _03092_ _03094_ _00174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09521_ _04507_ _04528_ _00479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06733_ _02150_ _02198_ _02162_ _02163_ _02199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_TAPCELL_ROW_108_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07315__A1 _02745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09452_ _02604_ _01778_ _04461_ _04462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06664_ _01825_ _02105_ _02128_ _02129_ _02130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_08403_ cpu.uart.receive_div_counter\[7\] _03581_ _03602_ _03583_ _03603_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05615_ _01061_ _01087_ _01088_ _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09383_ _01591_ _04388_ _04393_ _04394_ _04395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06595_ _02020_ _02061_ _02062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__05877__A1 _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08334_ cpu.uart.data_buff\[8\] _03528_ _03550_ _03551_ _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05546_ cpu.IO_addr_buff\[1\] _01020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08265_ _03438_ _03497_ _03441_ _03498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_74_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05477_ _00908_ _00952_ _00954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08196_ _03437_ _03443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07216_ _02560_ _02663_ _02664_ _02575_ _00038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09240__A1 _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07147_ _01101_ _02100_ _02600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07078_ _02537_ _02538_ _02539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_4
XTAP_TAPCELL_ROW_72_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06029_ _01346_ _01497_ _01501_ _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07583__I _01405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09543__A2 _04534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09719_ cpu.last_addr\[5\] _04698_ _04719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_6_0_wb_clk_i clknet_0_wb_clk_i clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_2_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_83_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06293__A1 cpu.timer_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08034__A2 _03262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10425_ _00298_ clknet_leaf_55_wb_clk_i cpu.orig_IO_addr_buff\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09231__A1 _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_17_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10356_ _00229_ clknet_leaf_43_wb_clk_i cpu.uart.dout\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07793__A1 cpu.regs\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10287_ _00160_ clknet_leaf_106_wb_clk_i cpu.regs\[6\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_29_Left_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07545__A1 _01407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_1_Left_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_56_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05400_ _00878_ _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_38_Left_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06380_ _01834_ _01847_ _01848_ _01849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_28_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05331_ cpu.PORTA_DDR\[5\] net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_16_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08050_ cpu.spi.data_out_buff\[4\] _03314_ _03324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05087__A2 net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05262_ _00762_ _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07001_ _02453_ _02459_ _02464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05193_ _00694_ _00697_ _00698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06587__A2 _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_47_Left_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08952_ _02779_ _04027_ _04029_ _00409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08499__I _03662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07903_ cpu.timer_div\[1\] _03185_ _03186_ cpu.timer_div\[5\] _03191_ _03192_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_08883_ _03209_ _03970_ _03975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10043__B _02683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07834_ _02429_ _02368_ _03133_ _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_79_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09289__A1 _01309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07765_ _03072_ _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_69_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09504_ _04238_ _04510_ _04511_ _04512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06716_ _02179_ _02181_ _02182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07696_ _02987_ _03036_ _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06647_ _02112_ _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XPHY_EDGE_ROW_56_Left_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09435_ _04443_ _04445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05651__I _01051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06511__A2 _01230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06578_ _01086_ _02044_ _02045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09366_ _04377_ _04378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05529_ _00993_ _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08317_ _02806_ _03521_ _03525_ _03537_ _03538_ _00265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_09297_ _04082_ _04308_ _04310_ _04311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09279__B _00593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08248_ _03396_ _03480_ _03484_ _03479_ _00250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08179_ _03423_ _03428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_65_Left_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10210_ _00083_ clknet_leaf_3_wb_clk_i _00001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07775__A1 cpu.regs\[4\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10141_ _00018_ clknet_leaf_117_wb_clk_i cpu.regs\[9\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10072_ _05002_ _05003_ _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_7_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_74_Left_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09033__I _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_qcpu_113 io_oeb[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xwrapped_qcpu_102 io_oeb[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_85_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06502__A2 _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07488__I cpu.uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10408_ _00281_ clknet_leaf_37_wb_clk_i cpu.uart.receive_div_counter\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10339_ _00212_ clknet_leaf_63_wb_clk_i cpu.spi.data_out_buff\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07230__A3 _02674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05880_ _01339_ _00858_ _01354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_105_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08268__B _03464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07550_ cpu.regs\[14\]\[3\] _02940_ _02944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06501_ net32 _01096_ _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07481_ cpu.uart.receive_div_counter\[9\] _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08494__A2 _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09220_ _04236_ _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06432_ _01871_ _01412_ _01900_ _01277_ _01901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_29_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09151_ _04185_ _00452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_60_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06363_ _00785_ _01832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_32_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08102_ _03351_ _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07398__I _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09082_ cpu.orig_IO_addr_buff\[6\] _04090_ _04133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05314_ _00779_ _00811_ _00812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10038__B net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08033_ _00624_ _01424_ _03310_ _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06294_ _01762_ _01763_ _01764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_25_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06009__A1 _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05245_ _00732_ _00746_ _00682_ _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_116_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05176_ _00681_ cpu.ROM_spi_mode net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_12_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09984_ _04928_ _04930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08935_ _04004_ _02755_ _04005_ _04017_ _04018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_4_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input21_I io_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08866_ _03207_ _03954_ _03961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08797_ _03901_ _03902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07817_ _01330_ _01404_ _03118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06732__A2 _02009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07748_ _03072_ _03073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07679_ _02971_ _03022_ _03026_ _00139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_109_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09418_ _04390_ _04415_ _04428_ _04392_ _04429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_10690_ _00562_ clknet_leaf_4_wb_clk_i cpu.regs\[15\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09349_ _04361_ _04362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08788__A3 _02763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_91_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10124_ cpu.regs\[15\]\[3\] _05045_ _05049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10055_ _04755_ _04751_ _04987_ _04760_ _04988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XPHY_EDGE_ROW_82_Left_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06487__A1 _01952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08535__C _03695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_91_Left_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06411__A1 _01877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06981_ _02427_ _02428_ _02445_ _02417_ _02446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_111_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_47_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_47_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08720_ _02800_ _03843_ _03848_ _03846_ _00358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05932_ _01405_ _01406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08164__A1 _03262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08651_ _03796_ _03799_ _03800_ _00337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05863_ _01336_ _01337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__05517__A3 _00609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07602_ _02967_ _02979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_37_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05794_ _01049_ _01268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08582_ cpu.toggle_ctr\[12\] _01738_ _03729_ cpu.toggle_ctr\[11\] _03736_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07533_ net15 _02931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_66_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06478__A1 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07464_ _02857_ _02824_ _02869_ _00081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06415_ _01883_ _01193_ _01191_ _01884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09203_ _04215_ _04224_ _04225_ _00464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_76_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09134_ _04172_ _00448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07395_ _02745_ _02811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_17_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06346_ _01723_ _01797_ _01802_ _01816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06277_ net10 _01226_ _01555_ _01747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_72_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09065_ _00926_ _04105_ _04118_ _04119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08016_ cpu.spi.div_counter\[6\] _03295_ _03297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05228_ _00722_ _00730_ _00731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_77_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09276__C _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05159_ _00666_ _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05376__I _00855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09967_ _04917_ _00536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08918_ _01456_ _04004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09898_ _00611_ _02536_ _04868_ _04869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__07591__I _01541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07902__A1 cpu.timer_div\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08849_ _03180_ _03947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05508__A3 _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08458__A2 _03643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10673_ _00545_ clknet_leaf_86_wb_clk_i cpu.PORTA_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05141__A1 _00647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07969__A1 _00613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05286__I _00785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05219__C _00707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10107_ _04454_ _05036_ _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10038_ _04955_ _02511_ net76 _04972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06200_ _01419_ _01669_ _01670_ _01671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_73_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06880__A1 _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07180_ _02107_ _02584_ _02631_ _02632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06131_ _01601_ _01602_ _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06062_ _01526_ _01533_ _01535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_113_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09821_ _04804_ _04807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09752_ _02562_ _04747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08703_ _03834_ _03835_ _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06964_ _02426_ _02429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09683_ _04434_ _04674_ _04683_ _04341_ _04684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_05915_ _00589_ _01382_ _01389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06895_ _02333_ _02360_ _02361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05846_ _01030_ _01320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08634_ _03182_ _03786_ _03787_ _03788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_89_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05777_ _01250_ _01037_ _01251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09637__A1 _04362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08565_ cpu.toggle_top\[4\] _03722_ _03723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07516_ _00664_ _02875_ _02916_ _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_76_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08496_ _00614_ _03674_ _03663_ _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07447_ _02824_ _02853_ _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_91_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07378_ _00979_ _02796_ _02798_ _02799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06871__A1 _00726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09117_ _00727_ _02859_ _04153_ _04160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06329_ _01796_ _01798_ _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09048_ _04081_ _04097_ _04104_ _00430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06623__A1 _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05834__I cpu.C vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09628__A1 _03703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09041__I _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06665__I net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10656_ _00528_ clknet_leaf_60_wb_clk_i net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05665__A2 _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10587_ _00459_ clknet_leaf_74_wb_clk_i cpu.last_addr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06614__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_10_Left_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_2_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05700_ _01047_ _01174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06680_ cpu.regs\[1\]\[1\] _02008_ _02146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05631_ _01104_ _01105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08350_ _03561_ _00275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_63_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09619__A1 _03701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05562_ _01030_ _01035_ _01036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07301_ _02734_ _02718_ _02735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08281_ _03507_ _03409_ _00239_ _03511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05493_ cpu.regs\[0\]\[5\] cpu.regs\[1\]\[5\] cpu.regs\[2\]\[5\] cpu.regs\[3\]\[5\]
+ _00829_ _00891_ _00969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_18_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07232_ _02675_ _02677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06853__A1 _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07163_ net12 _02593_ _02429_ _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06114_ _01584_ _01291_ _01585_ _01586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06605__A1 _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07339__C _02683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07094_ _02542_ _02552_ _02553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_62_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_62_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_100_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06081__A2 _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06045_ _00820_ _00821_ _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_112_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09804_ _02872_ _04792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_5_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07996_ cpu.spi.div_counter\[0\] _03164_ _03283_ _03284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09735_ _04733_ _02561_ _04734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07581__A2 _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06947_ _02398_ _02412_ _02413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09666_ _02414_ _04443_ _04667_ _04411_ _04668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10212__D _00085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08530__A1 _03136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08617_ _03766_ _03767_ _03768_ _03770_ _03771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_06878_ _02334_ _02343_ _02344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_09597_ _04478_ _04580_ _04582_ _04408_ _04601_ _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05829_ _00874_ _01302_ _01303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05195__I1 cpu.regs\[9\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08548_ cpu.toggle_clkdiv _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_25_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08479_ _03662_ _03663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10510_ _00383_ clknet_leaf_23_wb_clk_i cpu.timer\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05647__A2 _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10441_ _00314_ clknet_leaf_83_wb_clk_i cpu.orig_PC\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10372_ _00245_ clknet_leaf_32_wb_clk_i cpu.uart.div_counter\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06072__A2 _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05564__I _00993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_88_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05186__I1 _00689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_46_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10639_ _00511_ clknet_leaf_65_wb_clk_i cpu.ROM_spi_cycle\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07850_ net19 _03121_ _03145_ _03148_ _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA_clkbuf_leaf_85_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05413__I2 cpu.regs\[10\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06801_ _00709_ _00949_ _02267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07781_ cpu.regs\[4\]\[4\] _03093_ _03094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput3 io_in[11] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09520_ _04367_ _04524_ _04525_ _04527_ _04528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06732_ _00762_ _02009_ _02198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_108_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06519__B _01986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09451_ _04459_ _04419_ _04460_ _04461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06663_ cpu.regs\[2\]\[4\] _02129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08402_ _03601_ _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_93_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05614_ _00596_ _00649_ _01088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09382_ _04355_ _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06594_ _01312_ _01313_ _02059_ _02060_ _02061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_19_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05877__A2 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08333_ _03181_ _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_86_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05545_ _00995_ _01019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06238__C _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08264_ _03378_ _03493_ _03488_ _03489_ _03497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_62_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06826__A1 _00689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05476_ _00908_ _00952_ _00953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08195_ _03383_ _03438_ _03441_ _03442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_61_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07215_ _01779_ _02662_ _02664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_14_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07146_ _02591_ _02598_ _02599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07077_ _00626_ _00674_ _02538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_30_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06028_ _01345_ _01500_ _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07554__A2 _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07979_ cpu.spi.div_counter\[7\] cpu.spi.divisor\[7\] _03267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09718_ _04714_ _04716_ _04717_ _04718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_58_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08503__A1 _02848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09649_ cpu.regs\[2\]\[4\] _04403_ _04650_ _04651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05317__A1 _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10424_ _00297_ clknet_leaf_54_wb_clk_i cpu.orig_IO_addr_buff\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08034__A3 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06045__A2 _00821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10355_ _00228_ clknet_leaf_43_wb_clk_i cpu.uart.dout\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08990__A1 cpu.timer_div\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10129__A1 _01826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10286_ _00159_ clknet_leaf_106_wb_clk_i cpu.regs\[6\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_2_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08538__C _03695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05330_ cpu.PORTB_DDR\[5\] net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_7_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05087__A3 _00595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05261_ _00761_ _00762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05469__I _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05192_ cpu.regs\[12\]\[0\] cpu.regs\[13\]\[0\] cpu.regs\[14\]\[0\] cpu.regs\[15\]\[0\]
+ _00695_ _00696_ _00697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_07000_ cpu.regs\[2\]\[7\] _02128_ _02463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07233__A1 cpu.uart.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08951_ cpu.spi.divisor\[4\] _04028_ _04029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_102_Left_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08981__A1 cpu.timer_div\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07902_ cpu.timer_div\[5\] _03186_ cpu.timer_div_counter\[7\] _03187_ _03190_ _03191_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08882_ _03624_ _03974_ _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05418__B _00853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07833_ _02290_ _02366_ _02367_ _03133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XPHY_EDGE_ROW_81_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_55_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05932__I _01405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07764_ _03053_ _03074_ _03082_ _00168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09503_ cpu.orig_PC\[6\] _04374_ _04511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06715_ _02137_ _02180_ _02181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07695_ _01117_ _03035_ _03036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_94_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06646_ cpu.mem_cycle\[2\] _02112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_69_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09434_ _04438_ _04442_ _04444_ _00476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_111_Left_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06577_ cpu.timer_capture\[15\] _01255_ _02044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09365_ _04304_ _04377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05528_ _01001_ _01002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08316_ cpu.uart.data_buff\[4\] _03531_ _03538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09296_ cpu.orig_PC\[0\] _04099_ _04309_ _01288_ _04310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_47_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08247_ cpu.uart.div_counter\[10\] _03441_ _03483_ _03438_ _03484_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_90_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05459_ cpu.regs\[8\]\[4\] cpu.regs\[9\]\[4\] cpu.regs\[10\]\[4\] cpu.regs\[11\]\[4\]
+ _00932_ _00935_ _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__05379__I _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08178_ _02794_ _03427_ _00236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07129_ _02581_ _02113_ _02582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__07594__I _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08972__A1 _01546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10140_ _00017_ clknet_leaf_117_wb_clk_i cpu.regs\[9\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10071_ _04958_ _04950_ _05003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05538__A1 _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_qcpu_114 io_oeb[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xwrapped_qcpu_103 io_oeb[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_84_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09452__A2 _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06266__A2 _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09984__I _04928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09204__A2 _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07215__A1 _01779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10407_ _00280_ clknet_leaf_39_wb_clk_i cpu.uart.receive_div_counter\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10338_ _00211_ clknet_leaf_61_wb_clk_i cpu.spi.data_out_buff\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_119_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_119_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07009__I net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10269_ _00142_ clknet_leaf_118_wb_clk_i cpu.regs\[8\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_105_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07480_ cpu.uart.receive_div_counter\[5\] _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_88_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06500_ _01944_ _01958_ _01967_ net96 _01491_ _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XANTENNA__09691__A2 _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05701__A1 _01174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06431_ _01872_ _01417_ _01418_ _01899_ _01900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_90_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09150_ cpu.ROM_addr_buff\[10\] _04184_ _04181_ _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06362_ _01830_ _01137_ _01831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08101_ cpu.uart.receive_buff\[3\] _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06293_ cpu.timer_top\[4\] _01459_ _01264_ _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09081_ _04122_ _04131_ _04132_ _00435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05313_ cpu.regs\[8\]\[7\] cpu.regs\[9\]\[7\] cpu.regs\[10\]\[7\] cpu.regs\[11\]\[7\]
+ _00788_ _00789_ _00811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08032_ _02672_ _03310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_71_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05199__I _00703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05244_ cpu.regs\[4\]\[3\] cpu.regs\[5\]\[3\] cpu.regs\[6\]\[3\] cpu.regs\[7\]\[3\]
+ _00733_ _00734_ _00746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_32_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05175_ cpu.ROM_OEB _00681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07206__A1 _02654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08954__A1 _02784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09983_ _04928_ _04929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05148__B _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08934_ cpu.timer\[15\] _04006_ _04017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08865_ cpu.timer\[11\] _03960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08796_ _03898_ _03901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07816_ _00690_ _03116_ _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input14_I io_in[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07747_ _03071_ _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07678_ cpu.regs\[8\]\[1\] _03025_ _03026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09417_ _02860_ _04427_ _04428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06629_ _01403_ _02095_ _02096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09348_ _02762_ _04339_ _04361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07996__A2 _03164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09279_ _01372_ _01336_ _00593_ _04293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_90_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output82_I net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07257__C _02697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10123_ _01643_ _05044_ _05048_ _00561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10054_ _04753_ _02502_ _04754_ _04943_ _02482_ _04987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06184__A1 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_7_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07987__A2 cpu.spi.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09219__I _04087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08936__A1 cpu.timer_capture\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07739__A2 _03058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06980_ _02429_ _02444_ _02445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input6_I io_in[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05931_ _01330_ _01404_ _01405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08164__A2 _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08650_ cpu.toggle_ctr\[4\] _03797_ _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05862_ _01335_ _01336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_89_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07601_ _02967_ _02978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_37_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_87_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_87_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09113__A1 _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05793_ cpu.timer_top\[8\] _01170_ _01177_ _01266_ _01267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_49_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08581_ cpu.toggle_ctr\[14\] _03734_ _01871_ cpu.toggle_ctr\[13\] _03735_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07532_ cpu.uart.receive_counter\[2\] _02926_ _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08793__I _03898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_16_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_16_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_49_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07463_ _02858_ _02603_ _02868_ _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06414_ cpu.uart.divisor\[13\] _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09202_ cpu.ROM_addr_buff\[8\] _04220_ _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09133_ cpu.ROM_addr_buff\[6\] _04171_ _04169_ _04172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07394_ _02695_ _02801_ _02808_ _02810_ _00070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_8_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06345_ _01723_ _01802_ _01797_ _01815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06276_ net2 _01221_ _01745_ _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09064_ cpu.orig_IO_addr_buff\[3\] _04106_ _04118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08015_ _03280_ _03296_ _00205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_102_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05227_ _00694_ _00723_ _00729_ _00682_ _00730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_05158_ _00665_ _00666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_77_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08927__A1 cpu.timer_capture\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09966_ cpu.PORTB_DDR\[3\] _04907_ _04915_ _04916_ _04917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05089_ cpu.IO_addr_buff\[7\] cpu.IO_addr_buff\[6\] cpu.IO_addr_buff\[5\] _00600_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_09897_ _00673_ _00674_ _04867_ _00990_ _04868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08917_ _03985_ _04003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08848_ _03895_ _03945_ _03946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08779_ _02784_ _03883_ _03887_ _03886_ _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_67_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10672_ _00544_ clknet_leaf_59_wb_clk_i cpu.PORTA_DDR\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08208__I _03440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09039__I _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10106_ _05023_ _05024_ _05035_ _05036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10037_ _04957_ _04970_ _04971_ _03421_ _00552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08099__B _00679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09343__A1 _00989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05380__A2 _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08449__A3 _03638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06130_ _01120_ net92 _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06061_ _01526_ _01533_ _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_113_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08909__A1 _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09820_ _04805_ _04806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09751_ _04742_ _04746_ _02710_ _00491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05443__I0 cpu.regs\[0\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06963_ cpu.PC\[13\] _02413_ _02428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08702_ cpu.pwm_counter\[5\] _03832_ _03709_ _03835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05914_ _00907_ _01385_ _01387_ _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09682_ _04294_ _04676_ _04682_ _04386_ _04683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06894_ _02335_ _02343_ _02344_ _02357_ _02359_ _02360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_05845_ _01025_ _01016_ _01319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08633_ _03711_ _03751_ _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05776_ _01004_ _01250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08564_ _03713_ _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07515_ _02915_ _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_76_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08495_ _03658_ _03674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06257__B _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07446_ _02626_ _02849_ _02852_ _02589_ _02853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_45_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07377_ _01275_ _02797_ _02798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_79_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09116_ _04159_ _00443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06328_ _01396_ _01784_ _01797_ _01615_ _01798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_103_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09047_ _00568_ _04098_ _04103_ _04104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_20_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06259_ _01375_ _01725_ _01729_ _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05682__I0 cpu.regs\[12\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09949_ _04111_ _04904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09325__A1 cpu.uart.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06011__I cpu.Z vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_36_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08366__C _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09628__A2 _00880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10655_ _00527_ clknet_leaf_61_wb_clk_i net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_82_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10586_ _00458_ clknet_leaf_74_wb_clk_i cpu.last_addr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06630__B _02062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05630_ cpu.br_rel_dest\[0\] _01104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09619__A2 _04554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06077__B cpu.PORTA_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05561_ _00603_ _00996_ _01035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07300_ cpu.timer\[3\] _02734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_63_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08280_ _03508_ _03509_ _03510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05105__A2 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05492_ _00909_ _00967_ _00847_ _00968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_117_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07231_ _02675_ _02676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06853__A2 _00855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08055__A1 _02784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07162_ _02602_ _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_42_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06113_ _01513_ _01585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07093_ net19 _02543_ _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_42_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07802__A1 cpu.regs\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09835__C _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06044_ _00906_ _01340_ _01517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_74_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09803_ _02484_ _04790_ _04791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07995_ _03262_ _03264_ _03283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09734_ _02489_ _04733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_31_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_31_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06946_ _02411_ _02412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09665_ _04478_ _04649_ _04651_ _04408_ _04666_ _04667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06877_ _02312_ _02336_ _02339_ _02342_ _02343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_08616_ _03753_ _01872_ _01167_ _03751_ _03769_ _03770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_05828_ _01301_ _01302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_96_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09596_ _04326_ _04600_ _04601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08547_ _03432_ _03635_ _00323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05759_ cpu.uart.divisor\[8\] _01194_ _01200_ _01232_ _01233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08478_ _00677_ _03662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07429_ cpu.PC\[1\] _02837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10440_ _00313_ clknet_leaf_83_wb_clk_i cpu.orig_PC\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07597__I _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10371_ _00244_ clknet_leaf_28_wb_clk_i cpu.uart.div_counter\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09546__A1 _04529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08221__I _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06780__A1 _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05186__I2 _00690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10638_ _00510_ clknet_leaf_65_wb_clk_i cpu.ROM_spi_cycle\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10569_ _00441_ clknet_leaf_97_wb_clk_i cpu.base_address\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07456__B _02861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06800_ _02260_ _02261_ _02250_ _02266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_07780_ _03085_ _03093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10313__D _00186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput4 io_in[12] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06731_ _02195_ _02196_ _02197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_108_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09450_ _02402_ _01112_ _04460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08401_ cpu.uart.receive_div_counter\[7\] _03600_ _03601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06662_ _02104_ _02127_ _02128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05613_ _01065_ _01087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09381_ _04094_ _04370_ _04391_ _04392_ _04393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06593_ _01089_ _02021_ _02060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08332_ _02790_ _03540_ _03549_ _03550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05544_ _01012_ _01017_ _01018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08263_ _03494_ _03490_ _03496_ _03479_ _00253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_52_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05475_ _00951_ _00952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_07214_ _02662_ _02663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08194_ _03440_ _03441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07145_ _02593_ _02595_ _02597_ _02598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_112_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07076_ _00627_ _02536_ _02537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_30_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06027_ _01498_ _01499_ _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_30_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08200__A1 _03391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07978_ cpu.spi.div_counter\[6\] cpu.spi.divisor\[6\] _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09717_ cpu.last_addr\[4\] cpu.ROM_addr_buff\[4\] _04697_ _04717_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_58_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06929_ _02212_ _02372_ _02394_ _02395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09648_ _04404_ _04649_ _04650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_2_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09579_ _04498_ _04580_ _04583_ _04584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_108_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10423_ _00296_ clknet_leaf_48_wb_clk_i cpu.needs_interrupt vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10354_ _00227_ clknet_leaf_43_wb_clk_i cpu.uart.dout\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09519__A1 _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10285_ _00158_ clknet_4_2_0_wb_clk_i cpu.regs\[6\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06505__A1 cpu.PORTB_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08835__B _03894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05260_ cpu.regs\[1\]\[4\] _00761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05191_ _00001_ _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_51_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08950_ _04020_ _04028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_71_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05485__I _00960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07901_ cpu.timer_div\[0\] _03188_ cpu.timer_div_counter\[2\] _01546_ _03189_ _03190_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_08881_ cpu.timer_capture\[13\] _03930_ _03973_ _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08796__I _03898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07832_ _02935_ _02601_ _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09502_ _04509_ _04510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07763_ cpu.regs\[5\]\[6\] _03072_ _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_79_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_55_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06714_ _00761_ _00943_ _02180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07694_ _01124_ _02936_ _03035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06645_ _02110_ _02111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_69_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09433_ _02861_ _04443_ _04444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09364_ _04238_ _04371_ _04375_ _04376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08315_ cpu.uart.data_buff\[5\] _03537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06576_ _02041_ _02042_ _02043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_35_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05527_ _00569_ _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09295_ _02829_ _04099_ _04309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08246_ _03396_ _03480_ _03483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05458_ _00833_ _00935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08177_ _03425_ _03418_ _03426_ _03417_ _03427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07128_ _02110_ _02581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_70_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08480__B _03663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05389_ _00862_ _00864_ _00866_ _00868_ _00869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_113_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07059_ cpu.ROM_addr_buff\[11\] _02521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05395__I _00874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06983__A1 _01921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10070_ _04760_ _05000_ _05001_ _05002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_7_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_102_Right_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09921__A1 _02701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_qcpu_115 io_oeb[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xwrapped_qcpu_104 io_oeb[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__07115__I _02549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09988__A1 cpu.PORTA_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08390__B _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10406_ _00279_ clknet_leaf_39_wb_clk_i cpu.uart.receive_buff\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10337_ _00210_ clknet_leaf_61_wb_clk_i cpu.spi.data_out_buff\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08963__A2 _00979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10268_ _00141_ clknet_leaf_120_wb_clk_i cpu.regs\[8\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09912__A1 _02690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10199_ _00010_ clknet_leaf_86_wb_clk_i cpu.instr_cycle\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_105_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09140__A2 cpu.regs\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06430_ _01896_ _01897_ _01898_ _01899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09979__A1 _02790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06361_ _01829_ _01830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_32_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08100_ _03357_ _03352_ _03359_ _00227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_83_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06292_ cpu.timer_capture\[12\] _01460_ _01761_ _01464_ _01762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09080_ cpu.IO_addr_buff\[5\] _03446_ _04127_ _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_60_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05312_ _00808_ _00809_ _00787_ _00810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_114_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08031_ _03308_ _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05243_ _00737_ _00744_ _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05174_ _00629_ _00675_ _00680_ _00009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09982_ _01033_ _03712_ _04928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_40_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08933_ _04016_ _00403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_4_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08864_ _03898_ _03959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06193__A2 _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08795_ _03893_ _03896_ _03900_ _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07390__A1 _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07815_ _03115_ _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05164__B _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07746_ _02600_ _03036_ _03071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_79_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08475__B _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09416_ _04426_ _04427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07677_ _03020_ _03025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06628_ _02075_ _02090_ _02094_ net97 _01638_ _02095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_06559_ _02025_ _01202_ _00999_ _02026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09347_ _04326_ _04333_ _04358_ _04359_ _04360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09278_ _04243_ _04292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08229_ _03443_ _03470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output75_I net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_91_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10122_ cpu.regs\[15\]\[2\] _05045_ _05048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10053_ _04980_ _04985_ _04731_ _04986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09370__A2 _01120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06184__A2 _01221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05931__A2 _01404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08881__A1 cpu.timer_capture\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09995__I _04928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06947__A1 _02398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09897__B1 _04867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05930_ net26 _01334_ _01402_ _01403_ _01404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_05861_ _00641_ _01335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08580_ cpu.toggle_top\[14\] _03734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07600_ _01826_ _02977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_37_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07531_ cpu.uart.receive_counter\[2\] _02926_ _02929_ _00088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05792_ _01253_ _01259_ _01265_ _01266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_66_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07462_ _02589_ _02867_ _02827_ _02868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06413_ _01881_ _01428_ _01659_ _01882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09201_ cpu.last_addr\[8\] _04216_ _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07393_ _02809_ _02810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_45_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_56_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_56_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09132_ cpu.regs\[2\]\[6\] _02637_ _04167_ _04171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06344_ _01800_ _01788_ _01804_ _01625_ _01813_ _01814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_72_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06275_ _01228_ _01745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09063_ _04081_ _04116_ _04117_ _00432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08014_ cpu.spi.div_counter\[6\] _03295_ _03296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_4_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05226_ _00692_ _00728_ _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05157_ _00664_ _00665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_77_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09965_ _04111_ _04916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05088_ cpu.IO_addr_buff\[4\] _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08916_ _04002_ _00400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05673__I _00595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09896_ _01331_ _01133_ _04867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__05461__I1 cpu.regs\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08847_ _03943_ _03859_ _03891_ _03944_ _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07363__A1 _02784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_26_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08778_ cpu.timer_top\[13\] _03884_ _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07729_ _03034_ _03059_ _03061_ _00154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10671_ _00543_ clknet_leaf_59_wb_clk_i cpu.PORTA_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05677__A1 _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09040__B2 _01105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_65_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10105_ _01834_ _05027_ _05028_ _05034_ _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_10036_ net72 _04957_ _04971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09055__I _00677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06060_ _01309_ _01353_ _01351_ _01533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07593__A1 _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_103_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_103_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09750_ _04744_ _04745_ _04746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05443__I1 cpu.regs\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06962_ _02426_ _02427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09681_ _04416_ _04680_ _04681_ _04682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08701_ cpu.pwm_counter\[5\] _03832_ _03834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05913_ _01373_ _01386_ _01387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07345__A1 _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08632_ _03711_ _03785_ _03786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_06893_ _02344_ _02358_ _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05844_ _01229_ _01279_ _01063_ _01296_ _01318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_05775_ cpu.timer_capture\[0\] _01248_ _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08563_ _03713_ _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07514_ _02879_ _02884_ _02897_ _02914_ _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_89_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08494_ cpu.orig_flags\[3\] _03672_ _03673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07213__I _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07445_ _02427_ _02851_ _02852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07376_ _02795_ _02797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09115_ cpu.ROM_addr_buff\[1\] _04158_ _04155_ _04159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09270__A1 _01830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06327_ _01785_ _01797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_17_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09046_ _04102_ _04103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05668__I _01141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06258_ _01715_ _01727_ _01728_ _01729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05209_ cpu.regs\[0\]\[1\] _00710_ cpu.regs\[2\]\[1\] cpu.regs\[3\]\[1\] _00711_
+ _00712_ _00713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_06189_ _01658_ _01428_ _01659_ _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08979__I _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09948_ _02790_ _04895_ _04903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09325__A2 cpu.spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09879_ net74 _03786_ _04852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09089__A1 _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output38_I net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08836__A1 cpu.timer_capture\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10654_ _00526_ clknet_leaf_60_wb_clk_i net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_82_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10585_ _00457_ clknet_leaf_74_wb_clk_i cpu.last_addr\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09261__A1 _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_1_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_1_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_101_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10019_ _00608_ _04763_ _02472_ _04955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_47_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05433__S0 _00828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05889__A1 _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05560_ _01019_ _01023_ _01028_ _01033_ _01034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_59_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06550__A2 _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08827__A1 _03259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05491_ cpu.regs\[12\]\[5\] cpu.regs\[13\]\[5\] cpu.regs\[14\]\[5\] cpu.regs\[15\]\[5\]
+ _00918_ _00834_ _00967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_07230_ _01005_ _01023_ _02674_ _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_82_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09252__A1 _00951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07161_ _01920_ _02612_ _02613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06112_ _01089_ _01584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07092_ _02551_ _00027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09004__A1 _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08799__I _03898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06043_ _01511_ _01512_ _01514_ _01515_ _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_22_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09802_ _02513_ _04790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07566__A1 _01407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07994_ _03261_ _03265_ _03281_ _03282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_66_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09851__C _04792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09733_ _04732_ _00487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06112__I _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06945_ cpu.PC\[11\] _02410_ _02411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09664_ _04326_ _04665_ _04666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06876_ _02314_ _02341_ _02342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09595_ _04455_ _04580_ _04599_ _04502_ _04600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08615_ _03765_ _03764_ _03769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05827_ _01296_ _01284_ _01301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_71_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_71_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_82_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05758_ _01222_ _01227_ _01231_ _01232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_85_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08546_ _03707_ _03710_ _00322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_92_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08483__B _03663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08477_ cpu.orig_IO_addr_buff\[6\] _03655_ _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05689_ _01160_ _01162_ _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_25_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07428_ _02340_ _02824_ _02836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07359_ _02012_ _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_80_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09243__A1 _01822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10370_ _00243_ clknet_leaf_29_wb_clk_i cpu.uart.div_counter\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09029_ _04085_ _04086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07557__A1 _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06780__A2 _00873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06957__I _02104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05861__I _00641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05415__S0 _00830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05186__I3 cpu.regs\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10637_ _00509_ clknet_leaf_67_wb_clk_i cpu.ROM_spi_cycle\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_116_Right_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07796__A1 cpu.regs\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10568_ _00440_ clknet_leaf_97_wb_clk_i cpu.base_address\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10499_ _00372_ clknet_leaf_28_wb_clk_i cpu.timer_div_counter\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput5 io_in[13] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06730_ _02165_ _02167_ _02196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_108_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06661_ _02122_ _02126_ _02127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_36_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08400_ _03599_ _02881_ _03590_ _03600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_05612_ _01040_ _01085_ _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_59_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09380_ _04351_ _04392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06592_ _01392_ _01474_ _01584_ _02058_ _02059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05543_ _01013_ _01016_ _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08331_ cpu.uart.data_buff\[9\] _03539_ _03549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08262_ _03493_ _03441_ _03495_ _03438_ _03496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_6_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05474_ _00950_ _00951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_22_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07698__I _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07213_ _02661_ _02662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08193_ _03411_ _03439_ _03440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_61_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06039__A1 _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07144_ net1 _02596_ _02597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07075_ _00576_ _00615_ _00655_ _02536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_42_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09528__A2 _04534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06026_ _01487_ _00717_ _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07977_ _03262_ _03264_ _03265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06211__A1 _01680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09716_ cpu.last_addr\[3\] cpu.ROM_addr_buff\[3\] _04715_ _04716_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_58_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06928_ _02373_ _02393_ _02394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09647_ _04648_ _04649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_2_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06859_ _02320_ _02324_ _02325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09578_ cpu.orig_PC\[9\] _04088_ _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08529_ cpu.orig_PC\[9\] _03684_ _03698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09464__A1 _04454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06278__A1 _01744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07401__I _02755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10422_ _00295_ clknet_leaf_33_wb_clk_i cpu.uart.receive_div_counter\[15\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10353_ _00226_ clknet_leaf_42_wb_clk_i cpu.uart.dout\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09328__I _04340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06450__A1 _00946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10284_ _00157_ clknet_leaf_2_wb_clk_i cpu.regs\[6\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09772__B _02683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06202__A1 cpu.timer_capture\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06753__A2 _00973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06505__A2 _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10065__A2 _04731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06636__B _01926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05190_ _00000_ _00695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_24_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07900_ cpu.timer_div\[0\] _03188_ _03185_ cpu.timer_div\[1\] _03189_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08880_ _03209_ _03918_ _03894_ _03972_ _03973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07831_ _03130_ _03119_ _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_16_Left_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09501_ _02636_ _04508_ _04509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07762_ _03051_ _03074_ _03081_ _00167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06713_ _00798_ _00899_ _02179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07693_ _01405_ _03034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06644_ cpu.mem_cycle\[3\] _02110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09432_ _02531_ _04244_ _04443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_69_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06575_ cpu.timer_capture\[7\] _01419_ _01251_ _02042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09363_ cpu.orig_PC\[2\] _04374_ _04375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05526_ _00999_ _01000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_93_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08314_ _02804_ _03522_ _03526_ _03535_ _03536_ _00264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_35_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09294_ _04296_ _04301_ _04307_ _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_25_Left_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08245_ _02873_ _03481_ _03482_ _00249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05457_ _00909_ _00933_ _00934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08176_ _03425_ _03423_ _03426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06680__A1 cpu.regs\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05388_ _00843_ _00867_ _00853_ _00868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_27_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07127_ _02119_ _02580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07058_ _02501_ _02520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06009_ _00859_ _01481_ _01482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_7_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07891__I _00664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_34_Left_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07932__B2 cpu.timer_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07932__A1 cpu.timer_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08488__A2 _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_qcpu_105 io_oeb[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_EDGE_ROW_43_Left_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06671__A1 cpu.regs\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10405_ _00278_ clknet_leaf_38_wb_clk_i cpu.uart.receive_buff\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10336_ _00209_ clknet_leaf_61_wb_clk_i cpu.spi.data_out_buff\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_52_Left_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08897__I _01456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10267_ _00140_ clknet_leaf_119_wb_clk_i cpu.regs\[8\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10198_ _00009_ clknet_leaf_87_wb_clk_i cpu.instr_cycle\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_105_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_61_Left_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06360_ _00647_ _01829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06291_ _01759_ _01760_ _01761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_60_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05311_ cpu.regs\[4\]\[7\] cpu.regs\[5\]\[7\] cpu.regs\[6\]\[7\] cpu.regs\[7\]\[7\]
+ _00794_ _00795_ _00809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xinput30 sram_out[4] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08030_ _03307_ _03308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05242_ cpu.regs\[0\]\[3\] _00742_ _00743_ cpu.regs\[3\]\[3\] _00733_ _00734_ _00744_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06662__A1 _02104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_5_0_wb_clk_i clknet_0_wb_clk_i clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_05173_ cpu.instr_cycle\[1\] _00629_ _00679_ _00680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09600__A1 _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09981_ _04927_ _00540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_110_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08932_ cpu.timer_capture\[14\] _04003_ _04014_ _04015_ _04016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_4_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08863_ _03958_ _00391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_98_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08794_ cpu.timer_capture\[0\] _03899_ _03371_ _03900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07814_ _02422_ _02126_ _03114_ _03115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA_clkbuf_leaf_16_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07745_ _03014_ _03069_ _03070_ _00161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09415_ _01134_ _04426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07676_ _02964_ _03022_ _03024_ _00138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09419__A1 _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06627_ _01800_ _02070_ _02093_ _01629_ _02094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__10029__A2 _04963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06558_ net67 _02025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_81_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09346_ _03310_ _04325_ _04359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09277_ _04291_ _00472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05509_ cpu.instr_buff\[15\] _00983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06489_ _01132_ _01933_ _01946_ _01368_ _01956_ _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08228_ cpu.uart.div_counter\[6\] _03468_ _03469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08491__B _03663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08159_ _03412_ _03413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06405__A1 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_55_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10121_ _01542_ _05044_ _05047_ _00560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output68_I net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10052_ _02491_ _02500_ _04984_ _04985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08158__A1 _00676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07905__A1 _01546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07905__B2 cpu.timer_div\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08510__I _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09658__A1 _02398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08330__A1 _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07133__A2 _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_94_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10319_ _00192_ clknet_leaf_44_wb_clk_i cpu.spi.dout\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06947__A2 _02412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05860_ _01333_ _01334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05791_ cpu.timer_top\[0\] _01260_ _01264_ _01265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09649__A1 cpu.regs\[2\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07530_ _02922_ _02928_ cpu.uart.receive_counter\[2\] _02929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08321__A1 _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07461_ _02591_ _02863_ _02866_ _02867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06412_ cpu.uart.divisor\[5\] _01881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_91_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09200_ _04222_ _04203_ _04223_ _04038_ _00463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07392_ _02573_ _02809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09131_ _04170_ _00447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09121__I0 cpu.ROM_addr_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06343_ _01523_ _01791_ _01811_ _01812_ _01813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_17_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09062_ _01025_ _04112_ _04103_ _04117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_72_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06635__A1 _01101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06274_ net63 _01078_ _01208_ _01743_ _01225_ _01744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_72_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_96_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_96_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08013_ _03287_ _03294_ _03295_ _00204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xclkbuf_leaf_25_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_25_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05225_ cpu.regs\[0\]\[2\] _00726_ _00727_ cpu.regs\[3\]\[2\] _00695_ _00696_ _00728_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_114_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05156_ _00663_ _00664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_102_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09964_ _02775_ _04908_ _04915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05087_ _00571_ net98 _00595_ _00597_ _00598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_08915_ cpu.timer_capture\[11\] _03986_ _04001_ _03998_ _04002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09895_ _04853_ _04864_ _04865_ _04866_ _04792_ _00515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05461__I2 cpu.regs\[2\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08846_ _03943_ _03938_ _03944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08560__A1 _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05989_ _01459_ _01461_ _01462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08777_ _02779_ _03883_ _03885_ _03886_ _00377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_67_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07728_ cpu.regs\[6\]\[0\] _03060_ _03061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07659_ _03014_ _03015_ _03016_ _00129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10670_ _00542_ clknet_leaf_59_wb_clk_i cpu.PORTA_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05677__A2 _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09329_ _01126_ _04303_ _04342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_118_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_11_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05864__I _00703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09879__A1 net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08240__I _02809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10104_ _01800_ _05025_ _05023_ _01128_ _05033_ _05034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_10035_ _04769_ _04966_ _04969_ _04958_ _04970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_105_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09004__C _03853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05104__I _00613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06617__A1 _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_113_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05443__I2 cpu.regs\[2\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06961_ _02001_ _02425_ _02426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09680_ _04343_ _04671_ _04681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08700_ _03832_ _03833_ _00353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05912_ _00883_ _00822_ _01386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08631_ _03747_ _03772_ _03784_ _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06892_ _02352_ _02353_ _02355_ _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05843_ _01000_ _01082_ _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05774_ _01044_ _01248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08562_ _02806_ _03714_ _03720_ _03717_ _00328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07513_ _02898_ _02901_ _02905_ _02913_ _02914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08493_ _03654_ _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10101__A1 _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07444_ _02639_ _02351_ _02850_ _02641_ _02851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_36_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05949__I _01421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07375_ _02795_ _02796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_79_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09114_ _00670_ _03130_ _04157_ _04158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10076__B net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06326_ _00961_ _01391_ _01782_ _01384_ _01398_ _01796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_115_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09045_ _04095_ _04101_ _00628_ _00990_ _04102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_72_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06257_ _01715_ _01727_ _01635_ _01728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_32_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05208_ _00685_ _00712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06188_ _01198_ _01659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05139_ cpu.br_rel_dest\[4\] _00648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_8_Left_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09947_ _04902_ _00531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08781__A1 _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09878_ _04843_ _04851_ _00513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08829_ _03929_ _00386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06847__A1 _00689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10653_ _00525_ clknet_leaf_61_wb_clk_i net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_48_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10584_ _00456_ clknet_4_14_0_wb_clk_i cpu.last_addr\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09261__A2 _02315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08772__A1 _02776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05586__A1 _00991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07575__A2 _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10018_ net65 _04954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_47_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05338__A1 cpu.ROM_OEB vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05433__S1 _00910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05490_ _00913_ _00965_ _00966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07160_ _02611_ _02612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07263__A1 _02701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06111_ _01581_ _01582_ _01152_ _01583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09252__A2 _00946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07091_ _00957_ _02541_ _02550_ _02547_ _02551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_41_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06042_ net91 _00873_ _01395_ _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_74_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09801_ _02481_ _04783_ _04758_ _04764_ _04789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07993_ cpu.spi.div_counter\[0\] _03281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09732_ _04690_ _04692_ _04695_ _04731_ _04290_ _04732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_66_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06944_ cpu.PC\[10\] _02409_ _02410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09663_ _04361_ _04649_ _04664_ _04502_ _04665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06875_ _02340_ _01477_ _02292_ _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_82_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09594_ _04372_ _04584_ _04598_ _04471_ _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_05826_ _01299_ _01087_ _01088_ _01300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08614_ cpu.toggle_ctr\[7\] _03763_ _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08545_ _03708_ _03658_ _03709_ _03710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07224__I _01392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05757_ net6 _01229_ _01230_ _01231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_85_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08476_ _03656_ _03660_ _00302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_64_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05688_ _00823_ _01161_ _00007_ _01162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_18_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07427_ _02835_ _00078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_40_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_40_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07358_ _02779_ _02780_ _02782_ _02772_ _00062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_45_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06309_ _01778_ _01779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06057__A2 _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09243__A2 _01869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07289_ _02722_ _02715_ _02716_ _02724_ _02725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_5_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09028_ _01829_ _00649_ _01087_ _04085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_20_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07827__C _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07557__A2 _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06303__I _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output50_I net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05415__S1 _00835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05740__A1 net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10636_ _00508_ clknet_4_14_0_wb_clk_i cpu.ROM_spi_dat_out\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07245__A1 cpu.uart.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10567_ _00439_ clknet_leaf_97_wb_clk_i cpu.base_address\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10498_ _00371_ clknet_leaf_27_wb_clk_i cpu.timer_div_counter\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 io_in[14] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07472__C _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06660_ _02123_ _02125_ _02126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_108_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05611_ _01084_ _01006_ _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_59_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07720__A2 _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06591_ _01291_ _02021_ _02057_ _01474_ _02058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05542_ _01015_ _01016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_86_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08330_ _02813_ _03521_ _03525_ _03547_ _03548_ _00268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_74_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08261_ _03493_ _03488_ _03489_ _03495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_74_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05473_ _00949_ _00950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_22_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07212_ _02534_ _02583_ _02584_ _02539_ _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_61_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08192_ _01321_ _03415_ _03439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_89_Left_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07236__A1 _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06039__A2 _00873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07143_ _02123_ _02596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_112_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08984__A1 cpu.timer_div\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07074_ _02534_ _02535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__05798__A1 _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08603__I cpu.toggle_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06025_ _01104_ net90 _01498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07976_ _00585_ _00662_ _01424_ _03263_ _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XPHY_EDGE_ROW_98_Left_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_87_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09715_ cpu.last_addr\[2\] _04696_ _04715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06927_ _02391_ _02392_ _02393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_97_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09646_ _04646_ _04647_ _04648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_2_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06858_ _02293_ _02323_ _02324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05809_ _00643_ _01282_ _01283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09577_ cpu.regs\[2\]\[1\] _04403_ _04581_ _04582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06789_ _02244_ _02243_ _02255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_08528_ _03696_ _03693_ _03697_ _03695_ _00317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08267__A3 _03436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08459_ _01045_ _03642_ _03647_ _03646_ _00298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_65_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10421_ _00294_ clknet_leaf_33_wb_clk_i cpu.uart.receive_div_counter\[14\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07227__A1 _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10352_ _00225_ clknet_leaf_42_wb_clk_i cpu.uart.dout\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10283_ _00156_ clknet_leaf_3_wb_clk_i cpu.regs\[6\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06968__I _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05713__A1 _01186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_83_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05112__I _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10619_ _00491_ clknet_leaf_67_wb_clk_i cpu.mem_cycle\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07830_ cpu.regs\[2\]\[1\] _03130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_47_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07761_ cpu.regs\[5\]\[5\] _03072_ _03081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09500_ _02830_ _02620_ _04508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06712_ _02175_ _02176_ _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07692_ _03014_ _03032_ _03033_ _00145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06643_ _02108_ _02109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_69_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09431_ _04440_ _04422_ _04441_ _00742_ _04411_ _04442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06574_ _01248_ _02039_ _02040_ _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_09362_ _04272_ _04374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05525_ _00998_ _00999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08313_ cpu.uart.data_buff\[3\] _03531_ _03536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09446__A2 _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09293_ _04295_ _04306_ _04307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08244_ _03477_ _03474_ _03400_ _03482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05456_ cpu.regs\[12\]\[4\] cpu.regs\[13\]\[4\] cpu.regs\[14\]\[4\] cpu.regs\[15\]\[4\]
+ _00932_ _00910_ _00933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_27_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08175_ cpu.spi.counter\[2\] _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_104_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05387_ cpu.regs\[0\]\[1\] cpu.regs\[1\]\[1\] cpu.regs\[2\]\[1\] cpu.regs\[3\]\[1\]
+ _00831_ _00836_ _00867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__08333__I _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06562__B _01196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07126_ _02578_ _02569_ _02579_ _02575_ _00033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_30_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_45_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07057_ _02112_ _02519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08709__A1 _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06008_ _01089_ _01291_ _01481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_7_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06196__A1 cpu.spi.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05692__I _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07959_ _03235_ _03247_ _03248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05625__C _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_qcpu_106 io_oeb[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__08936__C _04015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09629_ _04416_ _04631_ _04632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07412__I _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09437__A2 _04446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_84_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06120__A1 _01591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10404_ _00277_ clknet_leaf_38_wb_clk_i cpu.uart.receive_buff\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08948__A1 _02776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10335_ _00208_ clknet_leaf_66_wb_clk_i cpu.spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08963__A4 _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07620__A1 _02964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10266_ _00139_ clknet_leaf_121_wb_clk_i cpu.regs\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10197_ _00008_ clknet_leaf_85_wb_clk_i net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_17_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_105_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07687__A1 _02981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06290_ cpu.timer_capture\[4\] _01569_ _01252_ _01760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_60_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06111__A1 _01581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05310_ cpu.regs\[0\]\[7\] _00807_ cpu.regs\[2\]\[7\] cpu.regs\[3\]\[7\] _00794_
+ _00795_ _00808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xinput20 io_in[3] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput31 sram_out[5] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05241_ cpu.regs\[2\]\[3\] _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_114_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05172_ _00678_ _00679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_24_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09980_ cpu.PORTB_DDR\[7\] _04918_ _04926_ _04098_ _04927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_58_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08931_ _03947_ _04015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08862_ cpu.timer_capture\[10\] _03902_ _03957_ _03948_ _03958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09364__A1 _04238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05225__I0 cpu.regs\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07813_ _02106_ _03113_ _03114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08793_ _03898_ _03899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07744_ cpu.regs\[6\]\[7\] _03069_ _03070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07675_ cpu.regs\[8\]\[0\] _03023_ _03024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_66_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09414_ _04351_ _04425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06626_ _02091_ _02092_ _02093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07232__I _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06350__B2 _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06350__A1 _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10079__B _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06557_ net47 _01429_ _01434_ _02024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_74_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09345_ _04335_ _04336_ _04337_ _04341_ _04357_ _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_114_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09276_ cpu.Z _02000_ _04264_ _04289_ _04290_ _04291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_47_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06488_ _01622_ _01939_ _01951_ _01955_ _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_05508_ net98 _00638_ _00981_ _00982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_117_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08227_ _03382_ _03462_ _03468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_63_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05439_ _00004_ _00917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__07850__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_1_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08158_ _00676_ _03411_ _03412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08089_ _03350_ _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06405__A2 _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07109_ _02109_ _02565_ _02566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_30_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10120_ cpu.regs\[15\]\[1\] _05045_ _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10051_ _04748_ _04982_ _04983_ _04984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_97_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09130__I1 _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09069__I _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10318_ _00191_ clknet_leaf_44_wb_clk_i cpu.spi.dout\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09346__A1 _03310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10249_ _00122_ clknet_leaf_119_wb_clk_i cpu.regs\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05790_ _01263_ _01264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_37_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06580__A1 _02046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06332__A1 net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07460_ _02135_ _02649_ _02865_ _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06411_ _01877_ _01878_ _01879_ _01880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07391_ cpu.toggle_top\[12\] _02802_ _02808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09130_ cpu.ROM_addr_buff\[5\] _04168_ _04169_ _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06342_ _01524_ _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_84_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09061_ _01591_ _04096_ _04115_ _04109_ _04116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_17_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08012_ cpu.spi.div_counter\[5\] _03293_ _03295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09200__C _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06273_ _01212_ _01739_ _01740_ _01742_ _01743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_72_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05224_ cpu.regs\[2\]\[2\] _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05155_ _00662_ _00663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_69_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06399__A1 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09963_ _04914_ _00535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_77_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05086_ _00596_ cpu.br_rel_dest\[4\] _00597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__06938__A3 cpu.PC\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_65_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_65_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_90_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08914_ _02733_ _03987_ _03988_ _04000_ _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_0_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09894_ cpu.pwm_counter\[0\] _03823_ cpu.pwm_counter\[3\] cpu.pwm_counter\[2\] _04866_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05461__I3 cpu.regs\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08845_ cpu.timer\[8\] _03943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08776_ _02771_ _03886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input12_I io_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05988_ cpu.timer_capture\[9\] _01460_ _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07727_ _03057_ _03060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06287__B _01647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07390__C _02697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07658_ cpu.regs\[10\]\[7\] _03015_ _03016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06609_ _02067_ _02076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07589_ cpu.regs\[12\]\[0\] _02969_ _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_36_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09328_ _04340_ _04341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_80_Left_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09259_ _01488_ _02345_ _02855_ _01600_ _04274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_31_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output80_I net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10103_ _01368_ _05029_ _05032_ _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09879__A2 _03786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10034_ _02497_ _04967_ _04968_ _04969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08551__A2 _03712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09264__B1 _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07600__I _01826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05120__I _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05443__I3 cpu.regs\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06960_ _02124_ _01336_ _01386_ _02425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input4_I io_in[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06891_ _02351_ _02356_ _02357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05911_ _00882_ _00634_ _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08542__A2 _03643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08630_ _03778_ _03747_ _03768_ _03782_ _03783_ _03784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_05842_ cpu.br_rel_dest\[0\] _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_89_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05773_ _01183_ _01185_ _01190_ _01246_ _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_55_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08561_ cpu.toggle_top\[3\] _03715_ _03720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07512_ cpu.uart.receive_div_counter\[0\] _02906_ _02908_ _02912_ _02913_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_08492_ _03670_ _03671_ _00307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06305__A1 _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_112_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_112_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07443_ _02348_ _02350_ _02850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08058__A1 _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09113_ _02838_ _04153_ _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07374_ _01012_ _02674_ _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_79_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06325_ _01701_ _01793_ _01794_ _01795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__07805__A1 _01921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09044_ _04099_ _04085_ _04100_ _04101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_45_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06256_ _01726_ _01717_ _01727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05207_ _00683_ _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06187_ cpu.uart.divisor\[3\] _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_96_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05138_ _00646_ _00647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05069_ cpu.startup_cycle\[6\] cpu.startup_cycle\[5\] cpu.startup_cycle\[4\] _00580_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_96_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09946_ net57 _04894_ _04901_ _04891_ _04902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09877_ cpu.ROM_spi_cycle\[4\] _04849_ _04851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_99_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08828_ cpu.timer_capture\[5\] _03902_ _03928_ _03924_ _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08759_ cpu.timer_div_counter\[7\] _03873_ _03874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_95_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05205__I cpu.regs\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_109_Left_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08049__A1 _02776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10652_ _00524_ clknet_leaf_66_wb_clk_i net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_75_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08516__I _03662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10583_ _00455_ clknet_leaf_77_wb_clk_i cpu.ROM_addr_buff\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_63_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_88_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09261__A3 _02297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09549__A1 _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_118_Left_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05586__A2 _00642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06783__A1 _00807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10017_ _03432_ _04953_ _00550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_97_Right_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08200__B _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05338__A2 cpu.ROM_spi_mode vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06110_ _00952_ _01302_ _01582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09252__A3 _00976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07090_ _02542_ _02549_ _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06041_ _01513_ _01390_ _01335_ _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_23_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09800_ _04786_ _04784_ _04788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07992_ _03279_ _03280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09731_ _04722_ _04725_ _04726_ _04730_ _04731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_5_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06943_ cpu.PC\[9\] _02408_ _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07505__I cpu.uart.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09662_ _04372_ _04653_ _04663_ _04340_ _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06874_ _00710_ _02340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_05825_ _01061_ _01299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08613_ _03760_ cpu.toggle_top\[2\] _03767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09593_ _04594_ _04597_ _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05756_ _01069_ _01013_ _01042_ _01230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_89_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08544_ _03662_ _03709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_85_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06565__B _01198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08475_ cpu.IO_addr_buff\[5\] _03659_ _03592_ _03660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05687_ cpu.regs\[4\]\[7\] cpu.regs\[5\]\[7\] cpu.regs\[6\]\[7\] cpu.regs\[7\]\[7\]
+ _00917_ _00890_ _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_92_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07426_ _02825_ _02834_ _02835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07357_ cpu.timer_top\[4\] _02781_ _02782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06308_ _01103_ _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_32_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_80_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_80_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_72_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07288_ _02723_ _02718_ _02724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09027_ _04083_ _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05695__I _01075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06239_ _01384_ _01689_ _01706_ _01709_ _01710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_32_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08203__A1 _03391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09929_ _02768_ _04888_ _04890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output43_I net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07190__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05740__A2 _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10077__A1 _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07478__C1 _02679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10635_ _00507_ clknet_leaf_71_wb_clk_i cpu.ROM_spi_dat_out\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10566_ _00438_ clknet_leaf_97_wb_clk_i cpu.base_address\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08993__A2 _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10497_ _00370_ clknet_leaf_27_wb_clk_i cpu.timer_div_counter\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09942__A1 _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10001__A1 cpu.PORTA_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput7 io_in[15] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06508__A1 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09170__A2 _00627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07325__I _02705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05610_ _01083_ _01084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_87_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06590_ _02052_ _02054_ _02056_ _02057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05541_ _00601_ _01014_ _01015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_86_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08260_ _03493_ _03494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_52_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05472_ _00948_ _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08191_ _03437_ _03438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07211_ _02660_ _00037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_70_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07142_ _02344_ _02594_ _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_42_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07073_ _00626_ _02534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_30_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_35_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06024_ _01381_ _01496_ _01497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_112_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09933__A1 net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07975_ _00643_ _01146_ _01281_ _03263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_09714_ _04710_ _04712_ _04713_ _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_87_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06926_ _02386_ _02387_ _02390_ _02392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__07235__I _01427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06857_ _02267_ _02322_ _02323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09645_ _02411_ _04446_ _04647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05808_ _01145_ _01281_ _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_2_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09576_ _04404_ _04580_ _04581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06788_ _02171_ _02253_ _02254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05739_ _01024_ _01213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_77_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08527_ cpu.orig_PC\[8\] _03668_ _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08458_ cpu.orig_IO_addr_buff\[1\] _03643_ _03647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_108_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_74_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07409_ _02576_ _02817_ _02577_ _02819_ _00076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_10420_ _00293_ clknet_leaf_33_wb_clk_i cpu.uart.receive_div_counter\[13\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_98_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08389_ _03445_ _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_18_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10351_ _00224_ clknet_leaf_47_wb_clk_i cpu.spi.data_in_buff\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05789__A2 _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10282_ _00155_ clknet_leaf_4_wb_clk_i cpu.regs\[6\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05374__B _00853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09152__A2 cpu.regs\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07163__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06910__A1 _00772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05477__A1 _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10618_ _00490_ clknet_leaf_67_wb_clk_i cpu.mem_cycle\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10549_ _00012_ clknet_leaf_40_wb_clk_i cpu.uart.clr_hb vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09915__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_119_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07760_ _03049_ _03074_ _03080_ _00166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05952__A2 _01424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06711_ _02175_ _02176_ _02177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09430_ _04407_ _04328_ _04441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07691_ cpu.regs\[8\]\[7\] _03032_ _03033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07154__A1 _02135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06642_ cpu.rom_data_dist _02108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_69_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06573_ cpu.timer_div\[7\] _01184_ _02040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09361_ _04372_ _04373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05524_ _00569_ _00993_ _00994_ _00997_ _00998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_82_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08312_ cpu.uart.data_buff\[4\] _03535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_19_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_19_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_35_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09292_ _02828_ _04305_ _04306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08243_ _03400_ _03453_ _03480_ _03470_ _03481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05455_ _00827_ _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_08174_ _03421_ _03422_ _03424_ _00235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05386_ _00826_ _00865_ _00866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07125_ _01646_ _02567_ _02579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07056_ _02473_ _02511_ _02514_ _02517_ _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_88_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09906__A1 _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06007_ _01473_ _01478_ _01479_ _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09445__I _04361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08590__B1 cpu.toggle_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07958_ _03238_ _03246_ _03247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07889_ cpu.spi.dout\[7\] _03174_ _03175_ cpu.spi.data_in_buff\[7\] _03179_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06909_ _02193_ _02205_ _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xwrapped_qcpu_107 io_oeb[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__08893__A1 cpu.timer_capture\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09628_ _03703_ _00880_ _04630_ _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09559_ _04383_ _04555_ _04565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06309__I _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08524__I _03645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10403_ _00276_ clknet_leaf_38_wb_clk_i cpu.uart.receive_buff\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10334_ _00207_ clknet_leaf_63_wb_clk_i net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06959__A1 _00773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10265_ _00138_ clknet_leaf_119_wb_clk_i cpu.regs\[8\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10196_ _00073_ clknet_leaf_12_wb_clk_i cpu.toggle_top\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07384__A1 _02800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05242__S0 _00733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09023__C _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08636__A1 _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput10 io_in[18] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 io_in[6] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_83_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05240_ _00741_ _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput32 sram_out[6] net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_109_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05171_ _00677_ _00678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_116_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09061__A1 _01591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08930_ _04004_ _02750_ _04005_ _04013_ _04014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_0_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08861_ _03259_ _03956_ _03904_ _03957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07812_ _02108_ _03112_ _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_4_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05225__I1 _00726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08792_ _01414_ _01262_ _03897_ _03898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__05925__A2 _01396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07743_ _03058_ _03069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08875__A1 cpu.timer_capture\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07674_ _03020_ _03023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09413_ _04378_ _04422_ _04423_ _04424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06625_ _01963_ _02078_ _02076_ _02092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05233__S0 _00733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06556_ _02022_ _01082_ _01649_ net38 _01432_ _02023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_75_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09344_ _04348_ _04356_ _04357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_35_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09275_ _00678_ _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06487_ _01952_ _01954_ _01812_ _01955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05507_ _00594_ _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08226_ _03382_ _03462_ _03467_ _03450_ _00245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_90_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05438_ _00912_ _00915_ _00916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08157_ cpu.uart.counter\[3\] _03410_ _03411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07108_ _02564_ _02565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__09052__A1 _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05369_ cpu.regs\[0\]\[0\] _00688_ cpu.regs\[2\]\[0\] cpu.regs\[3\]\[0\] _00832_
+ _00837_ _00849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_31_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08088_ _02916_ _03349_ _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07039_ _02492_ _02486_ _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_101_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10050_ _04960_ _02563_ _00574_ _04983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07366__A1 cpu.timer_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06169__A2 _01639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09903__I _04871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07669__A2 _03019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09291__A1 _01104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05852__A1 _01119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10317_ _00190_ clknet_leaf_44_wb_clk_i cpu.spi.dout\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10248_ _00121_ clknet_leaf_110_wb_clk_i cpu.regs\[11\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07357__A1 cpu.timer_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05118__I _00583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10179_ _00056_ clknet_leaf_30_wb_clk_i cpu.timer_capture\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05907__A2 _01380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05463__S0 _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06580__A2 _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06410_ net11 _01073_ _01555_ _01879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06332__A2 _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07390_ _02806_ _02801_ _02807_ _02697_ _00069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_57_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06341_ _01808_ _01810_ _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06272_ cpu.PORTB_DDR\[4\] _01039_ _01741_ _01742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09060_ _02684_ _04105_ _04114_ _04115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08011_ cpu.spi.div_counter\[5\] _03293_ _03294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_72_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05843__A1 _01000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05223_ _00725_ _00726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_69_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05154_ net25 _00662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_12_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09962_ cpu.PORTB_DDR\[2\] _04907_ _04913_ _04904_ _04914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_77_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05085_ cpu.br_rel_dest\[5\] _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08913_ _03960_ _03989_ _04000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07348__A1 _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09893_ cpu.pwm_counter\[5\] cpu.pwm_counter\[4\] cpu.pwm_counter\[7\] _03836_ _04865_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_08844_ _03942_ _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05987_ _01255_ _01460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08775_ cpu.timer_top\[12\] _03884_ _03885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_34_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_34_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07726_ _03058_ _03059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07520__A1 _00676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07657_ _03003_ _03015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06608_ _01943_ _02072_ _02074_ _02075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07588_ _02967_ _02969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09273__A1 cpu.Z vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09327_ _04339_ _04334_ _04340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06539_ _01155_ _01157_ _01160_ _01162_ _02007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_62_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09258_ _00632_ _01052_ _04273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_51_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08209_ cpu.uart.div_counter\[2\] cpu.uart.div_counter\[1\] cpu.uart.div_counter\[0\]
+ _03454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09189_ _03420_ _04215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05647__B _01097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output73_I net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10102_ _01130_ _05026_ _05031_ _01637_ _05032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07339__A1 _02760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10033_ cpu.ROM_addr_buff\[1\] _02494_ _02523_ cpu.ROM_addr_buff\[5\] cpu.ROM_addr_buff\[13\]
+ _04961_ _04968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_105_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06314__A2 _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09264__A1 _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09567__A2 _04315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07578__A1 _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09319__A2 _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05910_ _01383_ _01384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06890_ _02354_ _02355_ _02356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05841_ _01310_ _01312_ _01314_ _01315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05436__S0 _00828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05772_ _01237_ _01240_ _01245_ _01246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08560_ _02804_ _03714_ _03719_ _03717_ _00327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07511_ _02892_ cpu.uart.receive_div_counter\[8\] cpu.uart.receive_div_counter\[0\]
+ _02906_ _02911_ _02912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_89_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08491_ _00672_ _03659_ _03663_ _03671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06305__A2 _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07442_ _02846_ _02848_ _02849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07373_ _02793_ _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_76_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09112_ _04156_ _00442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09255__A1 _01359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06324_ _01701_ _01793_ _01342_ _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_79_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09007__A1 _04039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09043_ _00644_ _01282_ _04100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06255_ _01617_ _01633_ _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_111_Right_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_103_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06186_ _01654_ _01655_ _01656_ _01657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09558__A2 _04562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05206_ _00709_ _00710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05137_ _00645_ _00646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07238__I _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06241__A1 _00722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05068_ cpu.ROM_spi_cycle\[4\] cpu.ROM_spi_cycle\[0\] _00579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_96_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09945_ _02787_ _04895_ _04901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09876_ _04848_ _04850_ _00512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08827_ _03259_ _03927_ _03904_ _03928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08758_ cpu.timer_div_counter\[6\] _03870_ _03873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08689_ _03822_ _03823_ cpu.pwm_counter\[2\] _03825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07709_ _01734_ _03047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10651_ _00523_ clknet_leaf_66_wb_clk_i net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10582_ _00454_ clknet_leaf_77_wb_clk_i cpu.ROM_addr_buff\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05221__I cpu.regs\[1\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09261__A4 _02433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08532__I cpu.PC\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06783__A2 _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10016_ _04793_ _04949_ _04952_ cpu.ROM_OEB _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_116_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_47_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06299__A1 _01738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07611__I _02097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09237__A1 _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09252__A4 _02021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07799__A1 _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_25_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06040_ _01495_ _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07991_ _03261_ _03265_ _03278_ _03167_ _03279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06223__A1 _01112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09730_ _02521_ _04703_ _04727_ _04729_ _04730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__07971__A1 _02793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06774__A2 _00948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06942_ _02399_ _02407_ _02408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05409__S0 _00830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09661_ _04659_ _04662_ _04663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06873_ _02337_ _02338_ _02339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07723__A1 _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05824_ _01294_ _01295_ _01297_ _01298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08612_ cpu.toggle_ctr\[7\] _03763_ _03764_ _03765_ _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_09592_ _00884_ _04465_ _04596_ _04354_ _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05755_ _01228_ _01229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_82_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08543_ cpu.PC\[13\] _03708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_89_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10086__A2 _04087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08474_ _03658_ _03659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05686_ _00840_ _01159_ _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_64_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05501__A3 _00976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07425_ _01406_ _02614_ _02827_ _02833_ _02834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07356_ _02764_ _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07287_ cpu.timer\[1\] _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06307_ _01479_ _01775_ _01776_ _01589_ _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_45_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09026_ _04082_ _04083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06462__A1 _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06238_ _01707_ _01688_ _01708_ _00981_ _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_5_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06169_ _00982_ _01639_ _01640_ _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_111_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09928_ _02760_ _04887_ _04889_ _00525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09859_ _04835_ _04812_ _04805_ _04811_ _04838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_99_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09467__A1 _02605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output36_I net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10634_ _00506_ clknet_leaf_71_wb_clk_i cpu.ROM_spi_dat_out\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10565_ _00437_ clknet_leaf_19_wb_clk_i cpu.IO_addr_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10496_ _00369_ clknet_leaf_27_wb_clk_i cpu.timer_div_counter\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06205__A1 cpu.timer_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09093__I _04141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput8 io_in[16] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06508__A2 _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_108_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05540_ _00567_ _00568_ _01014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07341__I _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05471_ _00912_ _00915_ _00920_ _00922_ _00948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_08190_ _03407_ _03436_ _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07210_ _02648_ _02659_ _02660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_116_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07141_ _02358_ _02357_ _02594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05796__I _01009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07072_ _02471_ _02518_ _02530_ _02533_ _00025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_2_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06023_ _00717_ _01495_ _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_2_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07974_ _01320_ _01174_ _03262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09713_ cpu.last_addr\[2\] cpu.ROM_addr_buff\[2\] _04696_ _04713_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_87_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06925_ _02386_ _02387_ _02390_ _02391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06856_ _02321_ _00944_ _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09644_ cpu.PC\[12\] _04646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_97_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05807_ _00645_ _00648_ _01281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_2_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09575_ _04579_ _04580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06787_ _00709_ _00974_ _02253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05738_ _01211_ _01212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_65_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08526_ _02399_ _03696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_92_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08457_ _01046_ _03642_ _03644_ _03646_ _00297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05669_ _01142_ _01143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07408_ _02532_ _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_21_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08388_ _03588_ _03581_ _03590_ _03583_ _03591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_98_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07339_ _02760_ _02765_ _02767_ _02683_ _00058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09621__A1 _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10350_ _00223_ clknet_leaf_47_wb_clk_i cpu.spi.data_in_buff\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09009_ _03849_ _04066_ _04071_ _04070_ _00424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_10281_ _00154_ clknet_leaf_2_wb_clk_i cpu.regs\[6\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10117__I _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08188__A1 _03432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09688__A1 _04413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05410__A2 _00825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06910__A2 _02009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09160__I0 cpu.ROM_addr_buff\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05477__A2 _00952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10617_ _00489_ clknet_leaf_85_wb_clk_i cpu.mem_cycle\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10548_ _00421_ clknet_leaf_84_wb_clk_i cpu.rom_data_dist vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10479_ _00352_ clknet_leaf_102_wb_clk_i cpu.pwm_counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_71_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09679__A1 cpu.PC\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06710_ _02147_ _02148_ _02176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09551__I _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07690_ _03021_ _03032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_69_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06641_ _02106_ _02107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06572_ cpu.spi.dout\[7\] _01566_ _01421_ _02038_ _02039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__07071__I _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09360_ _04335_ _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05523_ _00995_ _00996_ _00997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08311_ _02800_ _03522_ _03526_ _03533_ _03534_ _00263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_75_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09291_ _01104_ _04304_ _04305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08242_ _03400_ _03477_ _03474_ _03480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_05454_ _00592_ _00931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_59_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_59_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_62_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08173_ _03162_ _03423_ _03417_ _03424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05385_ cpu.regs\[4\]\[1\] cpu.regs\[5\]\[1\] cpu.regs\[6\]\[1\] cpu.regs\[7\]\[1\]
+ _00831_ _00836_ _00865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_07124_ _02557_ _02578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07055_ _02515_ _02516_ _02517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_88_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06006_ _01300_ _01479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07957_ _03240_ _03245_ _03242_ _03246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06908_ _02199_ _02203_ _02374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07888_ _03178_ _00196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_69_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09461__I _04340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06353__B1 _01822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06839_ _02302_ _02304_ _02305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09627_ _04628_ _04609_ _04629_ _04630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xwrapped_qcpu_108 io_out[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09558_ _04560_ _04562_ _04563_ _04564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08509_ _03682_ _03683_ _00312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09489_ _04236_ _04498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_12_Left_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10402_ _00275_ clknet_leaf_38_wb_clk_i cpu.uart.receive_buff\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06408__A1 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10333_ _00206_ clknet_leaf_46_wb_clk_i cpu.spi.div_counter\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06959__A2 _02128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10264_ _00137_ clknet_leaf_108_wb_clk_i cpu.regs\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10195_ _00072_ clknet_leaf_12_wb_clk_i cpu.toggle_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05919__C2 _01392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08696__B _03709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_21_Left_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_105_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05147__A1 _00616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05242__S1 _00734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09133__I0 cpu.ROM_addr_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08636__A2 _03786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput11 io_in[19] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput22 io_in[7] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput33 sram_out[7] net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05170_ _00676_ _00677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08860_ _03207_ _03955_ _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07811_ _02116_ _02582_ _02561_ _03112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__08572__A1 _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05225__I2 _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_106_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_106_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08791_ _00623_ _01148_ _03263_ _03897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_79_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07742_ _03053_ _03060_ _03068_ _00160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07673_ _03021_ _03022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10131__A1 _01921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09412_ _04354_ _04423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06624_ _01963_ _02076_ _02078_ _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__05233__S1 _00734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09343_ _00989_ _04350_ _04353_ _04355_ _04356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06555_ net58 _02022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05506_ _00980_ net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09274_ _02000_ _04288_ _04289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06486_ _01937_ _01953_ _01954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08225_ cpu.uart.div_counter\[5\] _03453_ _03466_ _03448_ _03467_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05437_ _00913_ _00914_ _00846_ _00915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_99_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08156_ cpu.uart.counter\[0\] cpu.uart.counter\[1\] cpu.uart.counter\[2\] _03410_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_7_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05368_ _00843_ _00844_ _00847_ _00848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_31_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07107_ _02561_ _02563_ _02564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07063__A1 cpu.ROM_addr_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08087_ cpu.uart.receiving _03348_ _03349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06405__A4 _01084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05299_ cpu.regs\[1\]\[6\] _00798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07038_ _02499_ _02500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_3_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05216__I2 cpu.regs\[10\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08989_ _02706_ _04034_ _04056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10122__A1 cpu.regs\[15\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09115__I0 cpu.ROM_addr_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05224__I cpu.regs\[2\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_4_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_4_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10316_ _00189_ clknet_leaf_104_wb_clk_i cpu.regs\[2\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10247_ _00120_ clknet_leaf_118_wb_clk_i cpu.regs\[11\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10178_ _00055_ clknet_leaf_23_wb_clk_i cpu.timer_capture\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05463__S1 _00935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05134__I _00642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06340_ net94 _01809_ _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06271_ _01210_ _01741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08010_ _03287_ _03292_ _03293_ _00203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__05843__A2 _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05222_ _00724_ _00725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_114_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05153_ _00629_ _00660_ _00661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09961_ _02685_ _04908_ _04913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_77_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05084_ _00589_ _00593_ _00594_ _00595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__09209__C _03421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08912_ _03999_ _00399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08545__A1 _03708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09892_ _04856_ _04858_ _04863_ _04864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08843_ cpu.timer_capture\[7\] _03930_ _03941_ _03924_ _03942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05986_ _01086_ _01459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08774_ _03875_ _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10104__A1 _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07725_ _03057_ _03058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07656_ _02097_ _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_74_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_74_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07587_ _02967_ _02968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06607_ _01834_ _02073_ _02074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09326_ _04338_ _00651_ _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06538_ _02004_ _02005_ _01297_ _02006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09257_ _04236_ _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_106_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08208_ _03440_ _03453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06469_ _01936_ _01937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_106_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09188_ _04212_ _04203_ _04214_ _04038_ _00460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05685__I2 cpu.regs\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08139_ _02891_ _03375_ _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08784__A1 _00613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10101_ _01525_ _05030_ _05031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05647__C _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output66_I net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09914__I _04871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10032_ cpu.ROM_addr_buff\[9\] _02524_ _04967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_4_4_0_wb_clk_i clknet_0_wb_clk_i clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07511__A2 cpu.uart.receive_div_counter\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09264__A2 _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_15_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_113_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09096__I _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08775__A1 cpu.timer_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09045__B _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05840_ _01313_ _01314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05436__S1 _00910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07344__I _02771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07510_ _02909_ _02910_ _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05771_ _01241_ _01244_ _01188_ _01245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08490_ cpu.orig_flags\[2\] _03655_ _03670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_54_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07441_ _02847_ _02848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05364__I1 cpu.regs\[9\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07372_ _00678_ _02793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09111_ cpu.ROM_addr_buff\[0\] _04154_ _04155_ _04156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_57_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09255__A2 _01779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06323_ _01347_ _01788_ _01792_ _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_79_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09042_ _00646_ _01103_ _00571_ _04099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_06254_ _01723_ _01724_ _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06185_ net9 _01073_ _01197_ _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05205_ cpu.regs\[1\]\[1\] _00709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08766__A1 _02671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05136_ _00596_ _00645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_121_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_121_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05067_ _00577_ _00578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09944_ _04900_ _00530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06241__A2 _00730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09875_ _03551_ _04849_ _04850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08826_ cpu.timer\[5\] _03926_ _03927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07254__I _02694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_93_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07741__A2 _03058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05969_ cpu.uart.divisor\[9\] _01442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08757_ _03861_ _03872_ _00371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08794__B _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08688_ _03822_ _03823_ _03824_ _00350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07708_ _03045_ _03039_ _03046_ _00148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_95_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07639_ _03003_ _03004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10650_ _00522_ clknet_leaf_67_wb_clk_i net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_118_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07257__A1 _02695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09309_ _02831_ _04292_ _04322_ _04323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10581_ _00453_ clknet_leaf_77_wb_clk_i cpu.ROM_addr_buff\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07429__I cpu.PC\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10015_ _04760_ _04950_ _04951_ _04952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_47_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_4_Left_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07990_ _03277_ _03278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07971__A2 _03259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06941_ cpu.PC\[7\] _02400_ _02406_ _02407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_5_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09173__A1 cpu.ROM_addr_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05982__A1 cpu.timer_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09660_ _00931_ _04465_ _04661_ _04354_ _04662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05409__S1 _00835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07074__I _02534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08611_ cpu.toggle_ctr\[6\] _03765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06872_ _00741_ _00856_ _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05823_ _01296_ _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09591_ _04093_ _04579_ _04595_ _04467_ _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05754_ _01069_ _01071_ _01228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08542_ cpu.orig_PC\[13\] _03643_ _03707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07487__A1 cpu.uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08473_ _03657_ _03658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09476__A2 _00647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_59_Left_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05685_ cpu.regs\[0\]\[7\] cpu.regs\[1\]\[7\] cpu.regs\[2\]\[7\] cpu.regs\[3\]\[7\]
+ _00917_ _00890_ _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07424_ _02831_ _02591_ _02611_ _02832_ _02833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_92_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05322__I cpu.PORTB_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07355_ _02764_ _02780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08987__A1 cpu.timer_div\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07286_ _01585_ _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06306_ _00952_ _01584_ _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09025_ _01288_ _04082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06237_ _00925_ _01390_ _01708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07249__I _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06153__I _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06168_ net28 _01334_ _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05119_ _00626_ _00627_ _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_06099_ cpu.timer_capture\[2\] _01420_ _01252_ _01570_ _01571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_68_Left_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09927_ net79 _04888_ _02682_ _04889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09858_ _04835_ _04821_ _04823_ _04837_ _04792_ _00507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08911__A1 cpu.timer_capture\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07714__A2 _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09789_ _04778_ _04761_ _04779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05725__A1 cpu.uart.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08809_ cpu.timer_capture\[2\] _03899_ _03912_ _03913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08808__I _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05740__A4 _01084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_77_Left_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07712__I _01825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10077__A3 _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10633_ _00505_ clknet_leaf_70_wb_clk_i cpu.ROM_spi_dat_out\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08978__A1 _04047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08543__I cpu.PC\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10564_ _00436_ clknet_leaf_19_wb_clk_i cpu.IO_addr_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10495_ _00368_ clknet_leaf_27_wb_clk_i cpu.timer_div_counter\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05388__B _00853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07159__I _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07402__A1 _02053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08699__B _03709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08902__A1 cpu.timer_capture\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput9 io_in[17] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05851__B _01075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08130__A2 cpu.uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05470_ _00931_ _00946_ _00947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_116_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08969__A1 cpu.timer_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07140_ _02592_ _02593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_82_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07069__I _00619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07071_ _02532_ _02533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_2_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06022_ _01493_ _01494_ _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_100_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09394__A1 _02855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07973_ _00663_ _03166_ _03261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09712_ _04196_ _04711_ _04712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06924_ _02194_ _02388_ _02389_ _02390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_87_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05707__A1 _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09643_ _03703_ _04554_ _04641_ _04645_ _00484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06855_ _00689_ _02321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_96_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05806_ _01110_ _01118_ _00646_ _01280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_09574_ _03135_ _04577_ _04578_ _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08525_ _02654_ _03693_ _03694_ _03695_ _00316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06786_ _02251_ _02248_ _02252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05737_ _00993_ _01210_ _01211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_108_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08456_ _03645_ _03646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05668_ _01141_ _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08387_ _03588_ _03589_ _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_21_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07407_ _02571_ _02817_ _02572_ _02818_ _00075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_107_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05599_ _01072_ _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07338_ cpu.timer_top\[0\] _02766_ _02767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_98_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07269_ _02706_ _02691_ _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07632__A1 cpu.regs\[11\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09008_ _02909_ _04067_ _04071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10280_ _00153_ clknet_leaf_108_wb_clk_i cpu.regs\[7\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09924__A3 _03897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06199__A1 cpu.timer_div\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09137__A1 _02654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_85_Left_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07871__A1 _00620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10616_ _00488_ clknet_leaf_68_wb_clk_i cpu.mem_cycle\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08273__I _03503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_94_Left_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10547_ _00420_ clknet_leaf_31_wb_clk_i cpu.timer_div\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07623__A1 _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10478_ _00351_ clknet_leaf_101_wb_clk_i cpu.pwm_counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08222__B _03464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06640_ _00618_ _00583_ _02106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_69_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06362__A1 _01830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06571_ _02035_ _02036_ _02037_ _02038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05522_ cpu.IO_addr_buff\[2\] _00996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08310_ cpu.uart.data_buff\[2\] _03531_ _03534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09290_ _00905_ _04303_ _04304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08241_ _03477_ _03476_ _03478_ _03479_ _00248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05453_ _00930_ net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07862__A1 _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08172_ cpu.spi.counter\[0\] cpu.spi.counter\[1\] _03423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_103_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05384_ _00843_ _00863_ _00847_ _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_27_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07123_ _02576_ _02569_ _02577_ _02575_ _00032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_6_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07054_ cpu.spi_clkdiv _02472_ _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07090__A2 _02549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_99_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_99_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_28_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_28_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06005_ _01474_ _01285_ _01477_ _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09367__A1 cpu.PC\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_7_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05928__A1 _01337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07971__B cpu.needs_timer_interrupt vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07956_ _01463_ cpu.timer\[1\] _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input28_I sram_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06907_ _02208_ _02210_ _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_106_Right_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07887_ cpu.spi.dout\[6\] _03174_ _03175_ cpu.spi.data_in_buff\[6\] _03178_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_97_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07262__I _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06353__A1 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06838_ _02303_ _02299_ _02304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09626_ _03700_ _01127_ _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xwrapped_qcpu_109 io_out[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09557_ _04560_ _04562_ _04458_ _04563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06769_ _02232_ _02234_ _02235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08508_ _02861_ _03674_ _03677_ _03683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09488_ _04493_ _04496_ _04497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06105__A1 cpu.toggle_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08439_ _03570_ _03629_ _03632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_108_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_102_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06656__A2 _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05510__I net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10401_ _00274_ clknet_leaf_43_wb_clk_i cpu.uart.receive_buff\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06408__A2 _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10332_ _00205_ clknet_leaf_46_wb_clk_i cpu.spi.div_counter\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output96_I net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10263_ _00136_ clknet_leaf_110_wb_clk_i cpu.regs\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10194_ _00071_ clknet_leaf_13_wb_clk_i cpu.toggle_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06592__A1 _01392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06497__B _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06344__B2 _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06344__A1 _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput12 io_in[1] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_71_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05420__I _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput23 io_in[8] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05622__A3 _01051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08790_ _03895_ _03896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_4_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05225__I3 cpu.regs\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07810_ _02462_ _03110_ _03111_ _00185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07741_ cpu.regs\[6\]\[6\] _03058_ _03068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07672_ _03020_ _03021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09411_ _02860_ _04414_ _04422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06623_ _01625_ _02080_ _02089_ _02090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09342_ _04354_ _04355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06554_ _01929_ _02021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_114_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05505_ _00978_ _00979_ _00980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_47_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09273_ cpu.Z _04083_ _04263_ _04287_ _04288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06485_ net95 _01808_ _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08224_ cpu.uart.div_counter\[5\] _03461_ _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05330__I cpu.PORTB_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05436_ cpu.regs\[8\]\[3\] cpu.regs\[9\]\[3\] cpu.regs\[10\]\[3\] cpu.regs\[11\]\[3\]
+ _00828_ _00910_ _00914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_28_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08155_ _03408_ _03409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05367_ _00846_ _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09737__I _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07106_ _02562_ _02114_ _02496_ _02563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_70_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08086_ cpu.uart.receive_counter\[0\] cpu.uart.receive_counter\[1\] cpu.uart.receive_counter\[3\]
+ cpu.uart.receive_counter\[2\] _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_101_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05298_ _00787_ _00796_ _00797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07037_ _02494_ _02495_ _02498_ _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_30_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08988_ _04055_ _00419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07939_ cpu.timer\[5\] _03228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06326__A1 _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09609_ _03146_ _04427_ _04613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09115__I1 _04158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09276__B1 _04264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06629__A2 _02095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05240__I _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10315_ _00188_ clknet_leaf_104_wb_clk_i cpu.regs\[2\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06071__I _01141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10246_ _00119_ clknet_leaf_118_wb_clk_i cpu.regs\[11\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10177_ _00054_ clknet_leaf_23_wb_clk_i cpu.timer_capture\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_44_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06270_ net55 _01172_ _01213_ _01084_ _01740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_56_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05221_ cpu.regs\[1\]\[2\] _00724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05152_ _00658_ _00659_ _00660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09990__A1 cpu.PORTA_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09960_ _04912_ _00534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_69_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05083_ cpu.base_address\[3\] cpu.base_address\[2\] _00594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_90_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08911_ cpu.timer_capture\[10\] _03986_ _03997_ _03998_ _03999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_40_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09742__A1 _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09891_ _04859_ _04860_ _04861_ _04862_ _04863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__06556__B2 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_83_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08842_ _03895_ _03937_ _03940_ _03941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05985_ _01420_ _01455_ _01457_ _01458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08773_ _03875_ _03883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07724_ _02935_ _03036_ _03057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07655_ _02983_ _03005_ _03013_ _00128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05325__I cpu.PORTA_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Left_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06606_ _01848_ _01941_ _02072_ _02073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_87_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07586_ _02937_ _02966_ _02967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09325_ cpu.uart.busy cpu.spi.busy _04338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06537_ _01773_ _01294_ _02005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09256_ _01484_ _01289_ _04271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06468_ _00803_ _01936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_118_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_43_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_43_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08207_ _03379_ _03391_ _03452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09895__C _04792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05419_ _00889_ _00893_ _00895_ _00897_ _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_35_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09187_ cpu.ROM_addr_buff\[4\] _04213_ _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06399_ _01368_ _01851_ _01863_ _01867_ _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_08138_ cpu.uart.div_counter\[10\] _03392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08069_ cpu.spi.data_in_buff\[0\] _03334_ _03336_ cpu.spi.data_in_buff\[1\] _03338_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10040__B2 cpu.ROM_addr_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10040__A1 cpu.ROM_addr_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10100_ _00817_ _01952_ _05030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10031_ _02483_ _04966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07715__I _01920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06547__A1 _01924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output59_I net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08974__C _04015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08527__A2 _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10229_ _00102_ clknet_leaf_114_wb_clk_i cpu.regs\[13\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05770_ _01243_ _01244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_0_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07360__I _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08456__I _03645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07440_ _02837_ _02847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07371_ _02791_ _02780_ _02792_ _02786_ _00065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_45_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10636__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09110_ _04061_ _04155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_44_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06322_ _01347_ _01791_ _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09041_ _03445_ _04098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_79_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06253_ _01632_ _01704_ _01722_ _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_111_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06184_ net24 _01221_ _01229_ _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05748__C _01221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05204_ _00694_ _00704_ _00706_ _00707_ _00708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_25_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05135_ _00643_ _00644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05066_ cpu.ROM_spi_cycle\[3\] cpu.ROM_spi_cycle\[2\] cpu.ROM_spi_cycle\[1\] _00577_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_09943_ net56 _04894_ _04899_ _04891_ _04900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06241__A3 _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09874_ cpu.ROM_spi_cycle\[3\] _04846_ _04849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09191__A2 _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08825_ _03231_ _03858_ _03920_ _03926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA_input10_I io_in[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05968_ _01427_ _01428_ _01438_ _01439_ _01440_ _01441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08756_ _03193_ _03870_ _03872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10089__A1 _01310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08687_ _03822_ _03823_ _03371_ _03824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05899_ _00906_ _00877_ _01373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07707_ cpu.regs\[7\]\[2\] _03043_ _03046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07270__I _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07638_ _03002_ _03003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_82_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07569_ cpu.regs\[13\]\[2\] _02953_ _02956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09308_ _00625_ _04320_ _04321_ _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_36_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10580_ _00452_ clknet_leaf_77_wb_clk_i cpu.ROM_addr_buff\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09239_ _04252_ _04254_ _04251_ _00471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_35_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08969__C _04015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10014_ _02527_ _02485_ _04951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07193__A1 _02135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_63_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06524__I cpu.timer_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10004__A1 _02706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09945__A1 _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_74_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_105_Left_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06940_ cpu.PC\[5\] _02405_ _02406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input2_I io_in[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06871_ _00726_ _00871_ _02337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05822_ _01061_ _01064_ _01087_ _01296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08610_ cpu.toggle_top\[6\] _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__07184__A1 _02015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_84_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09590_ _03135_ _04426_ _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06931__A1 _02135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05753_ net21 _01225_ _01226_ _01227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_89_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08541_ _03705_ _03706_ _00321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08472_ _00624_ _00659_ _03638_ _03657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_49_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05684_ _01155_ _01157_ _01158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07423_ _02593_ _02347_ _02597_ _02630_ _02832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_114_Left_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07354_ _02778_ _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07285_ _02710_ _02721_ _00050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_72_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06305_ _01579_ _01769_ _01774_ _01775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XPHY_EDGE_ROW_93_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09024_ _02624_ _04081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06236_ _01341_ _01517_ _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06167_ _01610_ _01628_ _01636_ net92 _01638_ _01639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_05118_ _00583_ _00627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06098_ _01546_ _01422_ _01568_ _01569_ _01570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_111_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09926_ _04886_ _04888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09857_ cpu.ROM_spi_dat_out\[5\] _04790_ _04836_ _04771_ _04837_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09788_ _02474_ _04778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08808_ _02681_ _03912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_96_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08739_ _03860_ _03861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05513__I _00986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10632_ _00504_ clknet_leaf_71_wb_clk_i cpu.ROM_spi_dat_out\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_52_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10563_ _00435_ clknet_leaf_19_wb_clk_i cpu.IO_addr_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09927__A1 net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10494_ _00367_ clknet_leaf_29_wb_clk_i cpu.timer_div_counter\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06913__A1 _00807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05423__I _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07070_ _02531_ _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06021_ _00866_ _00868_ _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09918__A1 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09711_ cpu.last_addr\[0\] cpu.ROM_addr_buff\[0\] _04711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07085__I _00665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07972_ _03182_ _00616_ _03260_ _00198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06923_ _02197_ _02206_ _02389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_87_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09642_ _04411_ _04642_ _04644_ _04645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06854_ _02319_ _02312_ _02314_ _02320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_117_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05805_ _01059_ _01279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06785_ _00805_ _00855_ _02251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09573_ _02409_ _04479_ _04578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05736_ _00995_ _00604_ _01022_ _01210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_08524_ _03645_ _03695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_89_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05333__I cpu.PORTA_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08455_ _02573_ _03645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05667_ _01109_ _01140_ _01141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08409__B2 _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08386_ _02899_ _03582_ _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05598_ _01069_ _01071_ _01072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_21_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07406_ _02560_ _02817_ _02570_ _02818_ _00074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_07337_ _02764_ _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_116_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07268_ _02705_ _02706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_61_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09909__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09007_ _04039_ _04066_ _04069_ _04070_ _00423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06219_ _01688_ _01689_ _01690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07199_ net20 _02592_ _02649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09909_ net61 _04873_ _04877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07148__A1 _01116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output41_I net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06123__A2 _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07871__A2 _03167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10615_ _00487_ clknet_leaf_67_wb_clk_i cpu.mem_cycle\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09073__A1 _01779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_3_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10546_ _00419_ clknet_leaf_30_wb_clk_i cpu.timer_div\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10477_ _00350_ clknet_leaf_101_wb_clk_i cpu.pwm_counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_118_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09385__I _04340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07387__A1 _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06434__I0 cpu.regs\[8\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05493__S0 _00829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06362__A2 _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06570_ cpu.spi.divisor\[7\] _01243_ _01187_ _02037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_87_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05521_ cpu.IO_addr_buff\[3\] _00995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08240_ _02809_ _03479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05452_ _00908_ _00926_ _00929_ _00930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08171_ cpu.spi.counter\[1\] _03418_ _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07122_ _01591_ _02567_ _02577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05383_ cpu.regs\[8\]\[1\] cpu.regs\[9\]\[1\] cpu.regs\[10\]\[1\] cpu.regs\[11\]\[1\]
+ _00830_ _00835_ _00863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_42_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07053_ cpu.ROM_spi_cycle\[0\] _02515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_70_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05625__A1 _00989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06004_ _01475_ _01476_ _01477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_100_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07378__A1 _00979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05328__I cpu.PORTB_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_68_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_68_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07955_ _03226_ _03229_ _03241_ _03243_ _03244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06906_ _02238_ _02370_ _02371_ _02372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07886_ _03177_ _00195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_97_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05236__S0 _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07543__I _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09625_ _03701_ _01127_ _04628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06837_ _00771_ _00856_ _02303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09556_ _04529_ _01110_ _04561_ _04562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_06768_ _02233_ _02234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05719_ _01039_ _01013_ _01016_ _01193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08507_ cpu.orig_PC\[3\] _03672_ _03682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07302__A1 _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09487_ _01829_ _04350_ _04495_ _04423_ _04496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06105__A2 _01416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06699_ _02160_ _02164_ _02165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08438_ _03566_ _03630_ _03575_ _03631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_34_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08369_ _03574_ _03575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10400_ _00273_ clknet_leaf_43_wb_clk_i cpu.uart.receive_buff\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10331_ _00204_ clknet_leaf_46_wb_clk_i cpu.spi.div_counter\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05616__A1 _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10262_ _00135_ clknet_leaf_115_wb_clk_i cpu.regs\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07718__I _02015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10193_ _00070_ clknet_leaf_14_wb_clk_i cpu.toggle_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05238__I cpu.regs\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08869__A1 _03909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_34_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06069__I _01541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05855__A1 _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput13 io_in[20] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput24 io_in[9] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10529_ _00402_ clknet_leaf_25_wb_clk_i cpu.timer_capture\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_12_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_73_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06583__A2 _01049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07740_ _03051_ _03060_ _03067_ _00159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07671_ _01140_ _02965_ _03020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_59_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09410_ _04416_ _04420_ _04421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06622_ _01523_ _02063_ _02082_ _01367_ _02088_ _02089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_87_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09341_ _01331_ _01133_ _00957_ _04354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06553_ _01144_ _01314_ _01098_ _02020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09285__A1 cpu.PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08194__I _03440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05504_ _00859_ _00979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_118_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09272_ _04083_ _04286_ _04287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06484_ _00786_ _00804_ _01808_ _01952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xclkbuf_leaf_115_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_115_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_16_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08223_ _03463_ _03465_ _00244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05435_ _00840_ _00913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08154_ _03407_ _03408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05366_ _00845_ _00846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08085_ cpu.uart.receive_buff\[0\] _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07105_ cpu.mem_cycle\[5\] _02562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07036_ _02497_ _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09239__B _04251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05297_ cpu.regs\[4\]\[6\] cpu.regs\[5\]\[6\] cpu.regs\[6\]\[6\] cpu.regs\[7\]\[6\]
+ _00794_ _00795_ _00796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06023__A1 _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08987_ cpu.timer_div\[6\] _04046_ _04054_ _04050_ _04055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07273__I _02574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07938_ cpu.timer\[6\] _03227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05209__S0 _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07869_ cpu.spi.counter\[3\] cpu.spi.counter\[2\] cpu.spi.counter\[4\] _03162_ _03166_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_98_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09608_ _04378_ _04610_ _04611_ _04385_ _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_104_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09539_ _04093_ _04533_ _04545_ _04467_ _04546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_38_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09276__A1 cpu.Z vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_118_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09028__A1 _01829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06262__A1 net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07448__I _00726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10314_ _00187_ clknet_leaf_103_wb_clk_i cpu.regs\[2\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10245_ _00118_ clknet_leaf_119_wb_clk_i cpu.regs\[11\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10176_ _00053_ clknet_leaf_22_wb_clk_i cpu.timer_capture\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_66_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09267__A1 _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07817__A2 _01404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09019__A1 _02811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08490__A2 _03655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05220_ cpu.regs\[4\]\[2\] cpu.regs\[5\]\[2\] cpu.regs\[6\]\[2\] cpu.regs\[7\]\[2\]
+ _00711_ _00712_ _00723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_107_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05151_ cpu.instr_cycle\[3\] cpu.instr_cycle\[1\] _00659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_52_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_77_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05687__S0 _00917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05082_ _00590_ cpu.instr_buff\[14\] _00591_ _00592_ _00593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_90_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08910_ _03947_ _03998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09890_ cpu.pwm_top\[3\] cpu.pwm_counter\[3\] _04862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_0_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08841_ _03938_ _03939_ _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06556__A2 _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05984_ cpu.timer_capture\[1\] _01420_ _01456_ _01178_ _01457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_08772_ _02776_ _03876_ _03882_ _03879_ _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_79_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07723_ _03014_ _03055_ _03056_ _00153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08917__I _03985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07654_ cpu.regs\[10\]\[6\] _03003_ _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06605_ _01362_ _02063_ _02071_ _02072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07585_ _02965_ _02966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09324_ _04237_ _04331_ _04337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06536_ _01998_ _01999_ _02003_ _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09255_ _01359_ _01779_ _04268_ _04269_ _04270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__05819__A1 _00984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06467_ _00804_ _01934_ _01935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08206_ cpu.uart.div_counter\[2\] _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05418_ _00825_ _00896_ _00853_ _00897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09186_ _04201_ _04213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06398_ _01865_ _01866_ _01867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_31_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07268__I _02705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08137_ cpu.uart.div_counter\[0\] _03391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05349_ _00828_ _00829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_31_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08068_ _03331_ _03334_ _03336_ _03337_ _00217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_101_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_83_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_83_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06172__I _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07019_ cpu.startup_cycle\[5\] _02481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_101_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_12_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_12_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10030_ _04954_ _04957_ _04965_ _02818_ _00551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__06547__A2 _01926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09497__A1 _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05960__B _01203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06483__A1 _01395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10228_ _00101_ clknet_leaf_121_wb_clk_i cpu.regs\[13\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10159_ _00036_ clknet_leaf_99_wb_clk_i cpu.regs\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07370_ cpu.timer_top\[7\] _02781_ _02792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06321_ _00768_ _01790_ _01791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09040_ _04084_ _04092_ _04096_ _01105_ _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06252_ _01632_ _01722_ _01704_ _01723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05203_ _00003_ _00707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_06183_ _01650_ _01651_ _01653_ _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_4_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05134_ _00642_ _00643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_13_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05065_ _00574_ _00575_ _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09942_ _02783_ _04895_ _04899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09873_ cpu.ROM_spi_cycle\[3\] _04846_ _04848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08824_ _03925_ _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05336__I cpu.PORTA_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08755_ _03863_ _03870_ _03871_ _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05967_ _01198_ _01440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07706_ _01642_ _03045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08686_ cpu.pwm_counter\[1\] _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05898_ _00635_ _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_95_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07637_ _01140_ _02101_ _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07568_ _01543_ _02952_ _02955_ _00099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06519_ cpu.timer_div\[6\] _01185_ _01986_ _01182_ _01987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_76_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09307_ _00624_ cpu.instr_cycle\[1\] _01148_ _04321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07499_ cpu.uart.divisor\[11\] cpu.uart.receive_div_counter\[11\] _02900_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08454__A2 _03643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09238_ cpu.orig_flags\[2\] _04247_ _04249_ _04253_ _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_63_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09169_ cpu.last_addr\[0\] _04199_ _04200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_8_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output71_I net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07726__I _03058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10013_ _00575_ _04733_ _04950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_99_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_74_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06870_ _00726_ _00856_ _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05156__I _00663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05821_ cpu.C _01103_ _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05752_ _01072_ _01226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_82_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08540_ _02414_ _03658_ _03689_ _03706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08467__I _03645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08133__B2 _02679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08471_ cpu.orig_IO_addr_buff\[5\] _03655_ _03656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05683_ _00823_ _01156_ _00845_ _01157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_85_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07422_ _02830_ _02831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_85_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07353_ _00962_ _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09633__A1 _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07284_ cpu.timer_capture\[0\] _02712_ _02720_ _02721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06447__B2 _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06304_ _00925_ _01294_ _01302_ _01773_ _01774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06447__A1 _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09023_ _02815_ _04073_ _04080_ _04078_ _00429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06235_ _01519_ _01705_ _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_79_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06166_ _01637_ _01638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_111_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05117_ _00576_ _00626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06097_ _01248_ _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09925_ _04886_ _04887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09856_ _02504_ _02506_ _04836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08807_ _02729_ _03908_ _03910_ _03911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09787_ _04775_ _04777_ _02710_ _00496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_99_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06999_ _02097_ _02462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08738_ _00678_ _03859_ _03860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08669_ cpu.toggle_ctr\[10\] _03810_ _03813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06686__A1 _00762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10631_ _00503_ clknet_leaf_71_wb_clk_i cpu.ROM_spi_dat_out\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10562_ _00434_ clknet_leaf_54_wb_clk_i cpu.IO_addr_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09001__I _04065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10493_ _00366_ clknet_leaf_28_wb_clk_i cpu.timer_div_counter\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06360__I _00647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09671__I _04671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08236__B _03440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09846__I _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06020_ _00862_ _00864_ _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07929__A1 cpu.timer_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07971_ _02793_ _03259_ cpu.needs_timer_interrupt _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09710_ cpu.last_addr\[1\] cpu.ROM_addr_buff\[1\] cpu.last_addr\[0\] _04710_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06922_ _02207_ _02388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_87_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05168__A1 _00672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09641_ _04449_ _04627_ _04643_ _04439_ _04644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06853_ _00763_ _00855_ _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05804_ _01272_ _01274_ _01276_ _01277_ _01278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09572_ _03696_ _04531_ _04577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06784_ _02246_ _02249_ _02250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05263__S1 _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05735_ _01208_ _01209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_77_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08523_ cpu.orig_PC\[7\] _03668_ _03694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_26_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06668__A1 _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08454_ cpu.orig_IO_addr_buff\[0\] _03643_ _03644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05666_ _01117_ _01139_ _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_37_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08385_ cpu.uart.receive_div_counter\[4\] _03588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05597_ _01005_ _01070_ _01071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07405_ _02532_ _02818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_9_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09606__A1 _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07336_ _02764_ _02765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06445__I _01913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07093__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09006_ _03724_ _04070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07267_ _01166_ _02705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_103_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06218_ _00748_ _00951_ _01689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07198_ _02454_ _02587_ _02648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06149_ _01617_ _01620_ _01621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07276__I _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09908_ _04039_ _04872_ _04876_ _04875_ _00518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09839_ _04821_ _04822_ _04823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_29_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06659__A1 _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10614_ _00486_ clknet_leaf_89_wb_clk_i cpu.PC\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10545_ _00418_ clknet_leaf_30_wb_clk_i cpu.timer_div\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10476_ _00349_ clknet_leaf_101_wb_clk_i cpu.pwm_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05634__A2 _00986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_63_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05493__S1 _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05520_ _00599_ _00600_ _00994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_74_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09350__B _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05451_ _00881_ _00903_ _00928_ _00929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08170_ _03420_ _03421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_55_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06265__I _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07075__A1 _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07121_ _02552_ _02576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05382_ _00826_ _00861_ _00862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_112_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07052_ _02512_ _02513_ _00628_ _02514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_70_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06003_ _00895_ _00897_ _01476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07954_ _03239_ cpu.timer\[0\] _02723_ _01463_ _03242_ _03243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_07885_ cpu.spi.dout\[5\] _03174_ _03175_ cpu.spi.data_in_buff\[5\] _03177_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06905_ _02192_ _02211_ _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09624_ _04624_ _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05236__S1 _00734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06836_ _02219_ _02279_ _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_37_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_37_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_37_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09555_ _02653_ _01144_ _04539_ _04540_ _04561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_06767_ _02188_ _02189_ _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05718_ _01191_ _01192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08506_ _03680_ _03681_ _00311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09486_ _04427_ _04481_ _04494_ _04351_ _04495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06698_ _02162_ _02163_ _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_108_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08437_ _02890_ _03629_ _03630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05649_ _01119_ _00986_ _01122_ _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_102_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08368_ _02918_ _02931_ _03574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_92_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08299_ _03408_ _00239_ _03525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07319_ _01915_ _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10330_ _00203_ clknet_leaf_46_wb_clk_i cpu.spi.div_counter\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05616__A2 _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10261_ _00134_ clknet_leaf_115_wb_clk_i cpu.regs\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10192_ _00069_ clknet_leaf_15_wb_clk_i cpu.toggle_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08318__A1 _03407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10125__A1 _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09118__I0 cpu.ROM_addr_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05855__A2 _01328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput14 io_in[21] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_107_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput25 rst_n net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_25_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10528_ _00401_ clknet_leaf_25_wb_clk_i cpu.timer_capture\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08557__A1 _01413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10459_ _00332_ clknet_leaf_12_wb_clk_i cpu.toggle_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05429__I _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09109__I0 _00690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07670_ _02098_ _03019_ _00137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06621_ _02084_ _02085_ _02087_ _02088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09340_ _02848_ _04298_ _04351_ _04352_ _04353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06552_ _01142_ _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07296__A1 _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09271_ _04266_ _04270_ _04271_ _04283_ _04285_ _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_05503_ _00822_ _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09285__A2 _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08222_ cpu.uart.div_counter\[4\] _03460_ _03464_ _03465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06483_ _01395_ _01947_ _01948_ _01614_ _01950_ _01951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_23_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05113__B _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05434_ _00909_ _00911_ _00912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_31_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08153_ _03389_ _03406_ _03407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05365_ _00007_ _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08084_ _03346_ _00224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07104_ _02488_ _02118_ _02561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07035_ _02496_ _00574_ _02115_ _02497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_70_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05296_ _00775_ _00795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08986_ _02787_ _04034_ _04054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07220__A1 _01924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06023__A2 _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input33_I sram_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07937_ _02046_ _02756_ _02751_ _01992_ _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__10107__A1 _04454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07868_ _03164_ _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08720__A1 _02800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05129__A4 _00637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09607_ _04383_ _04604_ _04611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06819_ _02252_ _02258_ _02285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_07799_ _01643_ _03100_ _03105_ _00180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09538_ _04529_ _04426_ _04545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09469_ _04324_ _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_54_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10313_ _00186_ clknet_leaf_2_wb_clk_i cpu.regs\[2\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_115_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10244_ _00117_ clknet_leaf_120_wb_clk_i cpu.regs\[11\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10175_ _00052_ clknet_leaf_22_wb_clk_i cpu.timer_capture\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05150_ cpu.instr_cycle\[2\] _00658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__08778__A1 cpu.timer_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05159__I _00666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05081_ cpu.base_address\[4\] _00592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_100_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08840_ _02756_ _03932_ _03919_ _03939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05983_ _01016_ _01035_ _01456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08771_ cpu.timer_top\[11\] _03877_ _03882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07722_ cpu.regs\[7\]\[7\] _03055_ _03056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07653_ _02981_ _03005_ _03012_ _00127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06604_ _01362_ _02070_ _02071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09323_ cpu.orig_PC\[1\] _04099_ _04336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07584_ _01102_ _02100_ _02965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07269__A1 _02706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06535_ _01289_ _02002_ _02003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09254_ _02669_ _01290_ _01166_ _01280_ _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06466_ _01842_ _01934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_90_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08205_ _03379_ _03442_ _03449_ _03450_ _00241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09185_ cpu.last_addr\[4\] _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06492__A2 _00976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05417_ cpu.regs\[4\]\[2\] cpu.regs\[5\]\[2\] cpu.regs\[6\]\[2\] cpu.regs\[7\]\[2\]
+ _00829_ _00891_ _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_08136_ cpu.uart.div_counter\[7\] _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_71_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06453__I _01921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06397_ _01852_ _01864_ _01374_ _01866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05348_ _00827_ _00828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08067_ cpu.spi.data_in_buff\[0\] _03337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05279_ _00737_ _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07018_ cpu.startup_cycle\[6\] _02480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_110_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_52_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_52_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08969_ cpu.timer_div\[1\] _04035_ _04041_ _04015_ _04042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06180__A1 net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08472__A3 _03638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05688__B _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06363__I _00785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10227_ _00100_ clknet_leaf_0_wb_clk_i cpu.regs\[13\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08932__A1 cpu.timer_capture\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05746__B2 net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10158_ _00035_ clknet_leaf_99_wb_clk_i cpu.regs\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10089_ _01310_ _04100_ _05018_ _05019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_71_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06320_ _01693_ _01789_ _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06251_ _00722_ _00730_ _00902_ _01722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__07369__I _02790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05202_ _00692_ _00705_ _00706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_115_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06182_ _01652_ _01203_ _00999_ _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_52_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05133_ _00635_ _00638_ _00641_ _00642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_111_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09941_ _02779_ _04887_ _04898_ _00529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_96_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07974__A2 _01174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05064_ cpu.mem_cycle\[5\] cpu.mem_cycle\[4\] cpu.mem_cycle\[3\] cpu.mem_cycle\[2\]
+ _00575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__08702__B _03709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09872_ _04846_ _04847_ _00511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08923__A1 cpu.timer_capture\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05737__A1 _00993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08823_ cpu.timer_capture\[4\] _03902_ _03923_ _03924_ _03925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05966_ net7 _01073_ _01197_ _01439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08754_ cpu.timer_div_counter\[5\] _03868_ _03871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07705_ _03042_ _03039_ _03044_ _00147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_68_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08685_ _03822_ _00622_ _00349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05897_ _01308_ _01370_ _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_67_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07636_ _02985_ _03000_ _03001_ _00121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07567_ cpu.regs\[13\]\[1\] _02953_ _02955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06518_ _01983_ _01984_ _01985_ _01986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_76_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09306_ _02555_ _04319_ _04320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09100__A1 _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07498_ cpu.uart.receive_div_counter\[3\] _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09237_ _02728_ _04247_ _04253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07279__I _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06449_ _01479_ _01917_ _01589_ _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07662__A1 _01407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09168_ _04198_ _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08119_ net68 _03373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09099_ _02549_ _04143_ _04147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06217__A2 _00951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output64_I net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10012_ _04946_ _04947_ _04948_ _02507_ _04949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__08914__A1 _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07717__A2 _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05262__I _00762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07653__A1 _02981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08241__C _03479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06042__B _01395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05719__A1 _01039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08905__A1 _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05820_ _01293_ _01294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_19_Left_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05751_ _01224_ _01225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_106_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05172__I _00678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08470_ _03654_ _03655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05682_ cpu.regs\[12\]\[7\] cpu.regs\[13\]\[7\] cpu.regs\[14\]\[7\] cpu.regs\[15\]\[7\]
+ _00827_ _00890_ _01156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07421_ _02829_ _02830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07352_ _02776_ _02765_ _02777_ _02772_ _00061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06303_ _01772_ _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_18_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07283_ _02713_ _02715_ _02716_ _02719_ _02720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_28_Left_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09022_ cpu.uart.divisor\[15\] _04074_ _04080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06234_ _01704_ _01705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06165_ _00981_ _01637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_4_3_0_wb_clk_i clknet_0_wb_clk_i clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_05116_ _00624_ _00625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06096_ cpu.spi.dout\[2\] _01450_ _01422_ _01567_ _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__05958__A1 cpu.PORTA_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09149__A1 _03701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09924_ _01320_ _01080_ _03897_ _04886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_09855_ cpu.ROM_spi_dat_out\[6\] _04835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08806_ _02729_ _03908_ _03909_ _03910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_37_Left_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09786_ _04771_ _04776_ _04777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_14_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06998_ _02448_ _02449_ _02461_ _00023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_96_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05949_ _01421_ _01422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08737_ _03858_ _03859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09321__A1 _00651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08668_ cpu.toggle_ctr\[10\] _03810_ _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_49_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07619_ cpu.regs\[11\]\[0\] _02991_ _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10630_ _00502_ clknet_leaf_71_wb_clk_i cpu.ROM_spi_dat_out\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08599_ cpu.toggle_ctr\[5\] _03753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_48_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_46_Left_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10561_ _00433_ clknet_leaf_56_wb_clk_i cpu.IO_addr_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10492_ _00365_ clknet_leaf_27_wb_clk_i cpu.timer_div_counter\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08060__A1 _02791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06641__I _02106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_53_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Left_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10112__B _00666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_101_Right_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06088__I _00607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Left_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05720__I _01193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08051__A1 _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_73_Left_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07970_ _03258_ _03259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06921_ _02374_ _02375_ _02385_ _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_TAPCELL_ROW_87_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05168__A2 cpu.needs_interrupt vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08478__I _00677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09640_ _00743_ _04403_ _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07382__I _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06852_ _02312_ _02314_ _02317_ _02318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05803_ _01261_ _01058_ _01277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_09571_ _03696_ _04554_ _04576_ _00481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06783_ _00807_ _00858_ _02248_ _02249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05734_ _01201_ _01207_ _01208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_08522_ _03654_ _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09303__A1 _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08453_ _03640_ _03643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_58_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06668__A2 _02133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05665_ _01124_ _01138_ _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07404_ _02568_ _02817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08384_ _03504_ _03587_ _00283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_92_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05596_ _01020_ _00568_ _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09606__A2 _00880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07335_ _01085_ _02763_ _02764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_21_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07266_ cpu.uart.divisor\[7\] _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_98_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07093__A2 _02543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09005_ cpu.uart.divisor\[9\] _04067_ _04069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06217_ _00749_ _00951_ _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_14_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07197_ _02635_ _02646_ _02647_ _00036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06148_ _01618_ _01619_ _01620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06079_ net41 _01429_ _01077_ _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09907_ net60 _04873_ _04876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07148__A3 _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09838_ _02473_ _04801_ _04822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07292__I _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09769_ _02508_ _04763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_57_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06108__A1 _01277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_1_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09012__I _04065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10613_ _00485_ clknet_leaf_96_wb_clk_i cpu.PC\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10544_ _00417_ clknet_leaf_22_wb_clk_i cpu.timer_div\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07084__A2 _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10475_ _00348_ clknet_leaf_7_wb_clk_i cpu.toggle_ctr\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_118_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_71_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_7_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_7_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06434__I2 cpu.regs\[10\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05450_ _00927_ _00928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05381_ cpu.regs\[12\]\[1\] cpu.regs\[13\]\[1\] cpu.regs\[14\]\[1\] cpu.regs\[15\]\[1\]
+ _00831_ _00836_ _00861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_70_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07120_ _02571_ _02569_ _02572_ _02575_ _00031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_43_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07051_ _02472_ _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_81_Left_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06002_ _00889_ _00893_ _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_93_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07953_ cpu.timer_top\[2\] _03237_ _03242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07884_ _03176_ _00194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06904_ _02265_ _02368_ _02369_ _02370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09623_ cpu.orig_PC\[11\] _04238_ _04434_ _04625_ _04626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06835_ _02296_ _02300_ _02301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09554_ _03122_ _00978_ _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06766_ _02228_ _02230_ _02231_ _02232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05717_ _00607_ _01191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08505_ _02859_ _03674_ _03677_ _03681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09485_ _02621_ _04389_ _04494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06697_ _00771_ _00975_ _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08436_ _03625_ _03626_ _03629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06510__A1 _01975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_77_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_77_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_78_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06456__I _01119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05648_ _01121_ _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08367_ _03573_ _00280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05360__I _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07318_ _00621_ _02749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05579_ cpu.br_rel_dest\[7\] _01053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08298_ cpu.uart.data_buff\[1\] _03524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07249_ _02675_ _02691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05616__A3 _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10260_ _00133_ clknet_leaf_0_wb_clk_i cpu.regs\[0\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06577__A1 cpu.timer_capture\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10191_ _00068_ clknet_leaf_15_wb_clk_i cpu.toggle_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06501__A1 net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05270__I cpu.regs\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput15 io_in[23] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput26 sram_out[0] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10527_ _00400_ clknet_leaf_25_wb_clk_i cpu.timer_capture\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_12_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10458_ _00331_ clknet_leaf_11_wb_clk_i cpu.toggle_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10389_ _00262_ clknet_leaf_52_wb_clk_i cpu.uart.data_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09109__I1 _02831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06620_ _01396_ _02064_ _02086_ _01615_ _02087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_99_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06551_ _01408_ _02017_ _02018_ _00019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05502_ _00977_ net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09270_ _01830_ _01146_ _04268_ _04284_ _04285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_06482_ _01937_ _01511_ _01914_ _01949_ _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_08221_ _03445_ _03464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05433_ cpu.regs\[12\]\[3\] cpu.regs\[13\]\[3\] cpu.regs\[14\]\[3\] cpu.regs\[15\]\[3\]
+ _00828_ _00910_ _00911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08705__B _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08245__A1 _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08152_ _03395_ _03398_ _03402_ _03405_ _03406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_43_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05364_ cpu.regs\[8\]\[0\] cpu.regs\[9\]\[0\] cpu.regs\[10\]\[0\] cpu.regs\[11\]\[0\]
+ _00832_ _00837_ _00844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_08083_ cpu.spi.data_in_buff\[6\] _03333_ _03342_ cpu.spi.data_in_buff\[7\] _03346_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09993__A1 _02690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07103_ _02544_ _02560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05295_ _00774_ _00794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_113_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07034_ cpu.mem_cycle\[3\] cpu.mem_cycle\[2\] _02496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_43_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08440__B _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08985_ _04053_ _00418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07220__A2 _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07936_ _03202_ _03205_ _03216_ _03224_ _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA_input26_I sram_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05355__I _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10107__A2 _05036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07867_ _02531_ _03163_ _03164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06818_ _02281_ _02282_ _02283_ _02284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09606_ _03146_ _00880_ _04609_ _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_07798_ cpu.regs\[3\]\[2\] _03103_ _03105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_104_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09537_ _04458_ _04542_ _04543_ _04347_ _04544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06749_ _02187_ _02214_ _02215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09468_ _04477_ _00477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08419_ cpu.uart.receive_div_counter\[10\] _03613_ _03615_ _03611_ _03616_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09399_ _04410_ _04411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output94_I net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10312_ _00185_ clknet_leaf_104_wb_clk_i cpu.regs\[3\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_115_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08539__A2 _03643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10243_ _00116_ clknet_leaf_119_wb_clk_i cpu.regs\[11\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10174_ _00051_ clknet_leaf_21_wb_clk_i cpu.timer_capture\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08711__A2 _02674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08576__I cpu.toggle_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05080_ cpu.base_address\[5\] _00591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_110_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05764__A2 _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05982_ cpu.timer_div\[1\] _01422_ _01452_ _01454_ _01455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_08770_ _02804_ _03876_ _03881_ _03879_ _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05175__I cpu.ROM_OEB vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06961__A1 _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07721_ _03038_ _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10461__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07652_ cpu.regs\[10\]\[5\] _03003_ _03012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06603_ _02067_ _02069_ _02070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07583_ _01405_ _02964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_87_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09322_ _04334_ _04335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06534_ _00644_ _02001_ _02002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09253_ _01585_ _02684_ _04267_ _04268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06465_ _01930_ _01932_ _01933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08204_ _02809_ _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09184_ _04193_ _04210_ _04211_ _00459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_90_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06396_ _01838_ _01864_ _01865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05416_ _00894_ _00842_ _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08135_ _03377_ _03381_ _03385_ _03388_ _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05347_ _00004_ _00827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_71_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08066_ _03335_ _03336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05278_ _00776_ _00777_ _00750_ _00778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07017_ _02478_ _02479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05452__A1 _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09194__A2 _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06401__B1 _01869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08968_ _04039_ _04040_ _04041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08899_ _01254_ _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07919_ cpu.timer_top\[10\] _03207_ _03208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_79_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05813__I _00984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_21_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_21_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_66_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10016__B2 cpu.ROM_OEB vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07475__I cpu.uart.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10226_ _00099_ clknet_leaf_0_wb_clk_i cpu.regs\[13\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07196__A1 _02433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10157_ _00034_ clknet_leaf_99_wb_clk_i cpu.regs\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10088_ _00859_ _04240_ _05010_ _05012_ _05017_ _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__05723__I _01196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06250_ _01710_ _01711_ _01714_ _01720_ _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_115_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10007__A1 cpu.ROM_spi_mode vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09948__A1 _02790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05201_ cpu.regs\[8\]\[1\] cpu.regs\[9\]\[1\] cpu.regs\[10\]\[1\] cpu.regs\[11\]\[1\]
+ _00683_ _00685_ _00705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06181_ net62 _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05132_ _00639_ _00640_ _00641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_25_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09940_ net55 _04888_ _02682_ _04898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05063_ _00573_ _00574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_115_Right_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06503__B cpu.PORTA_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07385__I _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09871_ cpu.ROM_spi_cycle\[2\] _04844_ _04290_ _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07187__A1 _02637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08822_ _02546_ _03924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05965_ net22 _01000_ _01229_ _01437_ _01438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_08753_ cpu.timer_div_counter\[5\] _03868_ _03870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07704_ cpu.regs\[7\]\[1\] _03043_ _03044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08684_ cpu.pwm_counter\[0\] _03822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05896_ _01357_ _01370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07635_ cpu.regs\[11\]\[7\] _03000_ _03001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07566_ _01407_ _02952_ _02954_ _00098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06517_ cpu.spi.dout\[6\] _01450_ _01647_ _01985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09305_ _04293_ _04313_ _04318_ _04319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07497_ _02893_ _02894_ _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09236_ _00672_ _04245_ _04252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06448_ _01579_ _01901_ _01916_ _01917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09167_ _04197_ _04198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06379_ _01835_ _01846_ _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08118_ _03370_ _03353_ _03372_ _00232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09098_ _04146_ _00438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07414__A2 _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_43_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08049_ _02776_ _03308_ _03321_ _03323_ _00212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_3_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05276__I1 _00772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05976__A2 _01174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10011_ _04778_ _02482_ _04948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output57_I net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06639__I _02104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_82_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10209_ _00082_ clknet_leaf_7_wb_clk_i _00000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05750_ _01223_ _01195_ _01005_ _01224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__09353__C _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06549__I _02016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05681_ _00840_ _01154_ _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_85_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07420_ _02828_ _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07351_ cpu.timer_top\[3\] _02766_ _02777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06302_ _01770_ _01771_ _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07282_ _02717_ _02718_ _02719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09021_ _02701_ _04073_ _04079_ _04078_ _00428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06233_ _01690_ _01704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06164_ _01629_ _01631_ _01632_ _01634_ _01635_ _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_25_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05115_ _00623_ _00624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05407__A1 _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06095_ _01547_ _01564_ _01565_ _01566_ _01567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__06080__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05628__I _01101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09923_ _02706_ _04879_ _04885_ _04882_ _00524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09854_ _04834_ _00506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_4_12_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08805_ _03258_ _03909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09785_ _02476_ _02506_ _04776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06997_ net19 _02132_ _02450_ _02460_ _02419_ _02461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05948_ _01002_ _01250_ _01027_ _01421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08736_ _03196_ _03858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08667_ _03805_ _03810_ _03811_ _00342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05879_ _01352_ _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07618_ _02988_ _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08598_ cpu.toggle_ctr\[1\] _03750_ _01167_ _03751_ _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_24_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07549_ _01644_ _02939_ _02943_ _00092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_101_Left_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10560_ _00432_ clknet_leaf_56_wb_clk_i cpu.IO_addr_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07635__A2 _03000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09219_ _04087_ _04236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10491_ _00364_ clknet_leaf_20_wb_clk_i cpu.pwm_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07399__A1 cpu.toggle_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08849__I _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06374__A2 _01841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05273__I cpu.regs\[2\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07323__A1 cpu.timer_capture\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06126__A2 _01380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10689_ _00561_ clknet_leaf_5_wb_clk_i cpu.regs\[15\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05448__I _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06920_ _02374_ _02375_ _02385_ _02386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06851_ _02315_ _00858_ _02316_ _02317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06279__I cpu.uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09570_ _04367_ _04572_ _04573_ _04575_ _04576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05802_ _01275_ _01273_ _01276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06782_ _02245_ _02247_ _02248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_89_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05733_ _01206_ _01207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08521_ _03691_ _03692_ _00315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09303__A2 _04315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08452_ _03641_ _03642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07403_ _02815_ _02796_ _02816_ _02810_ _00073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__05876__A1 _01104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05664_ _01125_ _01132_ _01135_ _01137_ _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_08383_ cpu.uart.receive_div_counter\[3\] _03576_ _03586_ _03571_ _03587_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05595_ _00602_ _01069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_58_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07334_ _02761_ _02762_ _02763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_21_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07265_ _02703_ _00048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_98_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09004_ _03840_ _04066_ _04068_ _03853_ _00422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_84_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06216_ _01504_ _01608_ _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08578__B1 _01275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07196_ _02433_ _02633_ _02647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06147_ _01350_ _01526_ _01619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06078_ _01548_ _01081_ _01432_ _01549_ _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_09906_ _03840_ _04872_ _04874_ _04875_ _00517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__07573__I _02951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09837_ _04804_ _04821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09768_ _04752_ _04758_ _04761_ _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_57_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08719_ cpu.pwm_top\[1\] _03847_ _03848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09699_ cpu.last_addr\[6\] cpu.last_addr\[5\] _04698_ _04699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06108__A2 _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05867__A1 _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06659__A3 _01337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10612_ _00484_ clknet_leaf_93_wb_clk_i cpu.PC\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10543_ _00416_ clknet_leaf_22_wb_clk_i cpu.timer_div\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06292__A1 cpu.timer_capture\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10474_ _00347_ clknet_leaf_7_wb_clk_i cpu.toggle_ctr\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_118_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08033__A2 _01424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09781__A2 _04771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06044__A1 _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06434__I3 cpu.regs\[11\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05380_ _00822_ _00859_ _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07050_ cpu.spi_clkdiv _02512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05086__A2 cpu.br_rel_dest\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06001_ _01066_ _01474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08024__A2 _03164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07952_ _03232_ _03235_ _03238_ _03240_ _03241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07393__I _02809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07535__A1 _00620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07883_ cpu.spi.dout\[4\] _03174_ _03175_ cpu.spi.data_in_buff\[4\] _03176_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06903_ _02213_ _02237_ _02369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09622_ _04557_ _04624_ _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06834_ _02297_ _00857_ _02299_ _02300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09553_ _04557_ _04556_ _04558_ _04559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08504_ cpu.orig_PC\[2\] _03672_ _03680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_54_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09288__A1 cpu.Z vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06765_ _02226_ _02227_ _02231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05716_ cpu.spi.dout\[0\] _01189_ _01184_ _01190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_66_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09484_ _04385_ _04491_ _04492_ _04493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06696_ _02159_ _02161_ _02162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08435_ _03624_ _03628_ _00293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05647_ _01120_ _01092_ _01097_ _00878_ _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08366_ _03569_ _03571_ _03572_ _02708_ _03573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_58_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07317_ _02727_ _02748_ _00055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05578_ _00645_ _00649_ _01052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_116_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06274__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08297_ _03522_ _03523_ _00260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_46_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_46_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_104_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07248_ _00926_ _02690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_33_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09212__A1 _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07179_ _02592_ _02630_ _02614_ _02631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10190_ _00067_ clknet_leaf_15_wb_clk_i cpu.toggle_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput16 io_in[26] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput27 sram_out[1] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10526_ _00399_ clknet_leaf_25_wb_clk_i cpu.timer_capture\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10457_ _00330_ clknet_leaf_12_wb_clk_i cpu.toggle_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10388_ _00261_ clknet_leaf_51_wb_clk_i cpu.uart.data_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08190__A1 _03407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06550_ cpu.regs\[9\]\[6\] _01142_ _02018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_114_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05501_ _00957_ _00964_ _00976_ _00977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06481_ _01389_ _01914_ _00641_ _01949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08220_ cpu.uart.div_counter\[4\] _03456_ _03462_ _03444_ _03463_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05432_ _00833_ _00910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08151_ _02885_ cpu.uart.div_counter\[15\] _03403_ _02903_ _03404_ _03405_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_71_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07388__I _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09442__A1 _02315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05363_ _00842_ _00843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08082_ _03345_ _00223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07102_ _02559_ _00029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05294_ _00779_ _00792_ _00707_ _00793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07033_ _02493_ _02490_ _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_30_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06008__A1 _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09745__A2 _04731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08984_ cpu.timer_div\[5\] _04046_ _04052_ _04050_ _04053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07935_ _03220_ _03221_ _03223_ _03224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07866_ _03161_ cpu.spi.counter\[2\] cpu.spi.counter\[4\] _03162_ _03163_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_97_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09605_ _04585_ _04608_ _04609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_39_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input19_I io_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07797_ _01542_ _03100_ _03104_ _00179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06817_ _02278_ net117 _02283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_104_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09536_ _04489_ _04533_ _04543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06748_ cpu.regs\[1\]\[3\] _00942_ _02214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_78_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09467_ _02605_ _04445_ _04475_ _04476_ _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08418_ _02910_ _03614_ _03615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_109_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06679_ _00724_ _01927_ _02145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09398_ _01287_ _04410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08349_ cpu.uart.receive_buff\[3\] _03555_ _03557_ cpu.uart.receive_buff\[4\] _03561_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_80_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09433__A1 _02861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07995__A1 _03262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10311_ _00184_ clknet_leaf_105_wb_clk_i cpu.regs\[3\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_115_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output87_I net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05470__A2 _00946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10242_ _00115_ clknet_leaf_120_wb_clk_i cpu.regs\[11\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10173_ _00050_ clknet_leaf_21_wb_clk_i cpu.timer_capture\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08806__B _03909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08525__C _03695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10509_ _00382_ clknet_leaf_23_wb_clk_i cpu.timer\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05981_ _01422_ _01453_ _01454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07720_ _03053_ _03040_ _03054_ _00152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07651_ _02977_ _03005_ _03011_ _00126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07582_ _02098_ _02958_ _02963_ _00105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06602_ _01936_ _01914_ _02068_ _02069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10030__C _02818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06533_ _00663_ _02000_ _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09321_ _00651_ _04100_ _04334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_34_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09663__A1 _04361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06477__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09252_ _00951_ _00946_ _00976_ _02021_ _04267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_06464_ _01837_ _01839_ _01931_ _01932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09183_ cpu.ROM_addr_buff\[3\] _04206_ _04211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08203_ _03391_ _03448_ _03379_ _03449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06395_ _01815_ _01853_ _01864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05415_ cpu.regs\[0\]\[2\] cpu.regs\[1\]\[2\] cpu.regs\[2\]\[2\] cpu.regs\[3\]\[2\]
+ _00830_ _00835_ _00894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_08134_ _02880_ cpu.uart.div_counter\[13\] _03386_ cpu.uart.divisor\[11\] _03387_
+ _03388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_90_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05346_ _00825_ _00826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07977__A1 _03262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08065_ _03283_ _03333_ _03335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_33_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05277_ cpu.regs\[4\]\[5\] cpu.regs\[5\]\[5\] cpu.regs\[6\]\[5\] cpu.regs\[7\]\[5\]
+ _00774_ _00775_ _00777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07016_ _02477_ cpu.startup_cycle\[0\] _02478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05452__A2 _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06401__A1 net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05204__A2 _00704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08967_ _04033_ _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08898_ _03985_ _03988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07918_ cpu.timer\[10\] _03207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_07849_ _02410_ _03147_ _03120_ _03148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__07901__A1 cpu.timer_div\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07901__B2 _01546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09519_ _02556_ _04510_ _04526_ _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_61_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_61_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_93_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09301__I _04314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09406__A1 cpu.PC\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10225_ _00098_ clknet_leaf_1_wb_clk_i cpu.regs\[13\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08393__B2 _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10156_ _00033_ clknet_leaf_100_wb_clk_i cpu.br_rel_dest\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07491__I _02891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10087_ _04082_ _05015_ _05016_ _05017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_57_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08448__A2 _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05200_ cpu.regs\[12\]\[1\] cpu.regs\[13\]\[1\] cpu.regs\[14\]\[1\] cpu.regs\[15\]\[1\]
+ _00684_ _00686_ _00704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_25_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06180_ net42 _01212_ _01434_ _01651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_53_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05131_ cpu.base_address\[2\] _00640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05062_ cpu.mem_cycle\[1\] cpu.mem_cycle\[0\] _00573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07666__I _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09870_ cpu.ROM_spi_cycle\[2\] _04844_ _04846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_96_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08821_ _03231_ _03918_ _03895_ _03922_ _03923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09881__I net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_117_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05964_ _01431_ _01433_ _01435_ _01436_ _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_08752_ _03863_ _03868_ _03869_ _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08683_ _03742_ _03821_ _03790_ _00348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07703_ _03037_ _03043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07634_ _02989_ _03000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05895_ _01310_ _01353_ _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07565_ cpu.regs\[13\]\[0\] _02953_ _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07496_ _02885_ cpu.uart.receive_div_counter\[15\] _02888_ _02896_ _02897_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06516_ cpu.spi.divisor\[6\] _01547_ _01189_ _01984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09304_ _04293_ _04317_ _04318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09235_ _04246_ _04250_ _04251_ _00470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06447_ _00961_ _01294_ _01302_ _01915_ _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_17_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09166_ _00609_ _04196_ _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06378_ _01835_ _01846_ _01847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06870__A1 _00726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08117_ cpu.uart.dout\[7\] _03351_ _03371_ _03372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05329_ cpu.PORTA_DDR\[4\] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_71_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09097_ _00978_ _04142_ _04144_ _04145_ _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_44_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07414__A3 _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08048_ cpu.spi.data_out_buff\[2\] _03322_ _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05425__A2 _00887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06622__A1 _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05276__I2 _00773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10010_ _02496_ _02116_ _04733_ _04947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09999_ cpu.PORTA_DDR\[5\] _04937_ _04940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_99_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08127__B2 _02679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09875__A1 _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09031__I _04087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05664__A2 _01132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10208_ _00081_ clknet_leaf_103_wb_clk_i cpu.regs\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05975__I0 _01423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10139_ _00016_ clknet_leaf_121_wb_clk_i cpu.regs\[9\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09866__A1 _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05680_ cpu.regs\[8\]\[7\] cpu.regs\[9\]\[7\] cpu.regs\[10\]\[7\] cpu.regs\[11\]\[7\]
+ _00917_ _01153_ _01154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_85_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07350_ _02775_ _02776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_85_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06301_ _00970_ _00972_ _01771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09020_ cpu.uart.divisor\[14\] _04074_ _04079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_72_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07281_ _02714_ _02718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06232_ _01701_ _01702_ _01703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_25_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06163_ _00907_ _01340_ _01372_ _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_25_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05114_ _00585_ _00623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06604__A1 _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05407__A2 _00874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06094_ _01449_ _01566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09922_ net67 _04880_ _04885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09853_ cpu.ROM_spi_dat_out\[5\] _04807_ _04833_ _04829_ _04834_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09784_ _02476_ _04773_ _04775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08804_ _02717_ _02723_ _03907_ _03908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_08735_ _02791_ _03856_ _03857_ _02786_ _00364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06996_ _02452_ _02453_ _02459_ _02460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__09857__B2 _04771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05947_ _01419_ _01420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08666_ cpu.toggle_ctr\[9\] _03808_ _03811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10202__D _00075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05878_ _01350_ _01351_ _01352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08597_ cpu.toggle_ctr\[0\] _03751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09609__A1 _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07617_ _02989_ _02990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07548_ cpu.regs\[14\]\[2\] _02940_ _02943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06408__C _01225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09085__A2 _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07479_ _01883_ _02880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09218_ _00667_ _04234_ _04235_ _00469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10490_ _00363_ clknet_leaf_17_wb_clk_i cpu.pwm_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09149_ _03701_ _04063_ _04183_ _04184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05582__A1 _01051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08520__A1 _02637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08814__B _03912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06834__A1 _02297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10688_ _00560_ clknet_leaf_5_wb_clk_i cpu.regs\[15\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09000__A2 _03712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06850_ _02312_ _02314_ _02316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05801_ cpu.toggle_top\[8\] _01275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_93_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06781_ _00798_ _00869_ _02247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05732_ _00662_ _01147_ _01204_ _01205_ _01206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_08520_ _02637_ _03686_ _03689_ _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08451_ _03640_ _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05663_ _00987_ _01136_ _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_07402_ _02053_ _02797_ _02816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08382_ _02899_ _03582_ _03586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05594_ _01050_ _01056_ _01067_ _01068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_9_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07333_ _01147_ _01282_ _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_18_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07264_ cpu.uart.divisor\[6\] _02689_ _02702_ _02687_ _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_45_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_118_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_118_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_33_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09003_ _02891_ _04067_ _04068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06215_ _01646_ _01485_ _01685_ _01098_ _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_103_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07195_ _02587_ _02645_ _02646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05639__I _01112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06146_ _01487_ _00718_ _01618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07250__A1 _02690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06077_ _01171_ _01024_ _01083_ cpu.PORTA_DDR\[2\] _01549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_09905_ _04077_ _04875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07854__I cpu.PC\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09836_ _04820_ _00502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09767_ _04759_ _04760_ _04761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_57_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06979_ _02431_ _02443_ _02444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_29_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09698_ _04212_ _04697_ _04698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08718_ _03841_ _03847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_107_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08649_ cpu.toggle_ctr\[4\] _03797_ _03799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_1_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10611_ _00483_ clknet_leaf_93_wb_clk_i cpu.PC\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10542_ _00415_ clknet_leaf_50_wb_clk_i cpu.timer_div\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08569__A1 _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10473_ _00346_ clknet_leaf_6_wb_clk_i cpu.toggle_ctr\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_118_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08033__A3 _03310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08809__B _03912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08528__C _03695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09297__A2 _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08263__C _03479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06000_ _01410_ _01412_ _01472_ _01067_ _01473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_88_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07951_ _03239_ cpu.timer\[0\] cpu.timer\[1\] _01463_ _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07674__I _03020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06902_ _02290_ _02366_ _02367_ _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__10119__A1 _01406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07882_ _03168_ _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08732__A1 _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06833_ _02295_ _02298_ _02299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09621_ _03152_ _04623_ _04624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09552_ cpu.orig_PC\[8\] _04089_ _04558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06764_ _02218_ _02229_ _02230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05715_ _01188_ _01189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08503_ _02848_ _03651_ _03679_ _03653_ _00310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_54_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05922__I _01395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09483_ _04377_ _04481_ _04492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06695_ _00761_ _01928_ _02161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08434_ cpu.uart.receive_div_counter\[13\] _03613_ _03627_ _03583_ _03628_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05143__B _00651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05646_ cpu.br_rel_dest\[2\] _01120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08365_ _03569_ _02920_ _03572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05577_ _00991_ _01051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_46_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07316_ cpu.timer_capture\[5\] _02738_ _02747_ _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08296_ _03410_ _03519_ _02793_ cpu.uart.counter\[3\] _03523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_6_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06274__A2 _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07247_ _02675_ _02689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07178_ _02134_ _02630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06129_ _00722_ _00730_ _01600_ _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06026__A2 _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_86_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_86_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08971__A1 _00903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05785__A1 cpu.timer_capture\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_15_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_15_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_6_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09819_ _04804_ _04805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09732__C _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08723__A1 _03849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06663__I cpu.regs\[2\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput17 io_in[28] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput28 sram_out[2] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10525_ _00398_ clknet_leaf_26_wb_clk_i cpu.timer_capture\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10456_ _00329_ clknet_leaf_12_wb_clk_i cpu.toggle_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_20_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10387_ _00260_ clknet_leaf_51_wb_clk_i cpu.uart.counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08190__A2 _03436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06480_ _01930_ _01948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05500_ _00975_ _00976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_74_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05431_ _00823_ _00909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08150_ _02885_ cpu.uart.div_counter\[15\] cpu.uart.div_counter\[13\] _02880_ _03404_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_43_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07101_ _02556_ _02541_ _02558_ _02547_ _02559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05362_ _00841_ _00842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08081_ cpu.spi.data_in_buff\[5\] _03340_ _03342_ cpu.spi.data_in_buff\[6\] _03345_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05293_ cpu.regs\[8\]\[6\] cpu.regs\[9\]\[6\] cpu.regs\[10\]\[6\] cpu.regs\[11\]\[6\]
+ _00788_ _00789_ _00792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_113_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07032_ _02492_ _02493_ _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_clkbuf_leaf_23_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05189__I _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08983_ _02698_ _04034_ _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07934_ _03206_ cpu.timer\[8\] _03222_ _03223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07865_ cpu.spi.counter\[0\] cpu.spi.counter\[1\] _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09604_ _04586_ _04589_ _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_39_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07796_ cpu.regs\[3\]\[1\] _03103_ _03104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06816_ _02273_ _02275_ _02282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07072__C _02533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09535_ _04529_ _01110_ _04541_ _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06747_ _02170_ _02191_ _02213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_65_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09466_ _04410_ _04476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06678_ cpu.regs\[1\]\[1\] _01927_ _02144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_19_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10210__D _00083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08417_ _02882_ _03605_ _03601_ _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA_clkbuf_leaf_62_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05629_ _00648_ _01103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07692__A1 _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09397_ _04402_ _04371_ _04406_ _04408_ _04409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08348_ _03560_ _00274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09433__A2 _04443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08279_ _03499_ _03439_ _03509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07444__A1 _02639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07995__A2 _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10310_ _00183_ clknet_leaf_105_wb_clk_i cpu.regs\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_15_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10241_ _00114_ clknet_leaf_119_wb_clk_i cpu.regs\[11\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08944__A1 _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10172_ _00049_ clknet_leaf_40_wb_clk_i cpu.uart.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05758__A1 _01222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05930__A1 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09672__A2 _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07435__A1 _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10508_ _00381_ clknet_4_6_0_wb_clk_i cpu.timer\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10439_ _00312_ clknet_leaf_84_wb_clk_i cpu.orig_PC\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_107_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07738__A2 _03060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06410__A2 _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05980_ cpu.spi.dout\[1\] _01189_ _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08163__A2 _01424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07650_ cpu.regs\[10\]\[4\] _03007_ _03011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05472__I _00948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07581_ cpu.regs\[13\]\[7\] _02959_ _02963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06601_ _01947_ _01932_ _02068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06532_ _01204_ _02000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09320_ _02340_ _04328_ _04332_ _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_34_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09251_ _01829_ _01146_ _04265_ _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06517__B _01647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08202_ _03443_ _03448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_44_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06463_ _01836_ _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09182_ cpu.last_addr\[3\] _04199_ _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06394_ _01622_ _01844_ _01858_ _01862_ _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_05414_ _00842_ _00892_ _00847_ _00893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08133_ _02889_ cpu.uart.div_counter\[14\] cpu.uart.div_counter\[1\] _02679_ _03387_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_7_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05345_ _00824_ _00825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08064_ _03333_ _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07977__A2 _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07015_ cpu.startup_cycle\[1\] _02477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05988__A1 cpu.timer_capture\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05276_ cpu.regs\[0\]\[5\] _00772_ _00773_ cpu.regs\[3\]\[5\] _00774_ _00775_ _00776_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_113_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08926__A1 _02745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input31_I sram_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08966_ _02722_ _04039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08897_ _01456_ _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07917_ cpu.timer_top\[8\] _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07848_ _03146_ _02409_ _02625_ _03147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05912__A1 _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09518_ _02433_ _04441_ _04410_ _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07779_ _03085_ _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_38_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09449_ cpu.PC\[3\] cpu.br_rel_dest\[3\] _04459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_30_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_30_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_61_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06640__A2 _00583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10224_ _00097_ clknet_leaf_113_wb_clk_i cpu.regs\[14\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10155_ _00032_ clknet_leaf_100_wb_clk_i cpu.br_rel_dest\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10086_ cpu.orig_flags\[0\] _04087_ _05016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09645__A2 _04446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05130_ cpu.base_address\[3\] _00639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_25_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08271__C _03479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05061_ net25 _00572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08820_ _03919_ _03921_ _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05963_ _00998_ _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08751_ cpu.timer_div_counter\[4\] _03866_ _03869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_49_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08682_ cpu.toggle_ctr\[14\] _03818_ _03821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05894_ _01367_ _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07702_ _01541_ _03042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07895__A1 cpu.timer_div\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07633_ _02983_ _02991_ _02999_ _00120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09830__C _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07564_ _02951_ _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06515_ _01981_ _01982_ _01983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07495_ _02889_ _02890_ cpu.uart.receive_div_counter\[8\] _02892_ _02895_ _02896_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_48_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09303_ _02820_ _04315_ _04316_ _04317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09234_ _03503_ _04251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_61_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06446_ _01914_ _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_17_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09165_ _04194_ _04195_ _04196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_90_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08116_ _02681_ _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06377_ _01348_ _01840_ _01845_ _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05328_ cpu.PORTB_DDR\[4\] net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09096_ _04049_ _04145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08047_ _03300_ _03322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05425__A3 _00903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05259_ _00757_ _00759_ _00760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05276__I3 cpu.regs\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09572__A1 _03696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09998_ _04047_ _04936_ _04938_ _04939_ _00545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_08949_ _04020_ _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09312__I _04293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06310__A1 _01779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09563__A1 _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10207_ _00080_ clknet_leaf_99_wb_clk_i cpu.regs\[1\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10138_ _00015_ clknet_leaf_121_wb_clk_i cpu.regs\[9\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10069_ _04753_ _02502_ _04836_ _04813_ _05001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06129__A1 _00722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07629__A1 _02977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07280_ cpu.timer\[0\] _02717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06300_ _00966_ _00968_ _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06231_ _01687_ _01699_ _01361_ _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07677__I _03020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06162_ _01617_ _01633_ _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_13_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06093_ cpu.spi.divisor\[2\] _01547_ _01565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05113_ _00612_ _00617_ _00622_ _00011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07801__A1 _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09921_ _02701_ _04879_ _04884_ _04882_ _00523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09554__A1 _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09852_ _04831_ _04793_ _04805_ _04811_ _04833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09783_ _04772_ _04774_ _00495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08803_ _03197_ _03907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05415__I0 cpu.regs\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09157__I1 _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08734_ cpu.pwm_top\[7\] _03856_ _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06995_ _02456_ _02458_ _02459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05946_ _01248_ _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08665_ cpu.toggle_ctr\[9\] _03808_ _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05877_ _01316_ net90 _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08596_ cpu.toggle_top\[1\] _03750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07616_ _02988_ _02989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_62_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07547_ _01543_ _02939_ _02942_ _00091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_64_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07478_ cpu.uart.receive_div_counter\[5\] _01881_ _02876_ _02877_ _02679_ _02878_
+ _02879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_0_118_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09217_ cpu.ROM_addr_buff\[13\] _04213_ _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06429_ cpu.pwm_top\[5\] _01268_ _01270_ _01898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09148_ _04173_ cpu.regs\[3\]\[2\] _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07587__I _02967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09079_ _01830_ _04123_ _04130_ _04084_ _04131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_15_Left_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output62_I net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09545__B2 _04453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06359__A1 _01408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09751__B _02710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10149__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_24_Left_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07859__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06531__A1 cpu.toggle_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10091__A1 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_33_Left_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10687_ _00559_ clknet_leaf_4_wb_clk_i cpu.regs\[15\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06598__A1 _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05800_ _01273_ _01274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_42_Left_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06780_ _00800_ _00873_ _02245_ _02246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_26_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05731_ _00632_ _00992_ _01205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_26_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08450_ _03639_ _03640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05662_ _01000_ _01068_ _01074_ _01091_ _01136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_08381_ _03579_ _03580_ _03584_ _03585_ _00282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__06522__A1 cpu.timer_capture\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07401_ _02755_ _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07332_ _01149_ _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05593_ _01059_ _01063_ _01066_ _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XPHY_EDGE_ROW_51_Left_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07263_ _02701_ _02691_ _02702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_98_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10082__A1 _01392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08027__A1 _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09002_ _04065_ _04067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06214_ _01306_ _01683_ _01684_ _01313_ _01685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_5_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07194_ _02603_ _02644_ _02645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09775__A1 _02533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08578__A2 _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06145_ _01603_ _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06076_ net81 _01548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09904_ net59 _04873_ _04874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09835_ cpu.ROM_spi_dat_out\[1\] _04806_ _04819_ _04736_ _04820_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09766_ _00580_ _00582_ _04760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08966__I _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06978_ _02442_ _02443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_29_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09697_ cpu.last_addr\[3\] cpu.last_addr\[2\] _04696_ _04697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08717_ _03840_ _03843_ _03845_ _03846_ _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05929_ _01094_ _01403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_107_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08502__A2 _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08648_ _03796_ _03797_ _03798_ _00336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_1_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05390__I _00869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08579_ _03731_ _03732_ _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_76_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10610_ _00482_ clknet_leaf_96_wb_clk_i cpu.PC\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10541_ _00414_ clknet_leaf_22_wb_clk_i cpu.timer_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10472_ _00345_ clknet_leaf_6_wb_clk_i cpu.toggle_ctr\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_118_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09746__B _04251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09518__A1 _02433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_2_0_wb_clk_i clknet_0_wb_clk_i clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__06504__A1 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06807__A2 _00855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_13_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08116__I _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07950_ cpu.timer_top\[0\] _03239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05475__I _00951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06901_ _02239_ _02264_ _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07881_ _03164_ _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06832_ _00762_ _00870_ _02298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09620_ _02410_ _04479_ _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09551_ _04272_ _04557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06763_ _00806_ _00872_ _02217_ _02229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05714_ _01187_ _01188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08502_ cpu.orig_PC\[1\] _03668_ _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_54_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09482_ _04485_ _04488_ _04490_ _04491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06694_ _02145_ _02159_ _02151_ _02152_ _02160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_08433_ _03625_ _03626_ _03627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_52_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05645_ _01118_ _01119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08364_ _03570_ _03571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05576_ _01009_ _01041_ _01044_ _01049_ _01050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_62_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09996__A1 cpu.PORTA_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07315_ _02745_ _02739_ _02740_ _02746_ _02747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_6_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08295_ _03521_ _03522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08026__I _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07246_ _02688_ _00044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07177_ _02587_ _02628_ _02629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_112_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06128_ cpu.br_rel_dest\[2\] _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_06059_ _01500_ _01523_ _01525_ _01527_ _01531_ _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_6_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06982__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09818_ _02517_ _04803_ _04804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09920__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_91_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09749_ _04743_ _04740_ _04745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_55_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_55_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_68_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09987__A1 _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput18 io_in[29] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_107_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput29 sram_out[3] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10524_ _00397_ clknet_leaf_25_wb_clk_i cpu.timer_capture\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10455_ _00328_ clknet_leaf_15_wb_clk_i cpu.toggle_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10386_ _00259_ clknet_leaf_49_wb_clk_i cpu.uart.counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08962__A2 _00586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09911__A1 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05430_ _00907_ _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_55_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05361_ _00840_ _00841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_23_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07100_ _02542_ _02557_ _02558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08080_ _03344_ _00222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_99_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05292_ _00787_ _00790_ _00791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07031_ _02110_ _02112_ _02493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08982_ _04051_ _00417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07933_ cpu.timer_top\[9\] _03198_ _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07864_ cpu.spi.counter\[3\] _03161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09603_ _04557_ _04605_ _04606_ _04607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05519__A2 _00991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06815_ _02278_ _02280_ _02281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05933__I _01406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07795_ _03098_ _03103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_104_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09534_ _04539_ _04540_ _04541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06746_ _02192_ _02211_ _02212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09465_ _02556_ _04448_ _04452_ _04453_ _04474_ _04475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06677_ _00725_ _02008_ _02143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_19_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08416_ _03575_ _03613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05628_ _01101_ _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09396_ _04407_ _04408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07692__A2 _03032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08347_ cpu.uart.receive_buff\[2\] _03555_ _03557_ cpu.uart.receive_buff\[3\] _03560_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05559_ _01001_ _01030_ _01032_ _01033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_116_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08278_ _03507_ _03508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_102_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_102_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07229_ _02673_ _02674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_15_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10240_ _00113_ clknet_leaf_113_wb_clk_i cpu.regs\[12\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06432__C _01277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10171_ _00048_ clknet_leaf_40_wb_clk_i cpu.uart.divisor\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_110_Right_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09315__I _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10019__A1 _00608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09050__I _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_7_Left_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10507_ _00380_ clknet_leaf_11_wb_clk_i cpu.timer_top\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_69_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10438_ _00311_ clknet_leaf_84_wb_clk_i cpu.orig_PC\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07199__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10369_ _00242_ clknet_leaf_32_wb_clk_i cpu.uart.div_counter\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08935__A2 _02755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06849__I _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08163__A3 _03310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07371__A1 _02791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07580_ _02017_ _02958_ _02962_ _00104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06600_ _02064_ _02066_ _02067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06531_ cpu.toggle_top\[14\] _01274_ _01279_ _01999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09250_ _01778_ _00571_ _04239_ _04265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_16_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_0_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_0_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08201_ _03442_ _03447_ _00240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06462_ _00803_ _01929_ _01930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09181_ _04193_ _04208_ _04209_ _00458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06393_ _01615_ _01852_ _01859_ _01812_ _01861_ _01862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05413_ cpu.regs\[8\]\[2\] cpu.regs\[9\]\[2\] cpu.regs\[10\]\[2\] cpu.regs\[11\]\[2\]
+ _00829_ _00891_ _00892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_08132_ cpu.uart.div_counter\[11\] _03386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05344_ _00823_ _00824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08063_ _03299_ _00676_ _03332_ _03333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__08732__C _03853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05275_ _00753_ _00775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07014_ cpu.startup_cycle\[3\] _02476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08965_ _01183_ _04035_ _04037_ _04038_ _00413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_110_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07916_ cpu.timer_top\[15\] _03200_ _03204_ cpu.timer_top\[14\] _03205_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA_input24_I io_in[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08896_ _03985_ _03986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07847_ cpu.PC\[10\] _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07778_ _03047_ _03086_ _03091_ _00173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09517_ _04413_ _04315_ _04510_ _04525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06729_ _02160_ _02164_ _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08862__A1 cpu.timer_capture\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09448_ _04304_ _04458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_93_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09379_ _02846_ _04390_ _04391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05220__S0 _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07417__A2 _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09738__C _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output92_I net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10223_ _00096_ clknet_leaf_112_wb_clk_i cpu.regs\[14\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_70_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_70_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_30_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10154_ _00031_ clknet_leaf_100_wb_clk_i cpu.br_rel_dest\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10085_ _04277_ _05013_ _05014_ _04273_ _05015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_97_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05903__A2 _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06092__A1 cpu.spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05060_ _00570_ cpu.br_rel_dest\[6\] _00571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05962_ net60 _01434_ _01435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08750_ cpu.timer_div_counter\[4\] _03866_ _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_49_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08681_ _03790_ _03820_ _00347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05893_ _00589_ _01366_ _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07701_ _03034_ _03039_ _03041_ _00146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07632_ cpu.regs\[11\]\[6\] _02989_ _02999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09302_ _02830_ _04314_ _04316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09097__A1 _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07563_ _02951_ _02952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06514_ cpu.uart.dout\[6\] _01192_ _01665_ _01982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07494_ _02893_ _02894_ _02895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_36_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09233_ cpu.orig_flags\[3\] _04247_ _04248_ _04249_ _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_63_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06445_ _01913_ _01914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_29_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_15_0_wb_clk_i clknet_0_wb_clk_i clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09164_ _02561_ _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_90_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08115_ cpu.uart.receive_buff\[7\] _03370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06376_ _01348_ _01844_ _01845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05327_ cpu.PORTA_DDR\[3\] net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_44_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09095_ _02544_ _04143_ _04144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05658__I _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08046_ cpu.spi.data_out_buff\[3\] _03320_ _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05258_ _00737_ _00758_ _00759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_112_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09021__A1 _02701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05189_ _00002_ _00694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_101_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09997_ _02532_ _04939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08948_ _02776_ _04021_ _04026_ _00408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09324__A2 _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08879_ _03919_ _03971_ _03972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_88_Left_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05441__S0 _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09088__A1 _02755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05649__A1 _01119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06310__A2 _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08063__A2 _00676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09260__A1 _01105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_97_Left_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05821__A1 cpu.C vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10206_ _00079_ clknet_leaf_99_wb_clk_i cpu.regs\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_30_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10137_ _00014_ clknet_leaf_121_wb_clk_i cpu.regs\[9\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10068_ _02503_ _04999_ _05000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__05680__S0 _00917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06129__A2 _00730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09079__A1 _01830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08119__I net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06230_ _01700_ _01701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_5_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09251__A1 _01829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06161_ _01618_ _01534_ _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06092_ cpu.spi.busy _01235_ _01561_ _01563_ _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05112_ _00621_ _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_41_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09920_ net66 _04880_ _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09003__A1 _02891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05812__A1 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08789__I _03894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07693__I _01405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09851_ _04831_ _04821_ _04823_ _04832_ _04792_ _00505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09554__A2 _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06368__A2 _00976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09782_ _03551_ _04773_ _04774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08802_ _03906_ _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06994_ _02383_ _02439_ _02457_ _02458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05415__I1 cpu.regs\[1\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08733_ _03842_ _03856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_56_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05945_ _01411_ _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_95_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08664_ _03805_ _03808_ _03809_ _00341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05876_ _01104_ _01338_ _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08595_ _03748_ _01413_ _03749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07615_ _01117_ _01139_ _02987_ _02988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_76_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07546_ cpu.regs\[14\]\[1\] _02940_ _02942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07868__I _03164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07477_ cpu.uart.receive_div_counter\[1\] _02878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09216_ cpu.last_addr\[13\] _04198_ _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08293__A2 _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_107_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06428_ cpu.timer_top\[13\] _01465_ _01177_ _01897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09147_ _04182_ _00451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06359_ _01408_ _01827_ _01828_ _00017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09242__A1 _01639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09078_ _02745_ _04086_ _04129_ _04130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08029_ _03265_ _03303_ _03307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_73_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09545__A2 _04534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output55_I net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07271__C _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06295__A1 cpu.timer_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10686_ _00558_ clknet_leaf_64_wb_clk_i net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10091__A2 _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06598__A2 _01164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07547__A1 _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05730_ _00668_ _00658_ _00576_ _00583_ _01204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA_clkbuf_leaf_42_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05661_ _01134_ _01135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08380_ _02809_ _03585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_86_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07400_ _02813_ _02796_ _02814_ _02810_ _00072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07331_ _02670_ _02760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05592_ _01060_ _01064_ _01065_ _01066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_9_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07262_ _01915_ _02701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_45_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08027__A2 cpu.spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09001_ _04065_ _04066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09224__A1 _04238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06213_ _00613_ _01589_ _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07193_ _02135_ _02638_ _02643_ _02644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06144_ _01384_ _01595_ _01613_ _01615_ _01616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06075_ _01244_ _01547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09903_ _04871_ _04873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09834_ _04807_ _04818_ _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_81_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06210__A1 _00946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09765_ _00578_ _00579_ _04759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06977_ _02392_ _02441_ _02442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_29_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09696_ cpu.last_addr\[1\] cpu.last_addr\[0\] _04696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_69_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08716_ _03724_ _03846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05928_ _01337_ _01339_ _01365_ _01401_ _01402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_107_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08647_ cpu.toggle_ctr\[3\] _03793_ _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07091__C _02547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05859_ _01331_ _01332_ _01125_ _01333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_1_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08578_ cpu.toggle_ctr\[9\] _01410_ _01275_ cpu.toggle_ctr\[8\] _03732_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_37_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07529_ _02927_ _02928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10540_ _00413_ clknet_leaf_50_wb_clk_i cpu.timer_div\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09215__A1 _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10471_ _00344_ clknet_leaf_5_wb_clk_i cpu.toggle_ctr\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05315__I0 cpu.regs\[12\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10669_ _00541_ clknet_leaf_58_wb_clk_i cpu.PORTA_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06900_ _02310_ _02364_ _02365_ _02366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__06991__A2 _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07880_ _03173_ _00193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06831_ _00772_ _02297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07940__A1 cpu.timer_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07940__B2 cpu.timer_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09550_ _04555_ _04556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06762_ _02226_ _02227_ _02228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_05713_ _01186_ _01014_ _01187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08501_ _03676_ _03678_ _00309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_54_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09481_ _04485_ _04488_ _04489_ _04490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08432_ cpu.uart.receive_div_counter\[12\] _03617_ _03618_ _03626_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06693_ _00741_ _02008_ _02159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05644_ _01054_ _01118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08363_ _02919_ _03570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05575_ _01004_ _01047_ _01048_ _01049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_34_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08294_ _03519_ _03520_ _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07314_ cpu.timer\[5\] _02741_ _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_62_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06259__A1 _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07245_ cpu.uart.divisor\[2\] _02676_ _02686_ _02687_ _02688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_61_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07176_ _02614_ _02619_ _02627_ _02628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06127_ _01597_ _01598_ _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_112_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06431__A1 _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06058_ _01528_ _01529_ _01530_ _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_70_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07881__I _03164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08977__I _00962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09817_ _04761_ _04802_ _02516_ _04803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09748_ _04743_ _04740_ _04744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_69_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09684__A1 _04362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09679_ cpu.PC\[13\] _01340_ _04679_ _04680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__09601__I _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput19 io_in[2] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_107_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10523_ _00396_ clknet_leaf_9_wb_clk_i cpu.timer\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07121__I _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10454_ _00327_ clknet_leaf_16_wb_clk_i cpu.toggle_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10385_ _00258_ clknet_leaf_50_wb_clk_i cpu.uart.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_70_Left_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06422__A1 cpu.timer_div\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07922__A1 cpu.timer_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07922__B2 cpu.timer_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09675__A1 _03708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06489__B2 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06489__A1 _01132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09427__A1 _04413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05360_ _00006_ _00840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_31_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05291_ cpu.regs\[12\]\[6\] cpu.regs\[13\]\[6\] cpu.regs\[14\]\[6\] cpu.regs\[15\]\[6\]
+ _00788_ _00789_ _00790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07030_ _00574_ _02487_ _02492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05486__I _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08981_ cpu.timer_div\[4\] _04046_ _04048_ _04050_ _04051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_48_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07932_ cpu.timer_top\[11\] _03217_ _03210_ cpu.timer_top\[12\] _03221_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_07863_ _03116_ _03158_ _03159_ _03160_ _00189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_09602_ cpu.orig_PC\[10\] _04374_ _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07913__A1 _02046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05519__A3 _00642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06814_ _02279_ _02219_ _02280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_39_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09533_ cpu.PC\[6\] _01054_ _04515_ _04540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07794_ _01406_ _03100_ _03102_ _00178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_104_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09666__A1 _02414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06745_ _02208_ _02210_ _02211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_66_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09464_ _04454_ _04473_ _04474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06676_ _02136_ _02137_ _02138_ _02141_ _02142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_TAPCELL_ROW_19_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08415_ _03609_ _03612_ _00289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwire98 _00587_ net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_65_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09395_ _04293_ _04407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05627_ _00647_ _00987_ _01100_ _01101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08346_ _03559_ _00273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05558_ _01031_ _01032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08277_ cpu.uart.counter\[0\] _03507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05489_ cpu.regs\[8\]\[5\] cpu.regs\[9\]\[5\] cpu.regs\[10\]\[5\] cpu.regs\[11\]\[5\]
+ _00918_ _00891_ _00965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_34_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07228_ _02000_ _02672_ _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_61_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07159_ _02585_ _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10170_ _00047_ clknet_leaf_40_wb_clk_i cpu.uart.divisor\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_100_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05143__A1 cpu.uart.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10506_ _00379_ clknet_leaf_16_wb_clk_i cpu.timer_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07840__B1 _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10437_ _00310_ clknet_leaf_90_wb_clk_i cpu.orig_PC\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10368_ _00241_ clknet_leaf_32_wb_clk_i cpu.uart.div_counter\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10299_ _00172_ clknet_leaf_3_wb_clk_i cpu.regs\[4\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_108_Left_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_87_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06530_ cpu.toggle_top\[6\] _01417_ _01418_ _01997_ _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_87_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06461_ _01928_ _01929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_16_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08200_ _03391_ _03444_ _03446_ _03447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_44_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05412_ _00890_ _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_29_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_117_Left_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09180_ cpu.ROM_addr_buff\[2\] _04206_ _04209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09120__I0 _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06392_ _01511_ _01837_ _01860_ _01861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08131_ _03382_ cpu.uart.divisor\[5\] cpu.uart.divisor\[0\] _03383_ _03384_ _03385_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_71_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05343_ _00006_ _00823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08062_ _03163_ _03277_ _03332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_71_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05274_ _00751_ _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07013_ _02474_ _02475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_EDGE_ROW_96_Right_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_71_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08964_ _03420_ _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_110_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08139__A1 _02891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07915_ _03203_ _03204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05944__I _01416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08895_ _01046_ _01036_ _02673_ _03985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_07846_ _03143_ _03144_ _03145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_input17_I io_in[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09639__A1 _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07777_ cpu.regs\[4\]\[3\] _03087_ _03091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09516_ _04368_ _04510_ _04523_ _04400_ _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06728_ _02139_ _02193_ _02194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_93_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08311__A1 _02800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09447_ _04237_ _04448_ _04456_ _04457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06659_ _01287_ _02124_ _01337_ _01386_ _02125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__09111__I0 cpu.ROM_addr_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09378_ _04389_ _04390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08329_ cpu.uart.data_buff\[7\] _03527_ _03548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_76_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10222_ _00095_ clknet_leaf_117_wb_clk_i cpu.regs\[14\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10153_ _00030_ clknet_leaf_100_wb_clk_i cpu.br_rel_dest\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05600__A2 _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07274__C _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10084_ _04274_ _04278_ _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_97_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input9_I io_in[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05961_ _01077_ _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07700_ cpu.regs\[7\]\[0\] _03040_ _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_49_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08680_ _03743_ _03818_ _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05892_ _01344_ _01366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07631_ _02981_ _02991_ _02998_ _00119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08296__B _02793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07562_ _02600_ _02937_ _02951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06513_ _01979_ _01980_ _01981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_75_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09301_ _04314_ _04315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07493_ cpu.uart.receive_div_counter\[12\] _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_91_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09232_ _02761_ _04241_ _04249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_63_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06444_ _01907_ _01912_ _01913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_17_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09163_ _02496_ _02487_ _04194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06375_ _01842_ _01843_ _01844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08114_ _03368_ _03361_ _03369_ _00231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05326_ cpu.PORTB_DDR\[3\] net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__05939__I _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09094_ _04141_ _04143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08045_ _03313_ _03320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05257_ cpu.regs\[8\]\[4\] cpu.regs\[9\]\[4\] cpu.regs\[10\]\[4\] cpu.regs\[11\]\[4\]
+ _00752_ _00754_ _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_112_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05188_ _00687_ _00691_ _00692_ _00693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_101_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09996_ cpu.PORTA_DDR\[4\] _04937_ _04938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08780__A1 cpu.timer_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08947_ cpu.spi.divisor\[3\] _04022_ _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05594__A1 _01050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08878_ _03209_ _03970_ _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07335__A2 _02763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07829_ _03117_ _03129_ _00186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05441__S1 _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07099__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06846__A1 _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05649__A2 _00986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10205_ _00078_ clknet_leaf_104_wb_clk_i cpu.regs\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08771__A1 cpu.timer_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10136_ _00013_ clknet_leaf_120_wb_clk_i cpu.regs\[9\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10067_ _02479_ _04797_ _04796_ _04768_ _04757_ _04999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_89_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_32_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06160_ _01509_ _01630_ _01613_ _01632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_25_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05111_ _00620_ _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06091_ _01562_ _00012_ _01235_ _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09850_ cpu.ROM_spi_dat_out\[3\] _04790_ _04832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_71_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09781_ _04769_ _04771_ _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05576__A1 _01009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08801_ cpu.timer_capture\[1\] _03902_ _03905_ _02708_ _03906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06993_ _02435_ _02438_ _02457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05415__I2 cpu.regs\[2\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08732_ _02813_ _03844_ _03855_ _03853_ _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05944_ _01416_ _01417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08663_ cpu.toggle_ctr\[8\] _03806_ _03809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05875_ _01348_ _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_95_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08594_ cpu.toggle_ctr\[1\] _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07614_ _01102_ _02100_ _02987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_62_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07545_ _01407_ _02939_ _02941_ _00090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07476_ cpu.uart.receive_div_counter\[2\] _02877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06828__A1 _00710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06828__B2 _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09215_ _00667_ _04232_ _04233_ _00468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06427_ cpu.timer_top\[5\] _01459_ _01895_ _01264_ _01896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_9_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05669__I _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09146_ cpu.ROM_addr_buff\[9\] _04180_ _04181_ _04182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06358_ cpu.regs\[9\]\[4\] _01544_ _01828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09242__A2 _01731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06289_ cpu.timer_div\[4\] _01185_ _01758_ _01182_ _01759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09077_ cpu.orig_IO_addr_buff\[5\] _04090_ _04129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05309_ _00806_ _00807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08028_ _03261_ _03306_ _00208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_49_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_49_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_32_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09979_ _02790_ _04919_ _04926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07556__A2 _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08505__A1 _02859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07124__I _02557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_105_Right_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_84_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06184__B _01229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10685_ _00557_ clknet_leaf_96_wb_clk_i cpu.C vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08992__A1 _00586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10119_ _01406_ _05044_ _05046_ _00559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_117_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05660_ _01095_ _01133_ _00591_ _00637_ _01134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_58_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05591_ _01053_ _00630_ _01065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07330_ _02749_ _02759_ _00057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_85_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07261_ _02700_ _00047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09000_ _01017_ _03712_ _04065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_61_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06212_ _00903_ _01481_ _01682_ _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07192_ _02639_ _02640_ _02641_ _02642_ _02643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_26_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06143_ _01614_ _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08983__A1 _02698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06074_ cpu.timer_div\[2\] _01546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_6_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09902_ _04871_ _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09833_ cpu.ROM_spi_dat_out\[0\] _04812_ _04817_ _04818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08735__A1 _02791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07538__A2 _01108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09764_ _04753_ _02481_ _02474_ _04757_ _04758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_06976_ _02440_ _02441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_29_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09695_ _04690_ _04693_ _04694_ _04695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06269__B cpu.PORTA_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08715_ cpu.pwm_top\[0\] _03844_ _03845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05927_ _01368_ _01369_ _01377_ _01400_ _01401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_107_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05173__B _00679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08646_ cpu.toggle_ctr\[3\] _03793_ _03797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05858_ _00636_ _01332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_1_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05789_ _01261_ _01179_ _01262_ _01263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08577_ cpu.toggle_ctr\[11\] _03729_ _03730_ cpu.toggle_ctr\[10\] _03731_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_37_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07528_ _02874_ cpu.uart.receive_counter\[1\] _02875_ _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09463__A2 _04448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07459_ _02351_ _02356_ _02864_ _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10470_ _00343_ clknet_leaf_5_wb_clk_i cpu.toggle_ctr\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09129_ _04061_ _04169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_118_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08974__A1 cpu.timer_div\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07119__I _02574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05960__A1 cpu.PORTB_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10668_ _00540_ clknet_leaf_58_wb_clk_i cpu.PORTB_DDR\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07217__A1 _01830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10599_ _00471_ clknet_leaf_57_wb_clk_i cpu.IE vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08717__A1 _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06830_ _00763_ _00872_ _02295_ _02296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06761_ _02178_ _02182_ _02227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05712_ _01069_ _00605_ _01186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08500_ _02831_ _03674_ _03677_ _03678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_54_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09480_ _04304_ _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06692_ _02154_ _02157_ _02158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08431_ cpu.uart.receive_div_counter\[13\] _03625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05643_ _01116_ _01117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_92_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08362_ cpu.uart.receive_div_counter\[0\] _03569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05574_ _01019_ _01025_ _01006_ _01048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_58_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08293_ _01321_ _03264_ _03520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07313_ _02012_ _02745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_62_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07456__A1 _02859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07244_ _02546_ _02687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07175_ _02620_ _02623_ _02626_ _02627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_112_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10074__B net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08956__A1 _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06126_ _01339_ _01380_ _01496_ _01512_ _01598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__09863__B _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06057_ _01373_ _01518_ _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_70_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09816_ _04795_ _04796_ _04801_ _04802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05242__I0 cpu.regs\[0\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09747_ _02114_ _04743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06959_ _00773_ _02128_ _02424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09678_ _04677_ _04656_ _04678_ _04679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08629_ _03742_ _02053_ _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_81_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_64_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_64_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_64_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10522_ _00395_ clknet_leaf_9_wb_clk_i cpu.timer\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06018__I _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10453_ _00326_ clknet_leaf_12_wb_clk_i cpu.toggle_top\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06670__A2 _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08947__A1 cpu.spi.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10384_ _00257_ clknet_leaf_50_wb_clk_i cpu.uart.counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06422__A2 _01647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06186__A1 _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09124__A1 _02605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06110__A1 _00952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05290_ _00775_ _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07610__A1 _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08980_ _04049_ _04050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07931_ _03218_ _03219_ _03220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07862_ _00743_ _03116_ _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09601_ _04604_ _04605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06813_ _02240_ _02270_ _02268_ _02279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XTAP_TAPCELL_ROW_39_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09532_ cpu.PC\[6\] _01118_ _04539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07793_ cpu.regs\[3\]\[0\] _03101_ _03102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_104_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09666__A2 _04443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06744_ _02142_ _02169_ _02209_ _02210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_78_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09463_ _04455_ _04448_ _04472_ _04436_ _04473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06675_ _02139_ _02140_ _02141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_19_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06547__B _01970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08414_ _02882_ _03576_ _03610_ _03611_ _03612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_65_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09394_ _02855_ _04403_ _04405_ _04406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05626_ _01099_ _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08345_ cpu.uart.receive_buff\[1\] _03555_ _03557_ cpu.uart.receive_buff\[2\] _03559_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05557_ cpu.IO_addr_buff\[3\] cpu.IO_addr_buff\[2\] _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_80_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09418__A2 _04415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08276_ _03504_ _03506_ _00256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05488_ _00637_ _00962_ _00963_ _00964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_34_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07227_ _01147_ _01282_ _02672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_115_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07158_ _02610_ _00034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06109_ cpu.toggle_top\[10\] _01274_ _01578_ _01580_ _01581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__07892__I _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07089_ net12 _02543_ _02549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_clkbuf_4_4_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09354__A1 _02859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_111_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_111_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06168__A1 net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09106__A1 _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07668__A1 _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05143__A2 cpu.spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09409__A2 _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06340__A1 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06971__I _00807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10505_ _00378_ clknet_leaf_11_wb_clk_i cpu.timer_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07840__A1 _01541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10436_ _00309_ clknet_leaf_88_wb_clk_i cpu.orig_PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10367_ _00240_ clknet_leaf_28_wb_clk_i cpu.uart.div_counter\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08898__I _03985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10298_ _00171_ clknet_leaf_3_wb_clk_i cpu.regs\[4\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07307__I _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07659__A1 _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06460_ _01927_ _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05411_ _00833_ _00890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08130_ cpu.uart.div_counter\[4\] cpu.uart.divisor\[4\] _03384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_50_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06391_ _01773_ _01390_ _01836_ _01395_ _01335_ _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_16_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09120__I1 _02861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05342_ _00821_ _00822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08061_ net16 _03331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_113_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05273_ cpu.regs\[2\]\[5\] _00773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07831__A1 _03130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07012_ cpu.startup_cycle\[4\] _02474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08963_ _01414_ _00979_ _01180_ _04036_ _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_07914_ cpu.timer\[14\] _03203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_110_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08894_ _03984_ _00396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07845_ _02642_ _02370_ _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07776_ _03045_ _03086_ _03090_ _00172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_91_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09515_ _04373_ _04512_ _04522_ _04397_ _04523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06727_ _00806_ _00945_ _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_65_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09446_ cpu.orig_PC\[4\] _04272_ _04456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06658_ _00638_ _02124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_93_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05609_ _01079_ _01083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_81_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06589_ _01293_ _02055_ _02056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09377_ _01135_ _04389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08328_ cpu.uart.data_buff\[8\] _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08259_ cpu.uart.div_counter\[13\] _03493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07822__A1 _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06389__A1 _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10221_ _00094_ clknet_leaf_117_wb_clk_i cpu.regs\[14\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10152_ _00029_ clknet_leaf_94_wb_clk_i cpu.instr_buff\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09327__A1 _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10083_ _04278_ _04279_ _05013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06561__A1 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_22_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09263__B1 _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06616__A2 _01952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07813__A1 _02106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05110__I _00619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10419_ _00292_ clknet_leaf_34_wb_clk_i cpu.uart.receive_div_counter\[12\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_61_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05960_ cpu.PORTB_DDR\[1\] _01432_ _01203_ _01433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_49_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05891_ _01342_ _01360_ _01364_ _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_07630_ cpu.regs\[11\]\[5\] _02989_ _02998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07561_ _02098_ _02945_ _02950_ _00097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06512_ cpu.uart.divisor\[14\] _01440_ _00012_ _01980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09300_ _01398_ _01341_ _04314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07492_ cpu.uart.divisor\[12\] _02893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05107__A2 cpu.needs_timer_interrupt vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06304__A1 _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06304__B2 _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10100__A2 _01952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09231_ _02733_ _04247_ _04248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06443_ _01909_ _01911_ _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09162_ _03420_ _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06374_ _01832_ _01841_ _01843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08113_ cpu.uart.dout\[6\] _03351_ _03362_ _03369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05325_ cpu.PORTA_DDR\[2\] net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07804__A1 cpu.regs\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09093_ _04141_ _04142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08044_ _02773_ _03308_ _03318_ _03319_ _00211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05256_ _00682_ _00757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_31_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05187_ _00002_ _00692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__05955__I _01196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09995_ _04928_ _04937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09309__A1 _02831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09871__B _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08946_ _02773_ _04021_ _04025_ _00407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05433__I3 cpu.regs\[15\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08877_ _03960_ cpu.timer\[12\] _03961_ _03970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_99_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07828_ _03118_ _02105_ _03119_ _03128_ _03129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07759_ cpu.regs\[5\]\[4\] _03076_ _03080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_109_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07099__A2 _02543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_106_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09429_ _04439_ _04315_ _04324_ _04440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_54_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06059__B1 _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09548__A1 _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10204_ _00077_ clknet_leaf_103_wb_clk_i _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10135_ _02985_ _05050_ _05055_ _00566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10066_ _04946_ _04997_ _04955_ _04998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_89_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08523__A2 _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05110_ _00619_ _00620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_81_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06090_ cpu.uart.dout\[2\] _01562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_40_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08800_ _03259_ _03903_ _03904_ _03905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09780_ _04769_ _04771_ _04772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06992_ _02380_ _02455_ _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05415__I3 cpu.regs\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05943_ _01178_ _01415_ _01416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08731_ cpu.pwm_top\[6\] _03842_ _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08662_ cpu.toggle_ctr\[8\] _03806_ _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05874_ _01347_ _01348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07613_ _02985_ _02978_ _02986_ _00113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08593_ _03733_ _03741_ _03746_ _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_88_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07544_ cpu.regs\[14\]\[0\] _02940_ _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07475_ cpu.uart.divisor\[2\] _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_24_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09214_ cpu.ROM_addr_buff\[12\] _04213_ _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06426_ _01260_ _01893_ _01894_ _01895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_106_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06274__C _01225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09145_ _04060_ _04181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_71_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06357_ _01826_ _01827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06288_ _01756_ _01757_ _01758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09076_ _04122_ _04126_ _04128_ _00434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05308_ _00805_ _00806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08027_ _03305_ cpu.spi.busy _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05239_ _00740_ _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06439__S1 _00935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09950__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09978_ _04925_ _00539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_89_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_89_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08929_ _03203_ _04006_ _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_18_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_18_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07405__I _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10684_ _00556_ clknet_leaf_54_wb_clk_i net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_51_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10000__A1 _02698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09941__A1 _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10118_ cpu.regs\[15\]\[0\] _05045_ _05046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06507__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10049_ _02501_ _04961_ _04981_ _04982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_59_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_11_Left_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05590_ _00597_ _01064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07260_ cpu.uart.divisor\[5\] _02689_ _02699_ _02687_ _02700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_38_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06211_ _01680_ _01681_ _01152_ _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07191_ _02590_ _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06142_ _01382_ _01385_ _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06073_ _01143_ _01543_ _01545_ _00014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09901_ _01076_ _03712_ _04871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_41_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09832_ _04808_ _04813_ _04817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09763_ _04754_ _04756_ _04757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_clkbuf_4_9_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08714_ _03841_ _03844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06975_ _02432_ _02439_ _02440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_29_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09694_ _04691_ _04694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07225__I _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05926_ _01393_ _01399_ _01400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_107_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08645_ _03795_ _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05857_ _01095_ _01331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_1_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07171__A1 _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08576_ cpu.toggle_top\[10\] _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07527_ _02924_ _02925_ _02926_ _00087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09999__A1 cpu.PORTA_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05788_ _01048_ _01262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07458_ _02592_ _02357_ _02864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06409_ net3 _01221_ _01745_ _01878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07389_ cpu.toggle_top\[11\] _02802_ _02807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09128_ _00773_ _02622_ _04167_ _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_118_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09059_ cpu.orig_IO_addr_buff\[2\] _04106_ _04114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06985__A1 _02015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09923__A1 _02706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output60_I net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10667_ _00539_ clknet_leaf_58_wb_clk_i cpu.PORTB_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05476__A1 _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10598_ _00470_ clknet_leaf_55_wb_clk_i cpu.TIE vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05228__A1 _00722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput90 net90 sram_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06728__A1 _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06760_ _02220_ _02221_ _02225_ _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05711_ _01184_ _01185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06691_ _02155_ _02156_ _02157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08430_ _03503_ _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_77_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05642_ _01111_ _00986_ _01115_ _01116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__07153__A1 _02605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08361_ _03568_ _00279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_86_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05573_ _01045_ _01046_ _01047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08292_ _03408_ _03411_ _03519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07312_ _02727_ _02744_ _00054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_62_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07456__A2 _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07243_ _02685_ _02677_ _02686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06664__B1 _02128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07174_ _02625_ _02626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05449__B _00887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06125_ _01596_ _01597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_100_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06056_ _01354_ _01496_ _01529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09815_ _04798_ _04800_ _02503_ _04801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09435__I _04443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09746_ _04741_ _04742_ _04251_ _00490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05242__I1 _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06958_ _02422_ _02423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05909_ _01129_ _01382_ _01383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09677_ _04646_ _00879_ _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_96_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08628_ _03744_ _03781_ _03782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06889_ _02337_ _02338_ _02342_ _02355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__07144__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08892__A1 _03909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08559_ cpu.toggle_top\[2\] _03715_ _03719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10521_ _00394_ clknet_leaf_9_wb_clk_i cpu.timer\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05203__I _00003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10452_ _00325_ clknet_leaf_11_wb_clk_i cpu.toggle_top\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10383_ _00256_ clknet_leaf_39_wb_clk_i cpu.uart.has_byte vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_33_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_33_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_103_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07135__A1 _02315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05146__B1 cpu.needs_interrupt vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07438__A2 _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05449__A1 _00880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer1 _00898_ net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09060__A1 _02684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06949__A1 _02414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07930_ cpu.timer_top\[10\] _03207_ _03219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06879__I _00710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07861_ _01734_ _02423_ _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06812_ _02254_ _02255_ _02278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09600_ _03146_ _04578_ _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07792_ _03098_ _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_39_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09531_ _04498_ _04534_ _04537_ _04538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06743_ _02158_ _02168_ _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_104_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08874__A1 _03909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09462_ _04434_ _04457_ _04470_ _04471_ _04472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06674_ _00770_ _00944_ _02140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_19_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08413_ _03570_ _03611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_93_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09393_ _04404_ _04371_ _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05625_ _00989_ _01093_ _01098_ _00883_ _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08344_ _03558_ _00272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05556_ _01029_ _01030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_86_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06119__I _01120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09858__C _04792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08275_ _03353_ _03505_ _03506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05487_ _00947_ _00955_ _00963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07226_ _02670_ _02671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_1_0_wb_clk_i clknet_0_wb_clk_i clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_14_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07157_ _02588_ _02609_ _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06108_ _01277_ _01579_ _01580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_42_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07088_ _02548_ _00026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06039_ _00717_ _00873_ _01512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09354__A2 _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_12_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09729_ cpu.last_addr\[12\] cpu.ROM_addr_buff\[12\] _04728_ _04729_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__07668__A2 _03019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06628__B1 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10504_ _00377_ clknet_leaf_11_wb_clk_i cpu.timer_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10435_ _00308_ clknet_leaf_88_wb_clk_i cpu.orig_flags\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05603__A1 _00598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10366_ _00239_ clknet_leaf_49_wb_clk_i cpu.uart.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_51_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10297_ _00170_ clknet_leaf_13_wb_clk_i cpu.regs\[4\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09345__A2 _04336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08856__A1 cpu.timer_capture\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07659__A2 _03015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05410_ _00888_ _00825_ _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_16_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06390_ _01833_ _01808_ _01859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_90_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05341_ _00588_ _00821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08060_ _02791_ _03309_ _03330_ _00216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08154__I _03407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05272_ _00771_ _00772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_31_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07011_ _02472_ _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09584__A2 _04562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08962_ _00610_ _00586_ _02762_ _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_08893_ cpu.timer_capture\[15\] _03959_ _03983_ _03979_ _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07913_ _02046_ cpu.timer\[7\] _03199_ _03201_ _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_110_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07844_ _02265_ _02368_ _02369_ _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_EDGE_ROW_3_Left_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06570__A2 _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07775_ cpu.regs\[4\]\[2\] _03087_ _03090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09514_ _04518_ _04521_ _04522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06726_ _02170_ _02191_ _02192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09445_ _04361_ _04455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06657_ _01299_ _01064_ _01311_ _02123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_05608_ _01081_ _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_62_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06588_ _01284_ _01295_ _02055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09376_ _04350_ _04388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05539_ _00997_ _01013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08327_ _03546_ _00267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06086__A1 cpu.uart.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08258_ _03491_ _03492_ _00252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Left_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07209_ _02462_ _02614_ _02633_ _02658_ _02659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08189_ cpu.uart.counter\[3\] _03410_ _03436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_10220_ _00093_ clknet_leaf_121_wb_clk_i cpu.regs\[14\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10151_ _00028_ clknet_leaf_94_wb_clk_i cpu.instr_buff\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10082_ _01392_ _01280_ _05011_ _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07408__I _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_58_Left_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06561__A2 _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07143__I _02123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07510__A1 _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_67_Left_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09263__B2 _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09263__A1 _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07813__A2 _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09015__A1 _04047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10418_ _00291_ clknet_leaf_34_wb_clk_i cpu.uart.receive_div_counter\[11\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10349_ _00222_ clknet_leaf_47_wb_clk_i cpu.spi.data_in_buff\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07318__I _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_76_Left_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07329__A1 cpu.timer_capture\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05890_ _01357_ _01362_ _01363_ _01309_ _01364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_88_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07560_ cpu.regs\[14\]\[7\] _02946_ _02950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06511_ cpu.uart.divisor\[6\] _01230_ _01194_ _01978_ _01979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_75_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07491_ _02891_ _02892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05107__A3 _00616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09230_ _04240_ _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09689__B _04251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06442_ _00841_ _01910_ _00852_ _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_17_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09161_ _04192_ _00455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09254__A1 _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06373_ _01832_ _01841_ _01842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_16_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08112_ cpu.uart.receive_buff\[6\] _03368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05324_ cpu.PORTB_DDR\[2\] net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_09092_ _02535_ _03112_ _03113_ _02539_ _04141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_44_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08043_ cpu.spi.data_out_buff\[1\] _03301_ _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05255_ _00750_ _00755_ _00756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_112_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09557__A2 _04562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07568__A1 _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05186_ cpu.regs\[0\]\[0\] _00689_ _00690_ cpu.regs\[3\]\[0\] _00684_ _00686_ _00691_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_101_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09994_ _04928_ _04936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06240__A1 _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08945_ cpu.spi.divisor\[2\] _04022_ _04025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05594__A3 _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input22_I io_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08876_ _03969_ _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_98_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07827_ _02131_ _03121_ _03127_ _02105_ _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_07758_ _03047_ _03073_ _03079_ _00165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_67_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06709_ _02146_ _02171_ _02172_ _02174_ _02175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__07898__I cpu.timer_div\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07689_ _02983_ _03023_ _03031_ _00144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09428_ _04325_ _04439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_118_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09359_ _04370_ _04371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output90_I net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08522__I _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10203_ _00076_ clknet_leaf_103_wb_clk_i _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10134_ cpu.regs\[15\]\[7\] _05051_ _05055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10065_ _04194_ _04731_ _04734_ _04997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_89_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09720__A2 cpu.ROM_addr_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05417__S0 _00829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06198__B _01647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06534__A2 _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07495__B1 cpu.uart.receive_div_counter\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06298__A1 cpu.toggle_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10094__A2 _05019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09021__C _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09236__A1 _00672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07601__I _02967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09787__A2 _04777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07798__A1 cpu.regs\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_84_Left_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06222__A1 _01112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06991_ _02454_ _01165_ _02455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05942_ _01414_ _01008_ _01415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08730_ _02811_ _03844_ _03854_ _03853_ _00362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09711__A2 cpu.ROM_addr_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08661_ _03805_ _03806_ _03807_ _00340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05873_ _01346_ _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07612_ cpu.regs\[12\]\[7\] _02979_ _02986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_93_Left_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08592_ _03742_ _02053_ _03744_ _03745_ _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_76_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09475__A1 _02297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07543_ _02938_ _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07474_ cpu.uart.receiving _02875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06289__A1 cpu.timer_div\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09213_ cpu.last_addr\[12\] _04198_ _04232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06425_ cpu.timer_capture\[13\] _01256_ _01894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09144_ cpu.regs\[3\]\[1\] _03136_ _04167_ _04180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_16_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06356_ _01825_ _01826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06287_ cpu.spi.dout\[4\] _01566_ _01647_ _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09075_ cpu.IO_addr_buff\[4\] _04112_ _04127_ _04128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_71_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05307_ cpu.regs\[1\]\[7\] _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08026_ _02872_ _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05238_ cpu.regs\[1\]\[3\] _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05169_ _00663_ _00676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_73_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06213__A1 _00613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09977_ cpu.PORTB_DDR\[6\] _04918_ _04924_ _04916_ _04925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08928_ _04012_ _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_99_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08859_ _03858_ _03954_ _03955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_58_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_58_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_67_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10076__A2 _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10683_ _00555_ clknet_leaf_69_wb_clk_i net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09218__A1 _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06481__B _00641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_14_0_wb_clk_i clknet_0_wb_clk_i clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_10117_ _05043_ _05045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10048_ _02562_ _04743_ _04690_ _04978_ _04981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__06507__A2 _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07180__A2 _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05730__A3 _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06210_ _00946_ _01301_ _01681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10609__D _00481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07190_ net19 _02596_ _02641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06141_ _01597_ _01613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05786__I _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06072_ cpu.regs\[9\]\[1\] _01544_ _01545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09900_ _04870_ _00516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09831_ _04816_ _00501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10584__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09762_ _04755_ _04752_ _04756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07943__B2 cpu.timer_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07943__A1 cpu.timer_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06974_ _02435_ _02438_ _02439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08713_ _03842_ _03843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05925_ _01394_ _01396_ _01397_ _01353_ _01398_ _01399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09693_ _02489_ _02563_ _04693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_107_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08644_ _03789_ _03795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05856_ _01307_ _01315_ _01329_ _01330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05787_ _01250_ _01261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08575_ cpu.toggle_top\[11\] _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_1_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07526_ cpu.uart.receive_counter\[0\] cpu.uart.receive_counter\[1\] _02917_ _02926_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_77_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07241__I _01477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07457_ _02404_ _02862_ _02863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06408_ net64 _01078_ _01208_ _01876_ _01225_ _01877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_07388_ _02733_ _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_51_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09127_ _00669_ _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_60_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06339_ _01805_ _01807_ _01809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_105_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_105_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_118_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09058_ _04081_ _04110_ _04113_ _00431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_118_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08009_ cpu.spi.div_counter\[4\] _03291_ _03293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_9_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output53_I net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09631__I _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07151__I _02401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09787__B _02710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10666_ _00538_ clknet_leaf_58_wb_clk_i cpu.PORTB_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05476__A2 _00952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06990__I _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10597_ _00469_ clknet_leaf_74_wb_clk_i cpu.last_addr\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06425__A1 cpu.timer_capture\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05228__A2 _00730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08178__A1 _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput80 net80 io_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput91 net91 sram_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_37_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05710_ _01173_ _01028_ _01184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06690_ _02138_ _02141_ _02156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05641_ _01114_ _01115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08360_ _02931_ _03562_ _03567_ cpu.uart.receive_buff\[7\] _03568_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_86_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07311_ cpu.timer_capture\[4\] _02738_ _02743_ _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05572_ _01010_ _01046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_58_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_34_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_3_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_3_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_116_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08291_ _03412_ _03518_ _00259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_73_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07242_ _02684_ _02685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06664__B2 _02129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06664__A1 _01825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07173_ _02624_ _02425_ _02625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06124_ _01594_ _01595_ _01596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_41_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06055_ _01354_ _01507_ _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09814_ _02478_ _04799_ _04768_ _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07916__A1 cpu.timer_top\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07916__B2 cpu.timer_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09745_ _04692_ _04731_ _04742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09669__A1 _02398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05242__I2 _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06957_ _02104_ _02422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_05908_ _01126_ _00877_ _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06888_ _02352_ _02353_ _02354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09676_ _04646_ _00879_ _04677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_96_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08627_ _03735_ _03780_ _03781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05839_ _01136_ _01313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08558_ _02800_ _03714_ _03718_ _03717_ _00326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07509_ cpu.uart.receive_div_counter\[10\] _02910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__09841__A1 _04777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08489_ _01484_ _03651_ _03669_ _03653_ _00306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_92_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10520_ _00393_ clknet_leaf_9_wb_clk_i cpu.timer\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_30_Left_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_107_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10451_ _00324_ clknet_leaf_9_wb_clk_i cpu.toggle_clkdiv vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10382_ _00255_ clknet_leaf_31_wb_clk_i cpu.uart.div_counter\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_41_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_73_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_73_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08332__A1 _02790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09132__I0 cpu.regs\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_80_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05449__A2 _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10649_ _00521_ clknet_leaf_67_wb_clk_i net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xrebuffer2 _02280_ net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08938__A3 _03638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06949__A2 _02412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07860_ _03121_ _03156_ _03157_ _02422_ _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__07374__A2 _02674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06811_ _02272_ _02276_ _02277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07791_ _03099_ _03100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09530_ cpu.orig_PC\[7\] _04088_ _04537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06742_ _02194_ _02207_ _02208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_39_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09461_ _04340_ _04471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_104_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06673_ _00798_ _00950_ _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08412_ _02882_ _03607_ _03610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_80_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09392_ _04327_ _04404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05624_ _01097_ _01098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08343_ cpu.uart.receive_buff\[0\] _03555_ _03557_ cpu.uart.receive_buff\[1\] _03558_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05555_ _00994_ _01029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_80_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08274_ _01423_ cpu.uart.clr_hb _03505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06637__A1 _01116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07225_ _02669_ _02670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05486_ _00961_ _00962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_13_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07156_ _01825_ _02589_ _02599_ _02608_ _02586_ _02609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_115_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06107_ _01063_ _01066_ _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07087_ _00931_ _02541_ _02545_ _02547_ _02548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06038_ _01383_ _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_100_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08562__A1 _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07989_ _03272_ _03274_ _03275_ _03276_ _03277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_97_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09728_ cpu.last_addr\[11\] _04702_ _04728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08314__A1 _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_8_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09659_ _04389_ _04648_ _04660_ _04467_ _04661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10121__A1 _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05214__I _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_120_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_120_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_107_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06628__B2 _01638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10503_ _00376_ clknet_leaf_16_wb_clk_i cpu.timer_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10434_ _00307_ clknet_leaf_90_wb_clk_i cpu.orig_flags\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10365_ _00238_ clknet_leaf_65_wb_clk_i cpu.spi.counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09356__I _04361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10296_ _00169_ clknet_leaf_104_wb_clk_i cpu.regs\[5\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05340_ _00633_ _00820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_83_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05271_ _00770_ _00771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_113_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07010_ _00578_ _00579_ _02472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05794__I _01049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08961_ _04034_ _04035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08892_ _03909_ _03982_ _03901_ _03983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07912_ cpu.timer_top\[15\] _03200_ _03201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_110_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07843_ _00727_ _03116_ _03142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07774_ _03042_ _03086_ _03089_ _00171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07504__C1 _01427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09513_ _01924_ _04388_ _04520_ _04394_ _04521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06725_ _02186_ _02190_ _02191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10103__A1 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09444_ _04325_ _04454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06656_ _02107_ _02121_ _02122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05607_ _01038_ _01029_ _01080_ _01081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09375_ _04378_ _04382_ _04384_ _04386_ _04387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06587_ _02053_ _01273_ _01285_ _01279_ _02054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08326_ cpu.uart.data_buff\[6\] _03528_ _03545_ _03182_ _03546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05538_ _01011_ _01007_ _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XPHY_EDGE_ROW_104_Left_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06086__A2 _01230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08257_ _03488_ _03489_ _03464_ _03492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07283__A1 _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05469_ _00945_ _00946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08188_ _03432_ _03435_ _00238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07208_ _02603_ _02657_ _02658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_104_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07139_ _02123_ _02592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_83_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_76_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08783__A1 _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05597__A1 _01005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10150_ _00027_ clknet_leaf_94_wb_clk_i cpu.base_address\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10081_ _01359_ _01289_ _04265_ _05011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08535__A1 _03701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_113_Left_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_92_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09263__A2 _02855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09795__B _00666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07274__A1 _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10417_ _00290_ clknet_leaf_35_wb_clk_i cpu.uart.receive_div_counter\[10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07577__A2 _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10348_ _00221_ clknet_leaf_45_wb_clk_i cpu.spi.data_in_buff\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09019__C _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10279_ _00152_ clknet_leaf_105_wb_clk_i cpu.regs\[7\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_49_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05760__A1 _01186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06510_ _01975_ _01976_ _01977_ _01978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07490_ cpu.uart.divisor\[8\] _02891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06441_ cpu.regs\[0\]\[6\] cpu.regs\[1\]\[6\] cpu.regs\[2\]\[6\] cpu.regs\[3\]\[6\]
+ _01902_ _01153_ _01910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_29_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_100_Right_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_75_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09160_ cpu.ROM_addr_buff\[13\] _04191_ _04061_ _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06372_ net94 _01693_ _01789_ _01841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_29_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08111_ _03366_ _03361_ _03367_ _00230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09091_ _04122_ _04139_ _04140_ _00437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05323_ cpu.PORTA_DDR\[1\] net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06068__A2 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08042_ cpu.spi.data_out_buff\[2\] _03314_ _03318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05254_ cpu.regs\[12\]\[4\] cpu.regs\[13\]\[4\] cpu.regs\[14\]\[4\] cpu.regs\[15\]\[4\]
+ _00752_ _00754_ _00755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_24_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05185_ cpu.regs\[2\]\[0\] _00690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09993_ _02690_ _04929_ _04935_ _04932_ _00544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_08944_ _02769_ _04021_ _04024_ _00406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08517__A1 _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08875_ cpu.timer_capture\[12\] _03959_ _03968_ _03948_ _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07244__I _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07826_ _03120_ _03126_ _03127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input15_I io_in[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07740__A2 _03060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07757_ cpu.regs\[5\]\[3\] _03076_ _03079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06708_ _02144_ _02173_ _02174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_94_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07688_ cpu.regs\[8\]\[6\] _03021_ _03031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05699__I _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09427_ _04413_ _04437_ _04438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06639_ _02104_ _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09358_ _02846_ _04369_ _04370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_35_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08309_ cpu.uart.data_buff\[3\] _03533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06059__A2 _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09289_ _01309_ _00592_ _04302_ _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_105_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07419__I cpu.PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07559__A2 _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10202_ _00075_ clknet_4_2_0_wb_clk_i _00005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10133_ _02016_ _05050_ _05054_ _00565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08508__A1 _02861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10064_ _04977_ _04993_ _04996_ _02818_ _00554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_89_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05417__S1 _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05402__I _00880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06990_ _02436_ _02454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input7_I io_in[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05576__A4 _01049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05941_ _01002_ _01414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08660_ cpu.toggle_ctr\[7\] _03803_ _03807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05872_ _01345_ _01346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07611_ _02097_ _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_88_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08591_ cpu.toggle_ctr\[8\] _01275_ _03745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07542_ _02938_ _02939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07473_ cpu.uart.receive_counter\[0\] _02874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_62_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09212_ _00667_ _04230_ _04231_ _00467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06424_ cpu.timer_capture\[5\] _01569_ _01251_ _01892_ _01893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09143_ _04179_ _00450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06355_ _01485_ _01777_ _01824_ _01825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__08986__A1 _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05306_ _00804_ net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_06286_ cpu.spi.divisor\[4\] _01547_ _01189_ _01755_ _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09074_ _04102_ _04127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08025_ _03301_ _03302_ _03304_ _00207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05237_ _00737_ _00738_ _00707_ _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_31_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08738__A1 _00678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05168_ _00672_ cpu.needs_interrupt _00673_ _00674_ _00675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_TAPCELL_ROW_73_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05099_ _00577_ _00579_ _00580_ _00581_ _00609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_4
X_09976_ _02787_ _04919_ _04924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08927_ cpu.timer_capture\[13\] _04003_ _04011_ _03998_ _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08858_ cpu.timer\[9\] cpu.timer\[8\] _03938_ _03954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_98_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_4_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07809_ cpu.regs\[3\]\[7\] _03110_ _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08789_ _03894_ _03895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07702__I _01541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_98_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_98_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_94_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_27_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_27_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_23_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10682_ _00554_ clknet_leaf_68_wb_clk_i net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10116_ _05043_ _05044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10047_ _04690_ _04979_ _02564_ _04980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_89_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08901__A1 _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05730__A4 _00583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06140__A1 _01477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06140__B2 _01396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08968__A1 _04039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06140_ _01477_ _01391_ _01611_ _01396_ _01336_ _01612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_41_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06071_ _01141_ _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_111_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09830_ cpu.ROM_spi_dat_out\[0\] _04806_ _04815_ _04736_ _04816_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09761_ _02477_ _04755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06973_ _02434_ _02437_ _02438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08712_ _03841_ _03842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05924_ _01335_ _01398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09692_ _04691_ _04692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_107_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08643_ _03790_ _03793_ _03794_ _00335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05855_ _01316_ _01328_ _00987_ _01329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_95_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05786_ _01086_ _01260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08574_ _02815_ _03721_ _03728_ _03725_ _00332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_49_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07525_ _02875_ _02874_ _02922_ _02925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_76_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07456_ _02859_ _02838_ _02861_ _02862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06407_ _01212_ _01873_ _01874_ _01875_ _01876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_07387_ _02804_ _02801_ _02805_ _02697_ _00068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_17_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09126_ _04062_ _04165_ _04166_ _00446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_72_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06338_ _01781_ _01805_ _01807_ _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_17_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_31_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06269_ _01207_ _01217_ cpu.PORTA_DDR\[4\] _01739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09057_ _00567_ _04112_ _04103_ _04113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_60_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07631__A1 _02981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08008_ cpu.spi.div_counter\[4\] _03291_ _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_114_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09959_ cpu.PORTB_DDR\[1\] _04907_ _04911_ _04904_ _04912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07934__A2 cpu.timer\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output46_I net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_70_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10665_ _00537_ clknet_leaf_57_wb_clk_i cpu.PORTB_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_35_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10596_ _00468_ clknet_leaf_76_wb_clk_i cpu.last_addr\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput70 net70 io_out[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06189__A1 _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput81 net81 io_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput92 net92 sram_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09094__I _04141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_qcpu_99 io_oeb[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__07689__A1 _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05640_ _01113_ _01093_ _01097_ _00906_ _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05571_ _01020_ _01045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_4_13_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07310_ _02694_ _02739_ _02740_ _02742_ _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08290_ cpu.uart.counter\[2\] _03509_ _03517_ _03409_ _03518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07241_ _01477_ _02684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06664__A2 _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07861__A1 _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07172_ _01125_ _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_112_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07613__A1 _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06123_ _00731_ _00901_ _01595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_26_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06054_ _01350_ _01526_ _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_112_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_115_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09813_ _04770_ _04799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_6_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05927__A1 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09744_ _02111_ _04739_ _04740_ _04741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05242__I3 cpu.regs\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06956_ _02421_ _00021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09669__A2 _02412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09675_ _03708_ _04634_ _04425_ _04675_ _04676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06887_ _02321_ _00901_ _02349_ _02353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05907_ _01338_ _01380_ _01381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05838_ _01299_ _01088_ _01311_ _01312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08626_ _03779_ _03740_ _03780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_68_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06352__A1 _01337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05769_ _01186_ _01242_ _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_76_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08557_ _01413_ _03715_ _03718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07508_ cpu.uart.divisor\[10\] _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08488_ cpu.orig_flags\[1\] _03668_ _03669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_37_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07439_ _02403_ _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10450_ _00323_ clknet_leaf_48_wb_clk_i cpu.had_int vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09109_ _00690_ _02831_ _04153_ _04154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10381_ _00254_ clknet_leaf_29_wb_clk_i cpu.uart.div_counter\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07604__A1 _02977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05091__A1 _00598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09357__A1 _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05233__I3 cpu.regs\[15\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_42_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_42_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06487__B _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05146__A2 cpu.needs_timer_interrupt vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06343__B2 _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06343__A1 _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09798__B _03912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09132__I1 _02637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07843__A1 _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10648_ _00520_ clknet_leaf_66_wb_clk_i net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_3_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08938__A4 _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10579_ _00451_ clknet_leaf_85_wb_clk_i cpu.ROM_addr_buff\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_11_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08721__I _02685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09899__A2 _04869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09980__C _04098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06582__A1 cpu.timer_top\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06810_ _02273_ _02275_ _02276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07790_ _03098_ _03099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_39_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06741_ _02197_ _02206_ _02207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_64_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09460_ _04464_ _04469_ _04470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08411_ _03503_ _03609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_104_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06672_ _00805_ _00900_ _02138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09391_ _04329_ _04403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05623_ _01094_ _01096_ _01097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_19_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08342_ _03556_ _03557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05554_ _01001_ _01027_ _01028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08273_ _03503_ _03504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05485_ _00960_ _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06637__A2 _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08117__B _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07224_ _01392_ _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07155_ _02603_ _02607_ _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_115_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07086_ _02546_ _02547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06106_ _01575_ _01576_ _01577_ _01578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09339__A1 _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06037_ _01372_ _01373_ _01508_ _01509_ _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_100_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07247__I _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07988_ cpu.spi.div_counter\[3\] cpu.spi.divisor\[3\] _03276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06573__A1 cpu.timer_div\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_114_Right_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09727_ cpu.last_addr\[13\] _04723_ _04727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06939_ _02401_ _02404_ _02405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_96_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09658_ _02398_ _04426_ _04660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08609_ cpu.toggle_top\[7\] _03763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09589_ _04590_ _04592_ _04593_ _04347_ _04594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_65_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10502_ _00375_ clknet_leaf_16_wb_clk_i cpu.timer_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10433_ _00306_ clknet_leaf_90_wb_clk_i cpu.orig_flags\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10364_ _00237_ clknet_leaf_64_wb_clk_i cpu.spi.counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10295_ _00168_ clknet_leaf_105_wb_clk_i cpu.regs\[5\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05119__A2 _00627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05405__I _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08716__I _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07816__A1 _00690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05270_ cpu.regs\[1\]\[5\] _00770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_113_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08960_ _04033_ _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07911_ cpu.timer\[15\] _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08891_ cpu.timer\[15\] _03981_ _03982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_110_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07842_ _03141_ _00187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09512_ _04094_ _04509_ _04519_ _04392_ _04520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07773_ cpu.regs\[4\]\[1\] _03087_ _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_79_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06724_ _02188_ _02189_ _02190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06655_ _02109_ _02120_ _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_66_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09443_ _04407_ _04453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05606_ _01079_ _01080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09374_ _04385_ _04386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08325_ _02783_ _03540_ _03544_ _03545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06586_ cpu.toggle_top\[15\] _02053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05537_ cpu.IO_addr_buff\[1\] _01010_ _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__07807__A1 _02016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08256_ _03488_ _03453_ _03490_ _03470_ _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_61_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05468_ _00944_ _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_34_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08187_ _03416_ _03278_ _03434_ _03435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_6_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05294__A1 _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07207_ _02650_ _02652_ _02656_ _02630_ _02657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_05399_ _00877_ _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07138_ _02590_ _02591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_76_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05597__A2 _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07069_ _00619_ _02531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10080_ _01290_ _01166_ _05010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09732__B2 _04731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08536__I _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05285__A1 _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10416_ _00289_ clknet_leaf_34_wb_clk_i cpu.uart.receive_div_counter\[9\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10347_ _00220_ clknet_leaf_46_wb_clk_i cpu.spi.data_in_buff\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09971__A1 cpu.PORTB_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06005__B _01477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10278_ _00151_ clknet_leaf_106_wb_clk_i cpu.regs\[7\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06537__A1 _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05760__A2 _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10097__A1 _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06440_ _00824_ _01908_ _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_29_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07350__I _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06371_ _01838_ _01839_ _01840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_29_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08110_ cpu.uart.dout\[5\] _03358_ _03362_ _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05322_ cpu.PORTB_DDR\[1\] net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_09090_ cpu.IO_addr_buff\[7\] _03446_ _04127_ _04140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08041_ _02769_ _03309_ _03316_ _03317_ _00210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05253_ _00753_ _00754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05184_ _00688_ _00689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09992_ cpu.PORTA_DDR\[3\] _04930_ _04935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_110_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08943_ cpu.spi.divisor\[1\] _04022_ _04024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08874_ _03909_ _03967_ _03901_ _03968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07825_ _02642_ _03123_ _03124_ _03125_ _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_07756_ _03045_ _03073_ _03078_ _00164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_67_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10088__A1 _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06707_ cpu.regs\[1\]\[0\] _02007_ _02173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09426_ _04362_ _04415_ _04435_ _04436_ _04437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06585__B _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07687_ _02981_ _03023_ _03030_ _00143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06638_ _02101_ _02103_ _02104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06569_ cpu.uart.dout\[7\] _01560_ _01664_ _02036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09357_ _02838_ _02830_ _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08308_ _02671_ _03522_ _03526_ _03530_ _03532_ _00262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_62_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09288_ cpu.Z _00592_ _04302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08239_ _03448_ _03474_ _03477_ _03478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_62_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10126__I _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05409__I3 cpu.regs\[15\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10201_ _00074_ clknet_leaf_107_wb_clk_i _00004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output76_I net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10132_ cpu.regs\[15\]\[6\] _05051_ _05054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_100_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10063_ _04993_ _04994_ _04995_ _04996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__06519__A1 cpu.timer_div\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05664__B _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07192__A1 _02639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08266__I _03407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05940_ cpu.toggle_top\[1\] _01413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10508__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05871_ _01343_ _01344_ _01345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08590_ _03742_ cpu.toggle_top\[15\] cpu.toggle_top\[14\] _03743_ _03744_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07610_ _02983_ _02978_ _02984_ _00112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_109_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07541_ _02935_ _02937_ _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_118_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07486__A2 cpu.uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07080__I _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07472_ _02578_ _02870_ _02668_ _02873_ _00085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_8_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09211_ _02521_ _04220_ _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06423_ _01890_ _01891_ _01419_ _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08435__A1 _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09142_ cpu.ROM_addr_buff\[8\] _04178_ _04169_ _04179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06354_ _01780_ _01823_ _01824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05305_ _00803_ _00804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06285_ _01753_ _01754_ _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_21_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09073_ _01779_ _04123_ _04125_ _04109_ _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06997__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_114_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08024_ cpu.spi.data_out_buff\[7\] _03164_ _03303_ _03304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_102_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05236_ cpu.regs\[8\]\[3\] cpu.regs\[9\]\[3\] cpu.regs\[10\]\[3\] cpu.regs\[11\]\[3\]
+ _00711_ _00734_ _00738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_25_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05167_ _00584_ net18 _00674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_40_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05098_ _00573_ _00575_ _00608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_09975_ _04923_ _00538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08926_ _02745_ _04004_ _04005_ _04010_ _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08857_ _03896_ _03952_ _03953_ _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06299__C _01277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07808_ _03099_ _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08788_ _01414_ _01262_ _02763_ _03894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__09470__I _04446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07739_ cpu.regs\[6\]\[5\] _03058_ _03067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_109_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_60_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10681_ _00553_ clknet_leaf_68_wb_clk_i net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05488__A1 _00637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09409_ _02402_ _01806_ _04419_ _04420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_23_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_67_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_67_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_90_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05263__I1 _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10115_ _02937_ _02987_ _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_10046_ _04743_ _04978_ _02562_ _04979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_59_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06070_ _01542_ _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09917__A1 _04047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_105_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09760_ _02504_ _02505_ _04754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06972_ _02436_ _01929_ _02437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09691_ _02538_ _04058_ _02537_ _04691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08711_ _01175_ _02674_ _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05923_ _00822_ _01366_ _01397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_83_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08642_ cpu.toggle_ctr\[2\] _03791_ _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07156__A1 _01825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05854_ _01317_ _01318_ _01327_ _01328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_89_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05785_ cpu.timer_capture\[8\] _01256_ _01258_ _01259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08573_ cpu.toggle_top\[7\] _03722_ _03728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07524_ cpu.uart.receive_counter\[1\] _02924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_88_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07455_ _02860_ _02861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05323__I cpu.PORTA_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06406_ cpu.PORTB_DDR\[5\] _01039_ _01741_ _01875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_17_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07386_ cpu.toggle_top\[10\] _02802_ _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08959__A2 _02674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09125_ cpu.ROM_addr_buff\[4\] _04062_ _04166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06337_ _01806_ net93 _01807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_118_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09056_ _04111_ _04112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06268_ cpu.toggle_top\[12\] _01738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_08007_ _03287_ _03290_ _03291_ _00202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_102_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09908__A1 _04039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05493__I1 cpu.regs\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05219_ _00699_ _00719_ _00721_ _00707_ _00722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__05642__A1 _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06199_ cpu.timer_div\[3\] _01185_ _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09958_ _02768_ _04908_ _04911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09136__A2 cpu.regs\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08909_ _02728_ _03987_ _03988_ _03996_ _03997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09889_ cpu.pwm_top\[7\] cpu.pwm_counter\[7\] _04861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_114_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_114_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07147__A1 _01101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output39_I net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08972__C _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06122__A2 _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10664_ _00536_ clknet_leaf_57_wb_clk_i cpu.PORTB_DDR\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08544__I _03662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10595_ _00467_ clknet_leaf_73_wb_clk_i cpu.last_addr\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09072__A1 _02694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06999__I _02097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput60 net60 io_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07386__A1 cpu.toggle_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput71 net71 io_out[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput82 net82 io_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_101_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput93 net93 sram_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08583__B1 _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05936__A2 _01407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10029_ _04958_ _04963_ _04956_ _04964_ _04965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__05244__S0 _00733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05570_ _01004_ _01043_ _01027_ _01044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_46_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07310__A1 _02694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07240_ _02679_ _02676_ _02680_ _02683_ _00043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_54_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07171_ _02622_ _02405_ _02623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06122_ _00731_ _00901_ _01594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06053_ _01499_ _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07377__A1 _01275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09812_ _02477_ _04797_ _04798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_6_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09743_ _02580_ _02582_ _04691_ _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06955_ _02130_ _02420_ _02421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07533__I net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09674_ _04634_ _04671_ _04675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05906_ _01378_ _01379_ _01380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_06886_ _02336_ _02346_ _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_96_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05837_ _01144_ _00630_ _01311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08625_ _03731_ _03737_ _03736_ _03733_ _03779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_68_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08556_ _02671_ _03714_ _03716_ _03717_ _00325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07507_ _02902_ cpu.uart.divisor\[7\] _02903_ cpu.uart.receive_div_counter\[6\] _02907_
+ _02908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_81_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05768_ _00567_ _01046_ _01242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_49_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05699_ _01172_ _01173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08487_ _03640_ _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_80_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07852__A2 _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07438_ _01593_ _01641_ _02589_ _02845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07369_ _02790_ _02791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09054__A1 _00989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09108_ _00669_ _04153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10380_ _00253_ clknet_leaf_31_wb_clk_i cpu.uart.div_counter\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09039_ _04095_ _04096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06591__A2 _02021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_82_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_82_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_56_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_11_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_11_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_31_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10647_ _00519_ clknet_leaf_65_wb_clk_i net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_101_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09045__A1 _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10578_ _00450_ clknet_leaf_78_wb_clk_i cpu.ROM_addr_buff\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09348__A2 _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07618__I _02988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05209__I1 _00710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06740_ _02193_ _02205_ _02206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07353__I _00962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06671_ cpu.regs\[1\]\[5\] _00949_ _02137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08410_ _03606_ _03602_ _03608_ _03585_ _00288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05622_ _01095_ _00636_ _01051_ _01096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_09390_ _02555_ _04402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_19_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08341_ _02917_ _03348_ _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05553_ _01024_ _01026_ _01027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_59_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09284__A1 _00983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08272_ _00620_ _03503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08184__I _02793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06098__A1 _01546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05484_ _00958_ _00959_ _00960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06637__A3 _02102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07223_ _02578_ _02663_ _02668_ _02666_ _00041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_27_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07154_ _02135_ _02405_ _02606_ _02607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_115_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05757__B _01230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07085_ _00665_ _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_06105_ cpu.toggle_top\[2\] _01416_ _01418_ _01577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_42_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06270__A1 net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06036_ _01355_ _01371_ _01507_ _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_07987_ cpu.spi.div_counter\[1\] cpu.spi.divisor\[1\] _03275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__05456__S0 _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09726_ _04228_ cpu.ROM_addr_buff\[10\] _04701_ _04726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06938_ _02402_ _02403_ cpu.PC\[1\] _02404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__05492__B _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09899__B _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09657_ _04458_ _04657_ _04658_ _04296_ _04659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06869_ _02334_ _02335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_96_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08608_ _03755_ _03758_ _03761_ _03762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_09588_ _04489_ _04579_ _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08539_ cpu.orig_PC\[12\] _03643_ _03705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_38_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07212__B _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10501_ _00374_ clknet_leaf_16_wb_clk_i cpu.timer_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08822__I _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10432_ _00305_ clknet_leaf_90_wb_clk_i cpu.orig_flags\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10363_ _00236_ clknet_leaf_64_wb_clk_i cpu.spi.counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10294_ _00167_ clknet_leaf_105_wb_clk_i cpu.regs\[5\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08069__A2 _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10033__C1 cpu.ROM_addr_buff\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08792__A3 _03897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08890_ _03203_ _03197_ _03975_ _03981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07910_ cpu.timer_top\[9\] _03198_ _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07841_ _03131_ _03140_ _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07772_ _03034_ _03086_ _03088_ _00170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09511_ _02636_ _04390_ _04519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06723_ _02184_ _02185_ _02189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06654_ _02111_ _02113_ _02116_ _02119_ _02120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_78_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_65_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09442_ _02315_ _04449_ _04451_ _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05605_ _01011_ _01031_ _01079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06585_ cpu.toggle_top\[7\] _01416_ _01411_ _02051_ _02052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_09373_ _04296_ _04385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08324_ cpu.uart.data_buff\[7\] _03539_ _03544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05536_ cpu.IO_addr_buff\[0\] _01010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_46_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05331__I cpu.PORTA_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09009__A1 _03849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08255_ cpu.uart.div_counter\[12\] _03489_ _03490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05467_ _00943_ _00944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08186_ cpu.spi.counter\[4\] _03433_ _03434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_15_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05398_ cpu.base_address\[2\] _00877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07206_ _02654_ _02655_ _02656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07137_ _01150_ _02133_ _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07258__I _02012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_18_Left_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07068_ _00609_ _02526_ _02529_ _02518_ _02530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_2_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07991__B2 _03167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06019_ _01491_ net91 _01492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09709_ cpu.last_addr\[5\] cpu.ROM_addr_buff\[5\] _04698_ _04709_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__09496__B2 _04453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_27_Left_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_87_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09248__A1 _01638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07721__I _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05241__I cpu.regs\[2\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08471__A2 _03655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08552__I _03713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10415_ _00288_ clknet_leaf_35_wb_clk_i cpu.uart.receive_div_counter\[8\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_36_Left_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10346_ _00219_ clknet_leaf_45_wb_clk_i cpu.spi.data_in_buff\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06785__A2 _00855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07431__B1 _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10277_ _00150_ clknet_leaf_14_wb_clk_i cpu.regs\[7\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_49_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_45_Left_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09487__A1 _01829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_0_0_wb_clk_i clknet_0_wb_clk_i clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08727__I _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06370_ _01782_ _01787_ _01784_ _01839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05321_ _00818_ net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08040_ cpu.spi.data_out_buff\[0\] _03301_ _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_11_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_54_Left_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06473__A1 _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05252_ _00712_ _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05183_ cpu.regs\[1\]\[0\] _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09991_ _03849_ _04929_ _04934_ _04932_ _00543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_86_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07973__A1 _00663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08942_ _02760_ _04021_ _04023_ _00405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05984__B1 _01456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08873_ cpu.timer\[12\] _03966_ _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_63_Left_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07824_ _02310_ _02364_ _02365_ _03125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07755_ cpu.regs\[5\]\[2\] _03076_ _03078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07686_ cpu.regs\[8\]\[5\] _03021_ _03030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06706_ _00724_ _00973_ _02172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_50_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09425_ _04399_ _04436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06637_ _01116_ _01123_ _02102_ _02103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_118_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06568_ _02030_ _02032_ _02034_ _02035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_81_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05061__I net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09356_ _04361_ _04368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06157__I _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08307_ cpu.uart.data_buff\[1\] _03531_ _03532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_72_Left_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05519_ _00631_ _00991_ _00642_ _00992_ _00993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_06499_ _01629_ _01962_ _01963_ _01966_ _01967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_35_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09287_ _01316_ _04297_ _04300_ _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08238_ cpu.uart.div_counter\[8\] _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08169_ _00665_ _03420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10200_ _00011_ clknet_leaf_87_wb_clk_i cpu.instr_cycle\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10131_ _01921_ _05050_ _05053_ _00564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10062_ _02515_ _04812_ _00627_ _04980_ _04995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_101_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08141__B2 _03391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07451__I _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06455__A1 _01408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06207__A1 cpu.toggle_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10329_ _00202_ clknet_leaf_62_wb_clk_i cpu.spi.div_counter\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08231__B _03464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05870_ _00905_ _00640_ _01344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_109_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07540_ _01117_ _01124_ _02936_ _02937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_76_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09880__A1 _02533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07471_ _02576_ _02870_ _02667_ _02873_ _00084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_118_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09210_ cpu.last_addr\[11\] _04198_ _04230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06422_ cpu.timer_div\[5\] _01647_ _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_57_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09141_ _03696_ _04063_ _04177_ _04178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06353_ net30 _01096_ _01822_ _01094_ _01823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_71_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09072_ _02694_ _04105_ _04124_ _04125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05304_ _00791_ _00793_ _00797_ _00802_ _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_08023_ _03299_ _03277_ _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06284_ cpu.uart.dout\[4\] _01560_ _01665_ _01754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05235_ _00699_ _00737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05166_ _00614_ cpu.needs_timer_interrupt _00673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08920__I _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05097_ _00607_ _00012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09974_ cpu.PORTB_DDR\[5\] _04918_ _04922_ _04916_ _04923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08925_ cpu.timer\[13\] _04006_ _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input20_I io_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08856_ cpu.timer_capture\[9\] _03899_ _03912_ _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07807_ _02016_ _03101_ _03109_ _00184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08787_ _02717_ _03891_ _03892_ _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05999_ _01413_ _01417_ _01418_ _01471_ _01472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_79_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07738_ _03049_ _03060_ _03066_ _00158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_94_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07669_ _02017_ _03019_ _00136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10680_ _00552_ clknet_leaf_69_wb_clk_i net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05488__A2 _00962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09408_ cpu.PC\[2\] cpu.br_rel_dest\[2\] _04418_ _04419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_51_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09339_ _04298_ _04330_ _04352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_109_Right_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08830__I _03894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07937__A1 _02046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10114_ _05042_ _00558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_36_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_36_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05263__I2 cpu.regs\[2\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10045_ _02110_ _02519_ _02117_ _04978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_59_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07114__C _02533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06428__A1 cpu.timer_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09090__A2 _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05100__A1 _00608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06971_ _00807_ _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09690_ _02118_ _04690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08710_ _02670_ _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05922_ _01395_ _01396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05853_ _01186_ _01325_ _01203_ _01326_ _01327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_08641_ cpu.toggle_ctr\[2\] _03791_ _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_107_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05784_ _01257_ _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08572_ _02813_ _03721_ _03727_ _03725_ _00331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07523_ _02874_ _02917_ _02923_ _00086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07454_ _02402_ _02860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06667__A1 _00593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06405_ net56 _01172_ _01213_ _01084_ _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_64_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07385_ _02728_ _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09124_ _02605_ _00670_ _04164_ _04165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_60_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05890__A2 _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06336_ _01113_ _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_114_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09055_ _00677_ _04111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06267_ _01143_ _01736_ _01737_ _00016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08006_ cpu.spi.div_counter\[3\] _03289_ _03291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_114_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05493__I2 cpu.regs\[2\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05218_ _00002_ _00720_ _00721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05642__A2 _00986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06198_ cpu.spi.dout\[3\] _01450_ _01647_ _01668_ _01669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_05149_ cpu.instr_cycle\[3\] cpu.instr_cycle\[1\] _00652_ _00657_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_40_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09957_ _04910_ _00533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08908_ cpu.timer\[10\] _03989_ _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09888_ cpu.pwm_top\[6\] cpu.pwm_counter\[6\] _04860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_99_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08839_ cpu.timer\[7\] _03932_ _03938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_56_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09144__I0 cpu.regs\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10663_ _00535_ clknet_leaf_56_wb_clk_i cpu.PORTB_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_97_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10594_ _00466_ clknet_leaf_79_wb_clk_i cpu.last_addr\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07083__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06830__A1 _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput61 net61 io_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput50 net50 io_oeb[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_31_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput72 net72 io_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_101_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput94 net94 sram_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput83 net83 sram_addr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10028_ _04769_ _02483_ _04964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_106_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05424__I _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05244__S1 _00734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07170_ _02621_ _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06121_ _01588_ _01590_ _01592_ _01593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08470__I _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06052_ _01524_ _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_112_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07086__I _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09811_ _02504_ cpu.startup_cycle\[2\] _04797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08574__A1 _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09742_ _03305_ _04738_ _04739_ _00489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_10_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08326__B2 _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06954_ _02131_ _02132_ _02397_ _02418_ _02419_ _02420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09673_ _04557_ _04672_ _04673_ _04674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10133__A1 _02016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05905_ _00850_ _00854_ _01379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06885_ _02348_ _02350_ _02351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08624_ _03766_ _03777_ _03778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05836_ _01309_ _01310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05767_ cpu.spi.divisor\[0\] _01241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_68_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08555_ _03645_ _03717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07506_ _02883_ cpu.uart.receive_div_counter\[9\] cpu.uart.receive_div_counter\[3\]
+ _01658_ _02876_ cpu.uart.receive_div_counter\[2\] _02907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_TAPCELL_ROW_81_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08629__A2 _02053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05698_ _01171_ _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_76_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08486_ _01310_ _03651_ _03667_ _03653_ _00305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_49_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_13_0_wb_clk_i clknet_0_wb_clk_i clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_64_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07437_ _02844_ _00079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07852__A3 _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07368_ _02705_ _02790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06165__I _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06319_ _01694_ _01697_ _01789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09107_ _04152_ _00441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_103_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07299_ _00925_ _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_60_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08380__I _02809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09038_ _01800_ _04094_ _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_32_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_92_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08565__A1 cpu.toggle_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06114__B _01585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08317__A1 _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10124__A1 cpu.regs\[15\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09117__I0 _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08555__I _03645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06500__B1 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05303__A1 _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10646_ _00518_ clknet_leaf_66_wb_clk_i net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_101_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_51_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_51_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10577_ _00449_ clknet_leaf_81_wb_clk_i cpu.ROM_addr_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08556__A1 _02671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05209__I2 cpu.regs\[2\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08308__A1 _02671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06670_ _00799_ _00945_ _02136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05154__I net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05621_ _00590_ _01095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_86_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08340_ _03554_ _03555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05552_ _00995_ _01025_ _01026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08465__I _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08271_ cpu.uart.div_counter\[15\] _03498_ _03502_ _03479_ _00255_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_86_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05483_ _00939_ _00941_ _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07222_ _01111_ _02661_ _02668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_116_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07153_ _02605_ _02404_ _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06104_ cpu.pwm_top\[2\] _01269_ _01168_ _01576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07084_ _02542_ _02544_ _02545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06270__A2 _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06035_ _01355_ _01371_ _01507_ _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__08547__A1 _03432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05329__I cpu.PORTA_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07986_ cpu.spi.div_counter\[2\] _03269_ cpu.spi.div_counter\[4\] _03270_ _03273_
+ _03274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__05456__S1 _00910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09725_ cpu.ROM_addr_buff\[13\] _04724_ _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06937_ cpu.PC\[2\] _02403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09656_ _04489_ _04648_ _04658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08607_ _03759_ cpu.toggle_top\[3\] cpu.toggle_top\[2\] _03760_ _03761_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06868_ _02293_ _02323_ _02320_ _02334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__05533__A1 _01005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05819_ _00984_ _01288_ _01290_ _01293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09587_ _04343_ _04591_ _04592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06799_ _02239_ _02264_ _02265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08538_ _03703_ _03693_ _03704_ _03695_ _00320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_108_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08469_ _03639_ _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10500_ _00373_ clknet_leaf_16_wb_clk_i cpu.timer_top\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10431_ _00304_ clknet_leaf_101_wb_clk_i cpu.orig_IO_addr_buff\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10362_ _00235_ clknet_leaf_64_wb_clk_i cpu.spi.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06261__A2 _01731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10293_ _00166_ clknet_leaf_14_wb_clk_i cpu.regs\[5\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08538__A1 _03703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09266__A2 _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05383__S0 _00830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10629_ _00501_ clknet_leaf_73_wb_clk_i cpu.ROM_spi_dat_out\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08777__A1 _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07840_ _01541_ _02422_ _03132_ _03139_ _03115_ _03140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07364__I _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07771_ cpu.regs\[4\]\[0\] _03087_ _03088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09510_ _04378_ _04516_ _04517_ _04385_ _04518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06722_ _02140_ _02187_ _02181_ _02179_ _02188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_40_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06653_ _02117_ _02118_ _02119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_91_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09441_ _04450_ _04448_ _04451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05604_ _01077_ _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_65_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06584_ _02048_ _02049_ _02050_ _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09372_ _04383_ _04370_ _04384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08323_ _03543_ _00266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05535_ _01002_ _01004_ _01008_ _01009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_59_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08254_ _03399_ _03485_ _03489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05466_ _00942_ _00943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08185_ _03161_ _03425_ _03278_ _03428_ _03433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_05397_ _00876_ net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07205_ _02636_ _02620_ _02655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08768__A1 _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07136_ _02585_ _02589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07539__I _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07067_ _02506_ _02527_ _02483_ _02528_ _02529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_76_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06018_ _00981_ _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09708_ _04222_ cpu.ROM_addr_buff\[7\] _04699_ _04708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_07969_ _00613_ _03197_ _03257_ _03258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_69_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_87_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09639_ _02556_ _04627_ _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07259__A1 _02698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09248__A2 _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_41_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10414_ _00287_ clknet_leaf_35_wb_clk_i cpu.uart.receive_div_counter\[7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07431__A1 _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10345_ _00218_ clknet_leaf_46_wb_clk_i cpu.spi.data_in_buff\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05293__I0 cpu.regs\[8\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07431__B2 _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10276_ _00149_ clknet_leaf_2_wb_clk_i cpu.regs\[7\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_49_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07133__B _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05320_ _00817_ _00818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_29_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05251_ _00751_ _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07670__A1 _02098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07359__I _02012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05182_ cpu.regs\[4\]\[0\] cpu.regs\[5\]\[0\] cpu.regs\[6\]\[0\] cpu.regs\[7\]\[0\]
+ _00684_ _00686_ _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09990_ cpu.PORTA_DDR\[2\] _04930_ _04934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08941_ cpu.spi.divisor\[0\] _04022_ _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08872_ _03960_ _03907_ _03961_ _03966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08922__A1 _02694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07823_ _02642_ _02366_ _03124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08918__I _01456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09478__A2 cpu.br_rel_dest\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07754_ _03042_ _03073_ _03077_ _00163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07685_ _02977_ _03023_ _03029_ _00142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06705_ _00688_ _01928_ _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09424_ _04341_ _04431_ _04433_ _04434_ _04435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_35_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06636_ _01125_ _01131_ _01135_ _01926_ _02102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_59_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05342__I _00821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06567_ _02033_ _01193_ _00607_ _02034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09355_ _04326_ _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08306_ _03527_ _03531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08989__A1 _02706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05518_ cpu.br_rel_dest\[5\] cpu.br_rel_dest\[4\] _00992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06498_ _01959_ _01964_ _01965_ _01966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09286_ _04297_ _04299_ _04300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08237_ _03390_ _03473_ _03476_ _03450_ _00247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_90_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05449_ _00880_ _00902_ _00887_ _00927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08168_ _02794_ _03419_ _00234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_108_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_108_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08099_ cpu.uart.dout\[2\] _03358_ _00679_ _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07413__A1 _02106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07119_ _02574_ _02575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10130_ cpu.regs\[15\]\[5\] _05051_ _05053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10061_ _02527_ _04988_ _04994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09166__A1 _00609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07716__A2 _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08563__I _03713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06455__A2 _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06083__I _01196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08601__B1 cpu.toggle_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06207__A2 _01416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10328_ _00201_ clknet_leaf_63_wb_clk_i cpu.spi.div_counter\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05966__A1 net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_0_Left_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10259_ _00132_ clknet_leaf_0_wb_clk_i cpu.regs\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06391__A1 _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06391__B2 _01395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07470_ _02872_ _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06421_ _01566_ _01888_ _01889_ _01184_ _01890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_8_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09140_ _04173_ cpu.regs\[3\]\[0\] _04177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_6_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_6_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06352_ _01337_ _01781_ _01795_ _01821_ _01822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_16_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06283_ _01748_ _01750_ _01752_ _01753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09071_ cpu.orig_IO_addr_buff\[4\] _04106_ _04124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09632__A2 _04624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05303_ _00779_ _00801_ _00769_ _00802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08022_ _00621_ _03167_ net70 _03302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06207__B _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05234_ _00732_ _00735_ _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05165_ cpu.IE _00672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05096_ _00569_ _00606_ _00607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09973_ _02783_ _04919_ _04922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_73_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05957__A1 net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08924_ _04009_ _00401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08855_ cpu.timer\[9\] _03859_ _03891_ _03951_ _03952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_98_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08786_ _02717_ _03197_ _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07806_ cpu.regs\[3\]\[6\] _03099_ _03109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input13_I io_in[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05998_ _01467_ _01469_ _01470_ _01471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07552__I _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07737_ cpu.regs\[6\]\[4\] _03062_ _03066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09320__A1 _02340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07668_ _01922_ _03019_ _00135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06619_ _02076_ _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_07599_ _02975_ _02968_ _02976_ _00109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09407_ _04379_ _04344_ _04417_ _04380_ _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_118_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09338_ _04349_ _04351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_23_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09623__A2 _04238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05800__I _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09269_ _02669_ _02705_ _04284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09387__A1 _00983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output81_I net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06631__I _02097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10113_ net69 _05041_ _03334_ _05042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_101_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05247__I _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05263__I3 cpu.regs\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10044_ net78 _04977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_76_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_76_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_59_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05176__A2 cpu.ROM_spi_mode vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05100__A2 _00609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05157__I _00664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06970_ _02200_ _02434_ _02381_ _02379_ _02435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA_input5_I io_in[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05921_ _01343_ _01382_ _01395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_05852_ _01119_ _01299_ _01088_ _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08640_ _03790_ _03791_ _03792_ _00334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_83_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07372__I _00678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05167__A2 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05783_ _01250_ _01085_ _01257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08571_ cpu.toggle_top\[6\] _03722_ _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07522_ _02874_ _02922_ _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07453_ _02846_ _02859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06404_ _01207_ _01217_ cpu.PORTA_DDR\[5\] _01873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09123_ _00670_ _02129_ _04164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07384_ _02800_ _02801_ _02803_ _02697_ _00067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_8_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06335_ _01695_ _01718_ _01805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_17_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09054_ _00989_ _04096_ _04108_ _04109_ _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06266_ cpu.regs\[9\]\[3\] _01544_ _01737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08005_ cpu.spi.div_counter\[3\] _03289_ _03290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_103_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05217_ cpu.regs\[12\]\[2\] cpu.regs\[13\]\[2\] cpu.regs\[14\]\[2\] cpu.regs\[15\]\[2\]
+ _00683_ _00685_ _00720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08041__A1 _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06197_ _01663_ _01666_ _01667_ _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05493__I3 cpu.regs\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05148_ _00654_ _00656_ _00622_ _00010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_110_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09956_ cpu.PORTB_DDR\[0\] _04907_ _04909_ _04904_ _04910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08592__A2 _02053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05079_ cpu.instr_buff\[15\] _00590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08907_ _03995_ _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09887_ cpu.pwm_top\[0\] _03826_ _03828_ cpu.pwm_top\[2\] _04859_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_08838_ _02756_ _03859_ _03937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08895__A3 _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08769_ cpu.timer_top\[10\] _03877_ _03881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09144__I1 _03136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07855__A1 _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09002__I _04065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05530__I _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10662_ _00534_ clknet_leaf_55_wb_clk_i cpu.PORTB_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_118_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10593_ _00465_ clknet_leaf_78_wb_clk_i cpu.last_addr\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07607__A1 _02981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07083__A2 _02543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06361__I _01829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput51 net51 io_oeb[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput40 net40 io_oeb[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput73 net73 io_out[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput62 net62 io_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput84 net84 sram_addr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput95 net95 sram_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10027_ _04959_ _04962_ _04963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_90_Left_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_106_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05440__I _00917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06120_ _01591_ _01314_ _01098_ _01592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_112_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06051_ _01366_ _01385_ _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_117_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_99_Right_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09810_ _04755_ _04752_ _04796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09741_ _02519_ _02580_ _04694_ _04739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06953_ _02127_ _02419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05904_ _00839_ _00848_ _01378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08198__I _00677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09672_ cpu.orig_PC\[13\] _04089_ _04673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06337__A1 _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06884_ _02313_ _02349_ _02350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_89_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08623_ _03765_ _03764_ _03755_ _03775_ _03776_ _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05835_ _01308_ _01309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_27_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05766_ _01238_ _01239_ _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08554_ cpu.toggle_top\[0\] _03715_ _03716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07505_ cpu.uart.divisor\[0\] _02906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_81_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07830__I cpu.regs\[2\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07837__A1 _03136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05697_ _00598_ _01171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_65_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08485_ cpu.orig_flags\[0\] _03648_ _03667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_76_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05350__I _00829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06446__I _01914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07436_ _02836_ _02843_ _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_33_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07367_ _02788_ _02780_ _02789_ _02786_ _00064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_61_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09106_ _00908_ _04142_ _04151_ _04145_ _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_06318_ _01785_ _01787_ _01788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07298_ _02727_ _02732_ _00052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09037_ _04093_ _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06249_ _01132_ _01692_ _01719_ _01525_ _01720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_103_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06181__I net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09939_ _04897_ _00528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_99_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output44_I net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06328__A1 _01396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09117__I1 _02859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06500__B2 _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05260__I cpu.regs\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06356__I _01825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10645_ _00517_ clknet_leaf_60_wb_clk_i net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_106_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09667__I _04668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10576_ _00448_ clknet_leaf_81_wb_clk_i cpu.ROM_addr_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_91_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_91_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05209__I3 cpu.regs\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_20_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_20_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_30_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05620_ _01051_ _00593_ _00641_ _01094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_86_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05551_ _00604_ _01025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_80_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08270_ _03378_ _03500_ cpu.uart.div_counter\[15\] _03502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05170__I _00676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05482_ _00934_ _00937_ _00958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07221_ _02576_ _02663_ _02667_ _02666_ _00040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_30_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07152_ _02604_ _02605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06103_ cpu.timer_top\[10\] _01170_ _01468_ _01574_ _01575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__07097__I _00983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07083_ net1 _02543_ _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_42_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06034_ _01496_ _01507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07985_ cpu.spi.div_counter\[5\] cpu.spi.divisor\[5\] _03273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09724_ cpu.last_addr\[13\] _04723_ _04724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06936_ cpu.PC\[3\] _02402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_97_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05781__A2 _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06867_ _02325_ _02327_ _02318_ _02333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09655_ _04646_ _00879_ _04656_ _04657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_96_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05818_ _01278_ _01286_ _01291_ _01292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08606_ cpu.toggle_ctr\[2\] _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_96_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06798_ _02250_ _02262_ _02263_ _02264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09586_ _04585_ _04586_ _04589_ _04591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05749_ _01045_ _01010_ _01223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08537_ cpu.orig_PC\[11\] _03641_ _03704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06176__I _01421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08468_ _00599_ _03651_ _03652_ _03653_ _00301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_107_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07419_ cpu.PC\[0\] _02828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08399_ _02904_ _03599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_107_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10430_ _00303_ clknet_leaf_19_wb_clk_i cpu.orig_IO_addr_buff\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10361_ _00234_ clknet_leaf_63_wb_clk_i cpu.spi.counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10292_ _00165_ clknet_leaf_13_wb_clk_i cpu.regs\[5\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07470__I _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05524__A2 _00993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06721__A1 cpu.regs\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_114_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05383__S1 _00835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10628_ _00500_ clknet_leaf_76_wb_clk_i cpu.spi_clkdiv vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10033__A1 cpu.ROM_addr_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09974__A1 cpu.PORTB_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10559_ _00431_ clknet_leaf_54_wb_clk_i cpu.IO_addr_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07770_ _03085_ _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06721_ cpu.regs\[1\]\[4\] _00948_ _02187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_78_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09440_ _04329_ _04450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06652_ cpu.mem_cycle\[0\] _02118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07380__I _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05603_ _00598_ _01076_ _01077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_65_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06583_ cpu.pwm_top\[7\] _01049_ _01009_ _02050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09371_ _04377_ _04383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08322_ cpu.uart.data_buff\[5\] _03528_ _03542_ _03182_ _03543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05534_ _01007_ _01008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_47_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08253_ cpu.uart.div_counter\[12\] _03488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07204_ _02653_ _02654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_7_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05465_ _00934_ _00937_ _00939_ _00941_ _00942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_08184_ _02793_ _03432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05396_ _00820_ _00860_ _00875_ _00876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_42_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07135_ _02315_ _02587_ _02588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_113_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07066_ cpu.ROM_spi_dat_out\[7\] _02473_ _02528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06017_ _01483_ _01486_ _01489_ _01490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07968_ _03225_ _03244_ _03256_ _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09707_ cpu.last_addr\[8\] cpu.ROM_addr_buff\[8\] _04700_ _04707_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_4_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06919_ _02383_ _02384_ _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07899_ cpu.timer_div_counter\[0\] _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09638_ _04639_ _04640_ _04413_ _04641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_87_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09569_ _04402_ _04556_ _04574_ _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07223__C _02666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06482__A3 _01914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06634__I _01108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10413_ _00286_ clknet_leaf_36_wb_clk_i cpu.uart.receive_div_counter\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10344_ _00217_ clknet_leaf_46_wb_clk_i cpu.spi.data_in_buff\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07431__A2 _00979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10275_ _00148_ clknet_leaf_3_wb_clk_i cpu.regs\[7\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_49_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06170__A2 _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06544__I _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05250_ _00733_ _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07670__A2 _03019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05181_ _00685_ _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08940_ _04020_ _04022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07375__I _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08871_ _03965_ _00392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07822_ _03122_ _02407_ _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07753_ cpu.regs\[5\]\[1\] _03076_ _03077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_79_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07684_ cpu.regs\[8\]\[4\] _03025_ _03029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06704_ _02142_ _02169_ _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09423_ _04335_ _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06635_ _01101_ _02100_ _02101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09354_ _02859_ _03551_ _04292_ _04366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08438__A1 _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06566_ cpu.uart.divisor\[15\] _02033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08305_ cpu.uart.data_buff\[2\] _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_90_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05517_ _00662_ _00608_ _00609_ _00990_ _00991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_51_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06497_ _01959_ _01964_ _01625_ _01965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_35_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09285_ cpu.PC\[0\] _04298_ _04299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08236_ _03443_ _03475_ _03440_ _03476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05448_ _00925_ _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08167_ _03299_ _03418_ _03303_ _03419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09938__A1 net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07118_ _02573_ _02574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05379_ _00858_ _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_30_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08098_ _03350_ _03358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07049_ _02483_ _02485_ _02510_ _02511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_30_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10060_ _02514_ _04992_ _04993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_89_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07101__A1 _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09929__A1 _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10327_ _00200_ clknet_leaf_63_wb_clk_i cpu.spi.div_counter\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05966__A2 _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10258_ _00131_ clknet_leaf_1_wb_clk_i cpu.regs\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07923__I cpu.timer_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10189_ _00066_ clknet_leaf_15_wb_clk_i cpu.toggle_top\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_109_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06420_ cpu.spi.dout\[5\] _01188_ _01889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_118_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06351_ _01799_ _01814_ _01820_ _01821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_06282_ _01191_ _01751_ _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09070_ _04095_ _04123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05302_ cpu.regs\[0\]\[6\] _00800_ cpu.regs\[2\]\[6\] cpu.regs\[3\]\[6\] _00788_
+ _00789_ _00801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_114_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08021_ _03300_ _03301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05233_ cpu.regs\[12\]\[3\] cpu.regs\[13\]\[3\] cpu.regs\[14\]\[3\] cpu.regs\[15\]\[3\]
+ _00733_ _00734_ _00735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05654__A1 _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05164_ _00657_ _00661_ _00667_ _00671_ _00008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_40_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05095_ _00602_ _00605_ _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09972_ _04921_ _00537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05406__A1 _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05957__A2 _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09148__A2 cpu.regs\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08923_ cpu.timer_capture\[12\] _04003_ _04008_ _03998_ _04009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_110_Left_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08854_ _03198_ _03950_ _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08785_ _03890_ _03891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05997_ cpu.pwm_top\[1\] _01269_ _01168_ _01470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07805_ _01921_ _03101_ _03108_ _00183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07736_ _03047_ _03059_ _03065_ _00157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_94_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07667_ _01827_ _03019_ _00134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07598_ cpu.regs\[12\]\[3\] _02969_ _02976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06618_ _01165_ _01391_ _02065_ _01383_ _01398_ _02085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_09406_ cpu.PC\[2\] cpu.br_rel_dest\[2\] _04417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09084__A1 _01924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09337_ _04349_ _04350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06549_ _02016_ _02017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_23_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09268_ _04266_ _04281_ _04282_ _04283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08219_ _03461_ _03462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09199_ cpu.ROM_addr_buff\[7\] _04213_ _04223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09387__A2 _03310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05660__A4 _00637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output74_I net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10112_ _03416_ _05040_ _00666_ _05041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10043_ _04972_ _04976_ _02683_ _00553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07743__I _03058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06373__A2 _01841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_45_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_45_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_85_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07389__A1 cpu.toggle_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05495__S0 _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05920_ _01339_ _01380_ _01394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05851_ _01261_ _01324_ _01075_ _01257_ _01325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_107_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08570_ _02811_ _03721_ _03726_ _03725_ _00330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__07561__A1 _02098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07521_ _02919_ _02921_ _02922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05782_ _01255_ _01256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09302__A2 _04314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07452_ _01686_ _01732_ _01733_ _02858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09066__A1 _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06403_ cpu.toggle_top\[5\] _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07383_ cpu.toggle_top\[9\] _02802_ _02803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09122_ _04163_ _00445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06334_ _01797_ _01803_ _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05627__A1 _00647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09053_ _04083_ _04109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06265_ _01735_ _01736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08004_ _03287_ _03288_ _03289_ _00201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06196_ cpu.spi.divisor\[3\] _01244_ _01188_ _01667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05216_ cpu.regs\[8\]\[2\] cpu.regs\[9\]\[2\] cpu.regs\[10\]\[2\] cpu.regs\[11\]\[2\]
+ _00684_ _00712_ _00719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_05147_ _00616_ _00655_ _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_110_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09955_ _02670_ _04908_ _04909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05078_ cpu.base_address\[1\] _00588_ _00589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08906_ cpu.timer_capture\[9\] _03986_ _03994_ _03979_ _03995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09886_ cpu.pwm_top\[1\] _03827_ _03828_ cpu.pwm_top\[2\] _04857_ _04858_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08837_ _03936_ _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07563__I _02951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08768_ _02769_ _03876_ _03880_ _03879_ _00374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_95_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08699_ cpu.pwm_counter\[4\] _03830_ _03709_ _03833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_0_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_0_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07719_ cpu.regs\[7\]\[6\] _03038_ _03054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10661_ _00533_ clknet_leaf_56_wb_clk_i cpu.PORTB_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_36_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10592_ _00464_ clknet_leaf_80_wb_clk_i cpu.last_addr\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05618__A1 _01000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput52 net52 io_oeb[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput41 net41 io_oeb[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput74 net74 io_out[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput63 net63 io_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09780__A2 _04771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput85 net85 sram_addr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput96 net96 sram_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10026_ cpu.ROM_addr_buff\[4\] _02523_ _02524_ cpu.ROM_addr_buff\[8\] cpu.ROM_addr_buff\[12\]
+ _04961_ _04962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__10113__B _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_20_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07406__C _02818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06552__I _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06050_ _01522_ _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_117_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09740_ _02580_ _04692_ _02519_ _04738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08479__I _03662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06585__A2 _01416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06952_ _02413_ _02416_ _02417_ _02418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
.ends

