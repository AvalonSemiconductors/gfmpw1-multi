magic
tech gf180mcuD
magscale 1 10
timestamp 1753965644
<< metal1 >>
rect 1344 36874 38640 36908
rect 1344 36822 5876 36874
rect 5928 36822 5980 36874
rect 6032 36822 6084 36874
rect 6136 36822 15200 36874
rect 15252 36822 15304 36874
rect 15356 36822 15408 36874
rect 15460 36822 24524 36874
rect 24576 36822 24628 36874
rect 24680 36822 24732 36874
rect 24784 36822 33848 36874
rect 33900 36822 33952 36874
rect 34004 36822 34056 36874
rect 34108 36822 38640 36874
rect 1344 36788 38640 36822
rect 19182 36706 19234 36718
rect 19182 36642 19234 36654
rect 37606 36594 37658 36606
rect 33170 36542 33182 36594
rect 33234 36542 33246 36594
rect 37606 36530 37658 36542
rect 13694 36482 13746 36494
rect 17390 36482 17442 36494
rect 23550 36482 23602 36494
rect 10210 36402 10222 36454
rect 10274 36402 10286 36454
rect 12338 36430 12350 36482
rect 12402 36430 12414 36482
rect 13694 36418 13746 36430
rect 13906 36402 13918 36454
rect 13970 36402 13982 36454
rect 16146 36430 16158 36482
rect 16210 36430 16222 36482
rect 17390 36418 17442 36430
rect 19842 36402 19854 36454
rect 19906 36402 19918 36454
rect 22754 36430 22766 36482
rect 22818 36430 22830 36482
rect 27246 36482 27298 36494
rect 31054 36482 31106 36494
rect 23550 36418 23602 36430
rect 24546 36402 24558 36454
rect 24610 36402 24622 36454
rect 28578 36430 28590 36482
rect 28642 36430 28654 36482
rect 27246 36418 27298 36430
rect 30706 36402 30718 36454
rect 30770 36402 30782 36454
rect 35422 36482 35474 36494
rect 31054 36418 31106 36430
rect 32498 36402 32510 36454
rect 32562 36402 32574 36454
rect 35422 36418 35474 36430
rect 38334 36482 38386 36494
rect 38334 36418 38386 36430
rect 20862 36370 20914 36382
rect 3446 36314 3498 36326
rect 3446 36250 3498 36262
rect 4566 36314 4618 36326
rect 4566 36250 4618 36262
rect 5686 36314 5738 36326
rect 5686 36250 5738 36262
rect 6806 36314 6858 36326
rect 6806 36250 6858 36262
rect 7926 36314 7978 36326
rect 7926 36250 7978 36262
rect 8710 36314 8762 36326
rect 8710 36250 8762 36262
rect 9718 36314 9770 36326
rect 20862 36306 20914 36318
rect 36150 36370 36202 36382
rect 36150 36306 36202 36318
rect 9718 36250 9770 36262
rect 13358 36258 13410 36270
rect 13358 36194 13410 36206
rect 17054 36258 17106 36270
rect 17054 36194 17106 36206
rect 23942 36258 23994 36270
rect 23942 36194 23994 36206
rect 25902 36258 25954 36270
rect 25902 36194 25954 36206
rect 27582 36258 27634 36270
rect 27582 36194 27634 36206
rect 31390 36258 31442 36270
rect 31390 36194 31442 36206
rect 35086 36258 35138 36270
rect 35086 36194 35138 36206
rect 37998 36258 38050 36270
rect 37998 36194 38050 36206
rect 1344 36090 38800 36124
rect 1344 36038 10538 36090
rect 10590 36038 10642 36090
rect 10694 36038 10746 36090
rect 10798 36038 19862 36090
rect 19914 36038 19966 36090
rect 20018 36038 20070 36090
rect 20122 36038 29186 36090
rect 29238 36038 29290 36090
rect 29342 36038 29394 36090
rect 29446 36038 38510 36090
rect 38562 36038 38614 36090
rect 38666 36038 38718 36090
rect 38770 36038 38800 36090
rect 1344 36004 38800 36038
rect 11286 35922 11338 35934
rect 11286 35858 11338 35870
rect 30942 35922 30994 35934
rect 30942 35858 30994 35870
rect 8878 35810 8930 35822
rect 8878 35746 8930 35758
rect 20974 35810 21026 35822
rect 16270 35737 16322 35749
rect 20974 35746 21026 35758
rect 2494 35698 2546 35710
rect 2494 35634 2546 35646
rect 5798 35698 5850 35710
rect 5798 35634 5850 35646
rect 6190 35698 6242 35710
rect 6190 35634 6242 35646
rect 12238 35698 12290 35710
rect 12238 35634 12290 35646
rect 12350 35698 12402 35710
rect 12350 35634 12402 35646
rect 15710 35698 15762 35710
rect 15710 35634 15762 35646
rect 16046 35698 16098 35710
rect 17278 35698 17330 35710
rect 16270 35673 16322 35685
rect 16594 35646 16606 35698
rect 16658 35646 16670 35698
rect 16046 35634 16098 35646
rect 17278 35634 17330 35646
rect 23662 35698 23714 35710
rect 23662 35634 23714 35646
rect 24782 35698 24834 35710
rect 25218 35673 25230 35725
rect 25282 35673 25294 35725
rect 28018 35673 28030 35725
rect 28082 35673 28094 35725
rect 31278 35698 31330 35710
rect 24782 35634 24834 35646
rect 31278 35634 31330 35646
rect 31726 35698 31778 35710
rect 33058 35673 33070 35725
rect 33122 35673 33134 35725
rect 35758 35698 35810 35710
rect 31726 35634 31778 35646
rect 35758 35634 35810 35646
rect 36430 35698 36482 35710
rect 36430 35634 36482 35646
rect 9718 35586 9770 35598
rect 3266 35534 3278 35586
rect 3330 35534 3342 35586
rect 5170 35534 5182 35586
rect 5234 35534 5246 35586
rect 6962 35534 6974 35586
rect 7026 35534 7038 35586
rect 9718 35522 9770 35534
rect 10950 35586 11002 35598
rect 20582 35586 20634 35598
rect 24054 35586 24106 35598
rect 13122 35534 13134 35586
rect 13186 35534 13198 35586
rect 15026 35534 15038 35586
rect 15090 35534 15102 35586
rect 16482 35534 16494 35586
rect 16546 35534 16558 35586
rect 18050 35534 18062 35586
rect 18114 35534 18126 35586
rect 19954 35534 19966 35586
rect 20018 35534 20030 35586
rect 22866 35534 22878 35586
rect 22930 35534 22942 35586
rect 10950 35522 11002 35534
rect 20582 35522 20634 35534
rect 24054 35522 24106 35534
rect 11902 35474 11954 35486
rect 11902 35410 11954 35422
rect 24446 35474 24498 35486
rect 24446 35410 24498 35422
rect 26238 35474 26290 35486
rect 26238 35410 26290 35422
rect 29038 35474 29090 35486
rect 29038 35410 29090 35422
rect 32062 35474 32114 35486
rect 32062 35410 32114 35422
rect 34414 35474 34466 35486
rect 34414 35410 34466 35422
rect 36094 35474 36146 35486
rect 36094 35410 36146 35422
rect 36766 35474 36818 35486
rect 36766 35410 36818 35422
rect 1344 35306 38640 35340
rect 1344 35254 5876 35306
rect 5928 35254 5980 35306
rect 6032 35254 6084 35306
rect 6136 35254 15200 35306
rect 15252 35254 15304 35306
rect 15356 35254 15408 35306
rect 15460 35254 24524 35306
rect 24576 35254 24628 35306
rect 24680 35254 24732 35306
rect 24784 35254 33848 35306
rect 33900 35254 33952 35306
rect 34004 35254 34056 35306
rect 34108 35254 38640 35306
rect 1344 35220 38640 35254
rect 2942 35138 2994 35150
rect 2942 35074 2994 35086
rect 8766 35138 8818 35150
rect 8766 35074 8818 35086
rect 15374 35138 15426 35150
rect 15374 35074 15426 35086
rect 22318 35138 22370 35150
rect 22318 35074 22370 35086
rect 24334 35138 24386 35150
rect 24334 35074 24386 35086
rect 9494 35026 9546 35038
rect 9494 34962 9546 34974
rect 9942 35026 9994 35038
rect 19966 35026 20018 35038
rect 12786 34974 12798 35026
rect 12850 34974 12862 35026
rect 16706 34974 16718 35026
rect 16770 34974 16782 35026
rect 9942 34962 9994 34974
rect 19966 34962 20018 34974
rect 20806 35026 20858 35038
rect 25778 34974 25790 35026
rect 25842 34974 25854 35026
rect 20806 34962 20858 34974
rect 4062 34914 4114 34926
rect 4062 34850 4114 34862
rect 5518 34914 5570 34926
rect 9102 34914 9154 34926
rect 6290 34862 6302 34914
rect 6354 34862 6366 34914
rect 5518 34850 5570 34862
rect 9102 34850 9154 34862
rect 10110 34914 10162 34926
rect 13750 34914 13802 34926
rect 10882 34862 10894 34914
rect 10946 34862 10958 34914
rect 10110 34850 10162 34862
rect 13750 34850 13802 34862
rect 13918 34914 13970 34926
rect 13918 34850 13970 34862
rect 15934 34914 15986 34926
rect 15934 34850 15986 34862
rect 19630 34914 19682 34926
rect 23998 34914 24050 34926
rect 20290 34862 20302 34914
rect 20354 34862 20366 34914
rect 19630 34850 19682 34862
rect 8206 34802 8258 34814
rect 8206 34738 8258 34750
rect 18622 34802 18674 34814
rect 19954 34806 19966 34858
rect 20018 34806 20030 34858
rect 21522 34834 21534 34886
rect 21586 34834 21598 34886
rect 23998 34850 24050 34862
rect 25006 34914 25058 34926
rect 25006 34850 25058 34862
rect 28030 34914 28082 34926
rect 28030 34850 28082 34862
rect 28254 34914 28306 34926
rect 29038 34914 29090 34926
rect 31054 34914 31106 34926
rect 34638 34914 34690 34926
rect 28522 34862 28534 34914
rect 28586 34862 28598 34914
rect 30482 34862 30494 34914
rect 30546 34862 30558 34914
rect 31826 34862 31838 34914
rect 31890 34862 31902 34914
rect 28254 34850 28306 34862
rect 29038 34850 29090 34862
rect 31054 34850 31106 34862
rect 34638 34850 34690 34862
rect 35310 34914 35362 34926
rect 35310 34850 35362 34862
rect 35422 34914 35474 34926
rect 35422 34850 35474 34862
rect 18622 34738 18674 34750
rect 27694 34802 27746 34814
rect 27694 34738 27746 34750
rect 33742 34802 33794 34814
rect 33742 34738 33794 34750
rect 36374 34802 36426 34814
rect 36374 34738 36426 34750
rect 34302 34690 34354 34702
rect 34302 34626 34354 34638
rect 34974 34690 35026 34702
rect 34974 34626 35026 34638
rect 35758 34690 35810 34702
rect 35758 34626 35810 34638
rect 37830 34690 37882 34702
rect 37830 34626 37882 34638
rect 38278 34690 38330 34702
rect 38278 34626 38330 34638
rect 1344 34522 38800 34556
rect 1344 34470 10538 34522
rect 10590 34470 10642 34522
rect 10694 34470 10746 34522
rect 10798 34470 19862 34522
rect 19914 34470 19966 34522
rect 20018 34470 20070 34522
rect 20122 34470 29186 34522
rect 29238 34470 29290 34522
rect 29342 34470 29394 34522
rect 29446 34470 38510 34522
rect 38562 34470 38614 34522
rect 38666 34470 38718 34522
rect 38770 34470 38800 34522
rect 1344 34436 38800 34470
rect 5966 34354 6018 34366
rect 5966 34290 6018 34302
rect 10894 34354 10946 34366
rect 10894 34290 10946 34302
rect 15710 34354 15762 34366
rect 18790 34354 18842 34366
rect 15710 34290 15762 34302
rect 17950 34298 18002 34310
rect 18790 34290 18842 34302
rect 20414 34354 20466 34366
rect 20414 34290 20466 34302
rect 17950 34234 18002 34246
rect 28926 34242 28978 34254
rect 17838 34169 17890 34181
rect 28926 34178 28978 34190
rect 7086 34130 7138 34142
rect 8878 34130 8930 34142
rect 8586 34078 8598 34130
rect 8650 34078 8662 34130
rect 7086 34066 7138 34078
rect 8878 34066 8930 34078
rect 8990 34130 9042 34142
rect 8990 34066 9042 34078
rect 9438 34130 9490 34142
rect 11778 34105 11790 34157
rect 11842 34105 11854 34157
rect 14354 34105 14366 34157
rect 14418 34105 14430 34157
rect 17614 34130 17666 34142
rect 9438 34066 9490 34078
rect 17838 34105 17890 34117
rect 18162 34078 18174 34130
rect 18226 34078 18238 34130
rect 19058 34105 19070 34157
rect 19122 34105 19134 34157
rect 21870 34130 21922 34142
rect 28254 34130 28306 34142
rect 27458 34078 27470 34130
rect 27522 34078 27534 34130
rect 17614 34066 17666 34078
rect 21870 34066 21922 34078
rect 28254 34066 28306 34078
rect 31614 34130 31666 34142
rect 31614 34066 31666 34078
rect 31726 34130 31778 34142
rect 31726 34066 31778 34078
rect 32958 34130 33010 34142
rect 36262 34130 36314 34142
rect 33730 34078 33742 34130
rect 33794 34078 33806 34130
rect 32958 34066 33010 34078
rect 36262 34066 36314 34078
rect 37662 34130 37714 34142
rect 37662 34066 37714 34078
rect 38334 34130 38386 34142
rect 38334 34066 38386 34078
rect 32062 34018 32114 34030
rect 36710 34018 36762 34030
rect 12562 33966 12574 34018
rect 12626 33966 12638 34018
rect 22642 33966 22654 34018
rect 22706 33966 22718 34018
rect 24546 33966 24558 34018
rect 24610 33966 24622 34018
rect 25554 33966 25566 34018
rect 25618 33966 25630 34018
rect 30818 33966 30830 34018
rect 30882 33966 30894 34018
rect 35634 33966 35646 34018
rect 35698 33966 35710 34018
rect 32062 33954 32114 33966
rect 36710 33954 36762 33966
rect 37326 34018 37378 34030
rect 37326 33954 37378 33966
rect 37998 33906 38050 33918
rect 7410 33854 7422 33906
rect 7474 33903 7486 33906
rect 7746 33903 7758 33906
rect 7474 33857 7758 33903
rect 7474 33854 7486 33857
rect 7746 33854 7758 33857
rect 7810 33854 7822 33906
rect 37998 33842 38050 33854
rect 1344 33738 38640 33772
rect 1344 33686 5876 33738
rect 5928 33686 5980 33738
rect 6032 33686 6084 33738
rect 6136 33686 15200 33738
rect 15252 33686 15304 33738
rect 15356 33686 15408 33738
rect 15460 33686 24524 33738
rect 24576 33686 24628 33738
rect 24680 33686 24732 33738
rect 24784 33686 33848 33738
rect 33900 33686 33952 33738
rect 34004 33686 34056 33738
rect 34108 33686 38640 33738
rect 1344 33652 38640 33686
rect 16158 33570 16210 33582
rect 9034 33518 9046 33570
rect 9098 33518 9110 33570
rect 14746 33518 14758 33570
rect 14810 33518 14822 33570
rect 16158 33506 16210 33518
rect 18958 33570 19010 33582
rect 18958 33506 19010 33518
rect 22654 33570 22706 33582
rect 22654 33506 22706 33518
rect 25678 33570 25730 33582
rect 25678 33506 25730 33518
rect 10446 33458 10498 33470
rect 30588 33458 30640 33470
rect 12338 33406 12350 33458
rect 12402 33406 12414 33458
rect 10446 33394 10498 33406
rect 30588 33394 30640 33406
rect 31334 33402 31386 33414
rect 32498 33406 32510 33458
rect 32562 33406 32574 33458
rect 8766 33346 8818 33358
rect 8766 33282 8818 33294
rect 9326 33346 9378 33358
rect 9326 33282 9378 33294
rect 9438 33346 9490 33358
rect 9438 33282 9490 33294
rect 10054 33346 10106 33358
rect 10054 33282 10106 33294
rect 10782 33346 10834 33358
rect 10782 33282 10834 33294
rect 11454 33346 11506 33358
rect 11454 33282 11506 33294
rect 11902 33346 11954 33358
rect 13806 33346 13858 33358
rect 12450 33294 12462 33346
rect 12514 33294 12526 33346
rect 11902 33282 11954 33294
rect 12226 33238 12238 33290
rect 12290 33238 12302 33290
rect 13806 33282 13858 33294
rect 13918 33346 13970 33358
rect 13918 33282 13970 33294
rect 14254 33346 14306 33358
rect 14254 33282 14306 33294
rect 14478 33346 14530 33358
rect 22150 33346 22202 33358
rect 14478 33282 14530 33294
rect 15474 33266 15486 33318
rect 15538 33266 15550 33318
rect 17938 33266 17950 33318
rect 18002 33266 18014 33318
rect 21310 33290 21362 33302
rect 13514 33182 13526 33234
rect 13578 33182 13590 33234
rect 21310 33226 21362 33238
rect 21422 33290 21474 33302
rect 22150 33282 22202 33294
rect 22318 33346 22370 33358
rect 22318 33282 22370 33294
rect 22990 33346 23042 33358
rect 22990 33282 23042 33294
rect 25006 33346 25058 33358
rect 25284 33346 25336 33358
rect 25106 33294 25118 33346
rect 25170 33294 25182 33346
rect 27806 33346 27858 33358
rect 25006 33282 25058 33294
rect 25284 33282 25336 33294
rect 26450 33266 26462 33318
rect 26514 33266 26526 33318
rect 27806 33282 27858 33294
rect 29822 33346 29874 33358
rect 21422 33226 21474 33238
rect 21982 33234 22034 33246
rect 21982 33170 22034 33182
rect 24278 33234 24330 33246
rect 24278 33170 24330 33182
rect 29150 33234 29202 33246
rect 29306 33238 29318 33290
rect 29370 33238 29382 33290
rect 29822 33282 29874 33294
rect 30830 33346 30882 33358
rect 35534 33402 35586 33414
rect 31334 33338 31386 33350
rect 31726 33346 31778 33358
rect 30830 33282 30882 33294
rect 35534 33338 35586 33350
rect 37662 33346 37714 33358
rect 31726 33282 31778 33294
rect 29150 33170 29202 33182
rect 30064 33234 30116 33246
rect 30064 33170 30116 33182
rect 31502 33234 31554 33246
rect 31502 33170 31554 33182
rect 34414 33234 34466 33246
rect 34414 33170 34466 33182
rect 34862 33234 34914 33246
rect 35018 33238 35030 33290
rect 35082 33238 35094 33290
rect 34862 33170 34914 33182
rect 35776 33234 35828 33246
rect 35776 33170 35828 33182
rect 36990 33234 37042 33246
rect 37146 33238 37158 33290
rect 37210 33238 37222 33290
rect 37662 33282 37714 33294
rect 36990 33170 37042 33182
rect 37904 33234 37956 33246
rect 37904 33170 37956 33182
rect 8430 33122 8482 33134
rect 8430 33058 8482 33070
rect 11118 33122 11170 33134
rect 11118 33058 11170 33070
rect 23326 33122 23378 33134
rect 23326 33058 23378 33070
rect 24726 33122 24778 33134
rect 24726 33058 24778 33070
rect 36374 33122 36426 33134
rect 36374 33058 36426 33070
rect 1344 32954 38800 32988
rect 1344 32902 10538 32954
rect 10590 32902 10642 32954
rect 10694 32902 10746 32954
rect 10798 32902 19862 32954
rect 19914 32902 19966 32954
rect 20018 32902 20070 32954
rect 20122 32902 29186 32954
rect 29238 32902 29290 32954
rect 29342 32902 29394 32954
rect 29446 32902 38510 32954
rect 38562 32902 38614 32954
rect 38666 32902 38718 32954
rect 38770 32902 38800 32954
rect 1344 32868 38800 32902
rect 5686 32786 5738 32798
rect 5686 32722 5738 32734
rect 13022 32786 13074 32798
rect 13022 32722 13074 32734
rect 24278 32786 24330 32798
rect 29710 32786 29762 32798
rect 9606 32674 9658 32686
rect 9606 32610 9658 32622
rect 17502 32674 17554 32686
rect 18834 32678 18846 32730
rect 18898 32678 18910 32730
rect 24278 32722 24330 32734
rect 24614 32730 24666 32742
rect 2382 32562 2434 32574
rect 7186 32510 7198 32562
rect 7250 32510 7262 32562
rect 7746 32510 7758 32562
rect 7810 32510 7822 32562
rect 8082 32525 8094 32577
rect 8146 32525 8158 32577
rect 8430 32562 8482 32574
rect 2382 32498 2434 32510
rect 8430 32498 8482 32510
rect 8654 32562 8706 32574
rect 9874 32566 9886 32618
rect 9938 32566 9950 32618
rect 17502 32610 17554 32622
rect 19630 32674 19682 32686
rect 10110 32590 10162 32602
rect 10110 32526 10162 32538
rect 10334 32590 10386 32602
rect 10334 32526 10386 32538
rect 10490 32526 10502 32578
rect 10554 32526 10566 32578
rect 10882 32510 10894 32562
rect 10946 32510 10958 32562
rect 11106 32510 11118 32562
rect 11170 32510 11182 32562
rect 11666 32510 11678 32562
rect 11730 32510 11742 32562
rect 11890 32525 11902 32577
rect 11954 32525 11966 32577
rect 14142 32562 14194 32574
rect 14354 32510 14366 32562
rect 14418 32510 14430 32562
rect 14690 32510 14702 32562
rect 14754 32510 14766 32562
rect 15698 32510 15710 32562
rect 15762 32510 15774 32562
rect 15922 32525 15934 32577
rect 15986 32525 15998 32577
rect 16482 32525 16494 32577
rect 16546 32525 16558 32577
rect 17838 32562 17890 32574
rect 16706 32510 16718 32562
rect 16770 32510 16782 32562
rect 18050 32510 18062 32562
rect 18114 32510 18126 32562
rect 18386 32537 18398 32589
rect 18450 32537 18462 32589
rect 18734 32562 18786 32574
rect 8654 32498 8706 32510
rect 14142 32498 14194 32510
rect 17838 32498 17890 32510
rect 18734 32498 18786 32510
rect 19294 32562 19346 32574
rect 19450 32566 19462 32618
rect 19514 32566 19526 32618
rect 19630 32610 19682 32622
rect 22990 32674 23042 32686
rect 29710 32722 29762 32734
rect 24614 32666 24666 32678
rect 20672 32600 20724 32612
rect 19294 32498 19346 32510
rect 19742 32562 19794 32574
rect 19742 32498 19794 32510
rect 20022 32562 20074 32574
rect 20022 32498 20074 32510
rect 20414 32562 20466 32574
rect 20514 32510 20526 32562
rect 20578 32510 20590 32562
rect 20672 32536 20724 32548
rect 21422 32562 21474 32574
rect 20414 32498 20466 32510
rect 21422 32498 21474 32510
rect 21646 32562 21698 32574
rect 22586 32566 22598 32618
rect 22650 32566 22662 32618
rect 22990 32610 23042 32622
rect 23158 32618 23210 32630
rect 26294 32618 26346 32630
rect 31434 32622 31446 32674
rect 31498 32622 31510 32674
rect 22754 32510 22766 32562
rect 22818 32510 22830 32562
rect 23158 32554 23210 32566
rect 23650 32510 23662 32562
rect 23714 32510 23726 32562
rect 24770 32510 24782 32562
rect 24834 32510 24846 32562
rect 25666 32538 25678 32590
rect 25730 32538 25742 32590
rect 25890 32510 25902 32562
rect 25954 32510 25966 32562
rect 26294 32554 26346 32566
rect 26574 32562 26626 32574
rect 26674 32510 26686 32562
rect 26738 32510 26750 32562
rect 26832 32560 26844 32612
rect 26896 32560 26908 32612
rect 28018 32537 28030 32589
rect 28082 32537 28094 32589
rect 30942 32562 30994 32574
rect 21646 32498 21698 32510
rect 26574 32498 26626 32510
rect 30942 32498 30994 32510
rect 31166 32562 31218 32574
rect 31166 32498 31218 32510
rect 31950 32562 32002 32574
rect 31950 32498 32002 32510
rect 32174 32562 32226 32574
rect 32174 32498 32226 32510
rect 35198 32562 35250 32574
rect 35198 32498 35250 32510
rect 35310 32562 35362 32574
rect 35310 32498 35362 32510
rect 15318 32450 15370 32462
rect 21086 32450 21138 32462
rect 3154 32398 3166 32450
rect 3218 32398 3230 32450
rect 5058 32398 5070 32450
rect 5122 32398 5134 32450
rect 7366 32394 7418 32406
rect 8194 32398 8206 32450
rect 8258 32398 8270 32450
rect 7366 32330 7418 32342
rect 11230 32394 11282 32406
rect 12002 32398 12014 32450
rect 12066 32398 12078 32450
rect 16034 32398 16046 32450
rect 16098 32398 16110 32450
rect 16370 32398 16382 32450
rect 16434 32398 16446 32450
rect 14690 32342 14702 32394
rect 14754 32342 14766 32394
rect 15318 32386 15370 32398
rect 21086 32386 21138 32398
rect 26126 32450 26178 32462
rect 26126 32386 26178 32398
rect 27246 32450 27298 32462
rect 27246 32386 27298 32398
rect 34078 32450 34130 32462
rect 36082 32398 36094 32450
rect 36146 32398 36158 32450
rect 37986 32398 37998 32450
rect 38050 32398 38062 32450
rect 34078 32386 34130 32398
rect 8922 32286 8934 32338
rect 8986 32286 8998 32338
rect 11230 32330 11282 32342
rect 23494 32338 23546 32350
rect 21914 32286 21926 32338
rect 21978 32286 21990 32338
rect 32442 32286 32454 32338
rect 32506 32286 32518 32338
rect 23494 32274 23546 32286
rect 1344 32170 38640 32204
rect 1344 32118 5876 32170
rect 5928 32118 5980 32170
rect 6032 32118 6084 32170
rect 6136 32118 15200 32170
rect 15252 32118 15304 32170
rect 15356 32118 15408 32170
rect 15460 32118 24524 32170
rect 24576 32118 24628 32170
rect 24680 32118 24732 32170
rect 24784 32118 33848 32170
rect 33900 32118 33952 32170
rect 34004 32118 34056 32170
rect 34108 32118 38640 32170
rect 1344 32084 38640 32118
rect 3166 32002 3218 32014
rect 3166 31938 3218 31950
rect 11118 32002 11170 32014
rect 11118 31938 11170 31950
rect 14310 32002 14362 32014
rect 14310 31938 14362 31950
rect 22766 32002 22818 32014
rect 22766 31938 22818 31950
rect 25230 32002 25282 32014
rect 25230 31938 25282 31950
rect 9344 31890 9396 31902
rect 8598 31834 8650 31846
rect 4286 31778 4338 31790
rect 4286 31714 4338 31726
rect 4398 31778 4450 31790
rect 4398 31714 4450 31726
rect 4622 31778 4674 31790
rect 4622 31714 4674 31726
rect 7758 31778 7810 31790
rect 7086 31666 7138 31678
rect 7242 31670 7254 31722
rect 7306 31670 7318 31722
rect 7758 31714 7810 31726
rect 8000 31778 8052 31790
rect 9344 31826 9396 31838
rect 9830 31890 9882 31902
rect 34190 31890 34242 31902
rect 16706 31838 16718 31890
rect 16770 31838 16782 31890
rect 19954 31838 19966 31890
rect 20018 31838 20030 31890
rect 24210 31838 24222 31890
rect 24274 31838 24286 31890
rect 29138 31838 29150 31890
rect 29202 31838 29214 31890
rect 31490 31838 31502 31890
rect 31554 31838 31566 31890
rect 35914 31838 35926 31890
rect 35978 31838 35990 31890
rect 9830 31826 9882 31838
rect 34190 31826 34242 31838
rect 8598 31770 8650 31782
rect 9102 31778 9154 31790
rect 11790 31778 11842 31790
rect 8000 31714 8052 31726
rect 9102 31714 9154 31726
rect 10110 31750 10162 31762
rect 10558 31750 10610 31762
rect 10110 31686 10162 31698
rect 4890 31614 4902 31666
rect 4954 31614 4966 31666
rect 7086 31602 7138 31614
rect 8430 31666 8482 31678
rect 10322 31670 10334 31722
rect 10386 31670 10398 31722
rect 10714 31710 10726 31762
rect 10778 31710 10790 31762
rect 11666 31726 11678 31778
rect 11730 31726 11742 31778
rect 10558 31686 10610 31698
rect 11498 31670 11510 31722
rect 11562 31670 11574 31722
rect 11790 31714 11842 31726
rect 12126 31778 12178 31790
rect 14590 31778 14642 31790
rect 12674 31726 12686 31778
rect 12738 31726 12750 31778
rect 14030 31750 14082 31762
rect 12126 31714 12178 31726
rect 13470 31722 13522 31734
rect 13570 31670 13582 31722
rect 13634 31670 13646 31722
rect 13794 31670 13806 31722
rect 13858 31670 13870 31722
rect 14590 31714 14642 31726
rect 14814 31778 14866 31790
rect 14814 31714 14866 31726
rect 15822 31778 15874 31790
rect 15822 31714 15874 31726
rect 15934 31778 15986 31790
rect 17278 31778 17330 31790
rect 20302 31778 20354 31790
rect 16258 31726 16270 31778
rect 16322 31726 16334 31778
rect 15934 31714 15986 31726
rect 14030 31686 14082 31698
rect 16594 31682 16606 31734
rect 16658 31682 16670 31734
rect 18050 31726 18062 31778
rect 18114 31726 18126 31778
rect 17278 31714 17330 31726
rect 20302 31714 20354 31726
rect 22094 31778 22146 31790
rect 22374 31778 22426 31790
rect 22194 31726 22206 31778
rect 22258 31726 22270 31778
rect 22094 31714 22146 31726
rect 22374 31714 22426 31726
rect 23438 31778 23490 31790
rect 23438 31714 23490 31726
rect 23774 31778 23826 31790
rect 25566 31778 25618 31790
rect 36206 31778 36258 31790
rect 24322 31726 24334 31778
rect 24386 31726 24398 31778
rect 23774 31714 23826 31726
rect 24098 31670 24110 31722
rect 24162 31670 24174 31722
rect 25566 31714 25618 31726
rect 26002 31698 26014 31750
rect 26066 31698 26078 31750
rect 29250 31711 29262 31763
rect 29314 31711 29326 31763
rect 29474 31726 29486 31778
rect 29538 31726 29550 31778
rect 32274 31698 32286 31750
rect 32338 31698 32350 31750
rect 32834 31698 32846 31750
rect 32898 31698 32910 31750
rect 36206 31714 36258 31726
rect 36318 31778 36370 31790
rect 36318 31714 36370 31726
rect 37158 31778 37210 31790
rect 37158 31714 37210 31726
rect 37662 31778 37714 31790
rect 37662 31714 37714 31726
rect 13470 31658 13522 31670
rect 36990 31666 37042 31678
rect 15082 31614 15094 31666
rect 15146 31614 15158 31666
rect 15530 31614 15542 31666
rect 15594 31614 15606 31666
rect 8430 31602 8482 31614
rect 12562 31558 12574 31610
rect 12626 31558 12638 31610
rect 36990 31602 37042 31614
rect 37904 31666 37956 31678
rect 37904 31602 37956 31614
rect 20638 31554 20690 31566
rect 20638 31490 20690 31502
rect 1344 31386 38800 31420
rect 1344 31334 10538 31386
rect 10590 31334 10642 31386
rect 10694 31334 10746 31386
rect 10798 31334 19862 31386
rect 19914 31334 19966 31386
rect 20018 31334 20070 31386
rect 20122 31334 29186 31386
rect 29238 31334 29290 31386
rect 29342 31334 29394 31386
rect 29446 31334 38510 31386
rect 38562 31334 38614 31386
rect 38666 31334 38718 31386
rect 38770 31334 38800 31386
rect 1344 31300 38800 31334
rect 5742 31106 5794 31118
rect 7410 31110 7422 31162
rect 7474 31110 7486 31162
rect 11660 31106 11712 31118
rect 6570 31054 6582 31106
rect 6634 31054 6646 31106
rect 8026 31054 8038 31106
rect 8090 31054 8102 31106
rect 15206 31106 15258 31118
rect 1822 30994 1874 31006
rect 1978 30998 1990 31050
rect 2042 30998 2054 31050
rect 5742 31042 5794 31054
rect 11660 31042 11712 31054
rect 14366 31050 14418 31062
rect 16270 31106 16322 31118
rect 33164 31106 33216 31118
rect 1822 30930 1874 30942
rect 2494 30994 2546 31006
rect 2494 30930 2546 30942
rect 3054 30994 3106 31006
rect 3054 30930 3106 30942
rect 6078 30994 6130 31006
rect 6078 30930 6130 30942
rect 6302 30994 6354 31006
rect 7298 30957 7310 31009
rect 7362 30957 7374 31009
rect 8318 30994 8370 31006
rect 7634 30942 7646 30994
rect 7698 30942 7710 30994
rect 6302 30930 6354 30942
rect 8318 30930 8370 30942
rect 8542 30994 8594 31006
rect 8542 30930 8594 30942
rect 10054 30994 10106 31006
rect 11902 30994 11954 31006
rect 12394 30998 12406 31050
rect 12458 30998 12470 31050
rect 10210 30942 10222 30994
rect 10274 30942 10286 30994
rect 10054 30930 10106 30942
rect 10334 30938 10386 30950
rect 2736 30882 2788 30894
rect 9662 30882 9714 30894
rect 3826 30830 3838 30882
rect 3890 30830 3902 30882
rect 11902 30930 11954 30942
rect 12574 30994 12626 31006
rect 12574 30930 12626 30942
rect 13246 30994 13298 31006
rect 13526 30994 13578 31006
rect 13346 30942 13358 30994
rect 13410 30942 13422 30994
rect 14466 30998 14478 31050
rect 14530 30998 14542 31050
rect 15206 31042 15258 31054
rect 15710 31050 15762 31062
rect 14702 31022 14754 31034
rect 14366 30986 14418 30998
rect 14702 30958 14754 30970
rect 14926 31022 14978 31034
rect 21690 31054 21702 31106
rect 21754 31054 21766 31106
rect 16270 31042 16322 31054
rect 22878 31033 22930 31045
rect 33164 31042 33216 31054
rect 15710 30986 15762 30998
rect 19518 30994 19570 31006
rect 14926 30958 14978 30970
rect 16034 30942 16046 30994
rect 16098 30942 16110 30994
rect 13246 30930 13298 30942
rect 13526 30930 13578 30942
rect 16438 30938 16490 30950
rect 16930 30942 16942 30994
rect 16994 30942 17006 30994
rect 17490 30942 17502 30994
rect 17554 30942 17566 30994
rect 17826 30942 17838 30994
rect 17890 30942 17902 30994
rect 10334 30874 10386 30886
rect 13918 30882 13970 30894
rect 2736 30818 2788 30830
rect 9662 30818 9714 30830
rect 19518 30930 19570 30942
rect 19854 30994 19906 31006
rect 19854 30930 19906 30942
rect 19966 30994 20018 31006
rect 19966 30930 20018 30942
rect 20190 30994 20242 31006
rect 20190 30930 20242 30942
rect 21198 30994 21250 31006
rect 21198 30930 21250 30942
rect 21422 30994 21474 31006
rect 21422 30930 21474 30942
rect 22318 30994 22370 31006
rect 22318 30930 22370 30942
rect 22654 30994 22706 31006
rect 23774 30994 23826 31006
rect 22878 30969 22930 30981
rect 23314 30942 23326 30994
rect 23378 30942 23390 30994
rect 22654 30930 22706 30942
rect 23774 30930 23826 30942
rect 24110 30994 24162 31006
rect 26014 30994 26066 31006
rect 29038 30994 29090 31006
rect 25442 30942 25454 30994
rect 25506 30942 25518 30994
rect 25666 30942 25678 30994
rect 25730 30942 25742 30994
rect 26786 30942 26798 30994
rect 26850 30942 26862 30994
rect 24110 30930 24162 30942
rect 26014 30930 26066 30942
rect 29038 30930 29090 30942
rect 29262 30994 29314 31006
rect 30370 30969 30382 31021
rect 30434 30969 30446 31021
rect 33406 30994 33458 31006
rect 29262 30930 29314 30942
rect 34078 30994 34130 31006
rect 33406 30930 33458 30942
rect 33910 30938 33962 30950
rect 16438 30874 16490 30886
rect 21030 30882 21082 30894
rect 13918 30818 13970 30830
rect 16774 30770 16826 30782
rect 17714 30774 17726 30826
rect 17778 30774 17790 30826
rect 21030 30818 21082 30830
rect 22990 30882 23042 30894
rect 22990 30818 23042 30830
rect 24726 30882 24778 30894
rect 34078 30930 34130 30942
rect 34302 30994 34354 31006
rect 34302 30930 34354 30942
rect 36990 30994 37042 31006
rect 36990 30930 37042 30942
rect 37326 30994 37378 31006
rect 37326 30930 37378 30942
rect 24726 30818 24778 30830
rect 25790 30826 25842 30838
rect 28690 30830 28702 30882
rect 28754 30830 28766 30882
rect 29530 30830 29542 30882
rect 29594 30830 29606 30882
rect 33910 30874 33962 30886
rect 37662 30882 37714 30894
rect 35074 30830 35086 30882
rect 35138 30830 35150 30882
rect 37662 30818 37714 30830
rect 20458 30718 20470 30770
rect 20522 30718 20534 30770
rect 25790 30762 25842 30774
rect 16774 30706 16826 30718
rect 1344 30602 38640 30636
rect 1344 30550 5876 30602
rect 5928 30550 5980 30602
rect 6032 30550 6084 30602
rect 6136 30550 15200 30602
rect 15252 30550 15304 30602
rect 15356 30550 15408 30602
rect 15460 30550 24524 30602
rect 24576 30550 24628 30602
rect 24680 30550 24732 30602
rect 24784 30550 33848 30602
rect 33900 30550 33952 30602
rect 34004 30550 34056 30602
rect 34108 30550 38640 30602
rect 1344 30516 38640 30550
rect 3726 30434 3778 30446
rect 3726 30370 3778 30382
rect 8262 30434 8314 30446
rect 8262 30370 8314 30382
rect 12798 30434 12850 30446
rect 17950 30434 18002 30446
rect 12798 30370 12850 30382
rect 13526 30378 13578 30390
rect 9550 30322 9602 30334
rect 17950 30370 18002 30382
rect 22150 30434 22202 30446
rect 22150 30370 22202 30382
rect 31726 30434 31778 30446
rect 31726 30370 31778 30382
rect 13526 30314 13578 30326
rect 14944 30322 14996 30334
rect 9550 30258 9602 30270
rect 14198 30266 14250 30278
rect 1878 30210 1930 30222
rect 1878 30146 1930 30158
rect 2382 30210 2434 30222
rect 2382 30146 2434 30158
rect 2624 30210 2676 30222
rect 2624 30146 2676 30158
rect 4846 30210 4898 30222
rect 4846 30146 4898 30158
rect 6134 30210 6186 30222
rect 6134 30146 6186 30158
rect 6862 30210 6914 30222
rect 6862 30146 6914 30158
rect 7534 30210 7586 30222
rect 1710 30098 1762 30110
rect 7018 30102 7030 30154
rect 7082 30102 7094 30154
rect 7534 30146 7586 30158
rect 7776 30210 7828 30222
rect 10222 30210 10274 30222
rect 7776 30146 7828 30158
rect 8990 30182 9042 30194
rect 8530 30102 8542 30154
rect 8594 30102 8606 30154
rect 8754 30102 8766 30154
rect 8818 30102 8830 30154
rect 8990 30118 9042 30130
rect 9102 30154 9154 30166
rect 10098 30158 10110 30210
rect 10162 30158 10174 30210
rect 9932 30102 9944 30154
rect 9996 30102 10008 30154
rect 10222 30146 10274 30158
rect 10446 30210 10498 30222
rect 14944 30258 14996 30270
rect 17110 30322 17162 30334
rect 17110 30258 17162 30270
rect 36038 30322 36090 30334
rect 36038 30258 36090 30270
rect 10446 30146 10498 30158
rect 12126 30154 12178 30166
rect 12226 30158 12238 30210
rect 12290 30158 12302 30210
rect 13682 30158 13694 30210
rect 13746 30158 13758 30210
rect 14198 30202 14250 30214
rect 14702 30210 14754 30222
rect 12394 30102 12406 30154
rect 12458 30102 12470 30154
rect 14702 30146 14754 30158
rect 15542 30210 15594 30222
rect 15542 30146 15594 30158
rect 16046 30210 16098 30222
rect 16046 30146 16098 30158
rect 16288 30210 16340 30222
rect 16288 30146 16340 30158
rect 17614 30210 17666 30222
rect 17614 30146 17666 30158
rect 19630 30210 19682 30222
rect 19630 30146 19682 30158
rect 20190 30210 20242 30222
rect 20190 30146 20242 30158
rect 20302 30210 20354 30222
rect 20302 30146 20354 30158
rect 21310 30210 21362 30222
rect 21310 30146 21362 30158
rect 21422 30210 21474 30222
rect 22430 30210 22482 30222
rect 22878 30210 22930 30222
rect 21690 30158 21702 30210
rect 21754 30158 21766 30210
rect 22530 30158 22542 30210
rect 22594 30158 22606 30210
rect 21422 30146 21474 30158
rect 22430 30146 22482 30158
rect 9102 30090 9154 30102
rect 12126 30090 12178 30102
rect 14030 30098 14082 30110
rect 1710 30034 1762 30046
rect 14030 30034 14082 30046
rect 15374 30098 15426 30110
rect 22698 30102 22710 30154
rect 22762 30102 22774 30154
rect 22878 30146 22930 30158
rect 23774 30210 23826 30222
rect 26462 30210 26514 30222
rect 24546 30158 24558 30210
rect 24610 30158 24622 30210
rect 23774 30146 23826 30158
rect 26462 30146 26514 30158
rect 27078 30210 27130 30222
rect 27078 30146 27130 30158
rect 27694 30210 27746 30222
rect 27694 30146 27746 30158
rect 28030 30210 28082 30222
rect 28030 30146 28082 30158
rect 28142 30210 28194 30222
rect 28142 30146 28194 30158
rect 29486 30210 29538 30222
rect 29486 30146 29538 30158
rect 29598 30210 29650 30222
rect 37158 30210 37210 30222
rect 29866 30158 29878 30210
rect 29930 30158 29942 30210
rect 29598 30146 29650 30158
rect 32386 30130 32398 30182
rect 32450 30130 32462 30182
rect 35298 30130 35310 30182
rect 35362 30130 35374 30182
rect 37158 30146 37210 30158
rect 37662 30210 37714 30222
rect 37662 30146 37714 30158
rect 36990 30098 37042 30110
rect 19898 30046 19910 30098
rect 19962 30046 19974 30098
rect 15374 30034 15426 30046
rect 36990 30034 37042 30046
rect 37904 30098 37956 30110
rect 37904 30034 37956 30046
rect 10782 29986 10834 29998
rect 10782 29922 10834 29934
rect 11398 29986 11450 29998
rect 11398 29922 11450 29934
rect 11846 29986 11898 29998
rect 11846 29922 11898 29934
rect 19294 29986 19346 29998
rect 19294 29922 19346 29934
rect 28478 29986 28530 29998
rect 28478 29922 28530 29934
rect 34190 29986 34242 29998
rect 34190 29922 34242 29934
rect 1344 29818 38800 29852
rect 1344 29766 10538 29818
rect 10590 29766 10642 29818
rect 10694 29766 10746 29818
rect 10798 29766 19862 29818
rect 19914 29766 19966 29818
rect 20018 29766 20070 29818
rect 20122 29766 29186 29818
rect 29238 29766 29290 29818
rect 29342 29766 29394 29818
rect 29446 29766 38510 29818
rect 38562 29766 38614 29818
rect 38666 29766 38718 29818
rect 38770 29766 38800 29818
rect 1344 29732 38800 29766
rect 11230 29650 11282 29662
rect 11230 29586 11282 29598
rect 12126 29650 12178 29662
rect 12126 29586 12178 29598
rect 14534 29650 14586 29662
rect 14534 29586 14586 29598
rect 23774 29650 23826 29662
rect 13936 29538 13988 29550
rect 14914 29542 14926 29594
rect 14978 29542 14990 29594
rect 23774 29586 23826 29598
rect 29094 29650 29146 29662
rect 29094 29586 29146 29598
rect 33238 29650 33290 29662
rect 33238 29586 33290 29598
rect 8138 29486 8150 29538
rect 8202 29486 8214 29538
rect 2494 29426 2546 29438
rect 2494 29362 2546 29374
rect 4958 29426 5010 29438
rect 5450 29430 5462 29482
rect 5514 29430 5526 29482
rect 4958 29362 5010 29374
rect 5630 29426 5682 29438
rect 7298 29389 7310 29441
rect 7362 29389 7374 29441
rect 8430 29426 8482 29438
rect 7634 29374 7646 29426
rect 7698 29374 7710 29426
rect 5630 29362 5682 29374
rect 8430 29362 8482 29374
rect 8654 29426 8706 29438
rect 10782 29426 10834 29438
rect 9538 29374 9550 29426
rect 9602 29374 9614 29426
rect 9874 29374 9886 29426
rect 9938 29374 9950 29426
rect 8654 29362 8706 29374
rect 10782 29362 10834 29374
rect 10894 29426 10946 29438
rect 10894 29362 10946 29374
rect 12462 29426 12514 29438
rect 12462 29362 12514 29374
rect 13022 29426 13074 29438
rect 13178 29430 13190 29482
rect 13242 29430 13254 29482
rect 13936 29474 13988 29486
rect 19910 29538 19962 29550
rect 13022 29362 13074 29374
rect 13694 29426 13746 29438
rect 13694 29362 13746 29374
rect 15038 29426 15090 29438
rect 15250 29430 15262 29482
rect 15314 29430 15326 29482
rect 19182 29426 19234 29438
rect 19338 29430 19350 29482
rect 19402 29430 19414 29482
rect 19910 29474 19962 29486
rect 25510 29538 25562 29550
rect 32062 29538 32114 29550
rect 19630 29426 19682 29438
rect 15586 29374 15598 29426
rect 15650 29374 15662 29426
rect 19506 29374 19518 29426
rect 19570 29374 19582 29426
rect 15038 29362 15090 29374
rect 19182 29362 19234 29374
rect 19630 29362 19682 29374
rect 20526 29426 20578 29438
rect 20738 29430 20750 29482
rect 20802 29430 20814 29482
rect 25510 29474 25562 29486
rect 29262 29482 29314 29494
rect 22318 29426 22370 29438
rect 23438 29426 23490 29438
rect 21186 29374 21198 29426
rect 21250 29374 21262 29426
rect 21634 29374 21646 29426
rect 21698 29374 21710 29426
rect 22866 29374 22878 29426
rect 22930 29374 22942 29426
rect 26114 29401 26126 29453
rect 26178 29401 26190 29453
rect 32062 29474 32114 29486
rect 29262 29418 29314 29430
rect 29374 29426 29426 29438
rect 20526 29362 20578 29374
rect 22318 29362 22370 29374
rect 23438 29362 23490 29374
rect 33842 29374 33854 29426
rect 33906 29374 33918 29426
rect 36082 29401 36094 29453
rect 36146 29401 36158 29453
rect 38222 29426 38274 29438
rect 29374 29362 29426 29374
rect 38222 29362 38274 29374
rect 17558 29314 17610 29326
rect 7186 29262 7198 29314
rect 7250 29262 7262 29314
rect 3614 29202 3666 29214
rect 3614 29138 3666 29150
rect 4716 29202 4768 29214
rect 9650 29206 9662 29258
rect 9714 29206 9726 29258
rect 17558 29250 17610 29262
rect 18230 29314 18282 29326
rect 18230 29250 18282 29262
rect 18678 29314 18730 29326
rect 18678 29250 18730 29262
rect 20862 29314 20914 29326
rect 24726 29314 24778 29326
rect 20862 29250 20914 29262
rect 22710 29258 22762 29270
rect 4716 29138 4768 29150
rect 10446 29202 10498 29214
rect 21522 29206 21534 29258
rect 21586 29206 21598 29258
rect 24726 29250 24778 29262
rect 28758 29314 28810 29326
rect 30146 29262 30158 29314
rect 30210 29262 30222 29314
rect 28758 29250 28810 29262
rect 22710 29194 22762 29206
rect 26798 29202 26850 29214
rect 10446 29138 10498 29150
rect 26798 29138 26850 29150
rect 36766 29202 36818 29214
rect 36766 29138 36818 29150
rect 1344 29034 38640 29068
rect 1344 28982 5876 29034
rect 5928 28982 5980 29034
rect 6032 28982 6084 29034
rect 6136 28982 15200 29034
rect 15252 28982 15304 29034
rect 15356 28982 15408 29034
rect 15460 28982 24524 29034
rect 24576 28982 24628 29034
rect 24680 28982 24732 29034
rect 24784 28982 33848 29034
rect 33900 28982 33952 29034
rect 34004 28982 34056 29034
rect 34108 28982 38640 29034
rect 1344 28948 38640 28982
rect 7086 28866 7138 28878
rect 7086 28802 7138 28814
rect 8374 28866 8426 28878
rect 8374 28802 8426 28814
rect 11342 28866 11394 28878
rect 11342 28802 11394 28814
rect 12126 28866 12178 28878
rect 12126 28802 12178 28814
rect 16886 28866 16938 28878
rect 16886 28802 16938 28814
rect 19872 28866 19924 28878
rect 19872 28802 19924 28814
rect 22262 28866 22314 28878
rect 5798 28754 5850 28766
rect 3042 28702 3054 28754
rect 3106 28702 3118 28754
rect 4946 28702 4958 28754
rect 5010 28702 5022 28754
rect 5798 28690 5850 28702
rect 6582 28754 6634 28766
rect 6582 28690 6634 28702
rect 10222 28754 10274 28766
rect 10222 28690 10274 28702
rect 12742 28754 12794 28766
rect 12742 28690 12794 28702
rect 13638 28754 13690 28766
rect 17390 28754 17442 28766
rect 20514 28758 20526 28810
rect 20578 28758 20590 28810
rect 22262 28802 22314 28814
rect 25454 28866 25506 28878
rect 25454 28802 25506 28814
rect 30960 28866 31012 28878
rect 30960 28802 31012 28814
rect 34750 28866 34802 28878
rect 34750 28802 34802 28814
rect 13638 28690 13690 28702
rect 16326 28698 16378 28710
rect 2270 28642 2322 28654
rect 2270 28578 2322 28590
rect 6750 28642 6802 28654
rect 11678 28642 11730 28654
rect 6750 28578 6802 28590
rect 7634 28575 7646 28627
rect 7698 28575 7710 28627
rect 7970 28590 7982 28642
rect 8034 28590 8046 28642
rect 8654 28614 8706 28626
rect 8654 28550 8706 28562
rect 8878 28614 8930 28626
rect 9214 28607 9266 28619
rect 8878 28550 8930 28562
rect 9046 28586 9098 28598
rect 9214 28543 9266 28555
rect 10054 28586 10106 28598
rect 10434 28590 10446 28642
rect 10498 28590 10510 28642
rect 9046 28522 9098 28534
rect 10054 28522 10106 28534
rect 10782 28586 10834 28598
rect 11678 28578 11730 28590
rect 11790 28642 11842 28654
rect 11790 28578 11842 28590
rect 16158 28642 16210 28654
rect 22766 28754 22818 28766
rect 17390 28690 17442 28702
rect 19126 28698 19178 28710
rect 16326 28634 16378 28646
rect 16606 28642 16658 28654
rect 18062 28642 18114 28654
rect 21702 28698 21754 28710
rect 16158 28578 16210 28590
rect 17938 28590 17950 28642
rect 18002 28590 18014 28642
rect 18722 28590 18734 28642
rect 18786 28590 18798 28642
rect 19126 28634 19178 28646
rect 19630 28642 19682 28654
rect 21534 28642 21586 28654
rect 20402 28590 20414 28642
rect 20466 28590 20478 28642
rect 20626 28590 20638 28642
rect 20690 28590 20702 28642
rect 22766 28690 22818 28702
rect 24502 28754 24554 28766
rect 28466 28702 28478 28754
rect 28530 28702 28542 28754
rect 24502 28690 24554 28702
rect 37158 28698 37210 28710
rect 21702 28634 21754 28646
rect 21982 28642 22034 28654
rect 16606 28578 16658 28590
rect 10782 28522 10834 28534
rect 16494 28530 16546 28542
rect 17772 28534 17784 28586
rect 17836 28534 17848 28586
rect 18062 28578 18114 28590
rect 19630 28578 19682 28590
rect 21534 28578 21586 28590
rect 21982 28578 22034 28590
rect 23102 28642 23154 28654
rect 23102 28578 23154 28590
rect 24782 28642 24834 28654
rect 25060 28642 25112 28654
rect 24882 28590 24894 28642
rect 24946 28590 24958 28642
rect 24782 28578 24834 28590
rect 25060 28578 25112 28590
rect 25790 28642 25842 28654
rect 29262 28642 29314 28654
rect 26562 28590 26574 28642
rect 26626 28590 26638 28642
rect 25790 28578 25842 28590
rect 29262 28578 29314 28590
rect 29598 28642 29650 28654
rect 29598 28578 29650 28590
rect 30214 28642 30266 28654
rect 30214 28578 30266 28590
rect 30718 28642 30770 28654
rect 30718 28578 30770 28590
rect 32062 28642 32114 28654
rect 7646 28474 7698 28486
rect 16494 28466 16546 28478
rect 18958 28530 19010 28542
rect 18958 28466 19010 28478
rect 21870 28530 21922 28542
rect 21870 28466 21922 28478
rect 31390 28530 31442 28542
rect 31546 28534 31558 28586
rect 31610 28534 31622 28586
rect 32062 28578 32114 28590
rect 32846 28642 32898 28654
rect 32846 28578 32898 28590
rect 33070 28642 33122 28654
rect 37158 28634 37210 28646
rect 37662 28642 37714 28654
rect 33070 28578 33122 28590
rect 36418 28562 36430 28614
rect 36482 28562 36494 28614
rect 37662 28578 37714 28590
rect 7646 28410 7698 28422
rect 18566 28418 18618 28430
rect 18566 28354 18618 28366
rect 23494 28418 23546 28430
rect 30258 28422 30270 28474
rect 30322 28422 30334 28474
rect 31390 28466 31442 28478
rect 32304 28530 32356 28542
rect 36990 28530 37042 28542
rect 33338 28478 33350 28530
rect 33402 28478 33414 28530
rect 32304 28466 32356 28478
rect 36990 28466 37042 28478
rect 37904 28530 37956 28542
rect 37904 28466 37956 28478
rect 23494 28354 23546 28366
rect 1344 28250 38800 28284
rect 1344 28198 10538 28250
rect 10590 28198 10642 28250
rect 10694 28198 10746 28250
rect 10798 28198 19862 28250
rect 19914 28198 19966 28250
rect 20018 28198 20070 28250
rect 20122 28198 29186 28250
rect 29238 28198 29290 28250
rect 29342 28198 29394 28250
rect 29446 28198 38510 28250
rect 38562 28198 38614 28250
rect 38666 28198 38718 28250
rect 38770 28198 38800 28250
rect 1344 28164 38800 28198
rect 9718 28082 9770 28094
rect 9718 28018 9770 28030
rect 13022 28082 13074 28094
rect 13022 28018 13074 28030
rect 14814 28082 14866 28094
rect 14814 28018 14866 28030
rect 18286 28082 18338 28094
rect 18286 28018 18338 28030
rect 22150 28082 22202 28094
rect 22150 28018 22202 28030
rect 28142 28082 28194 28094
rect 7646 27970 7698 27982
rect 2986 27918 2998 27970
rect 3050 27918 3062 27970
rect 7646 27906 7698 27918
rect 8560 27970 8612 27982
rect 3278 27858 3330 27870
rect 3278 27794 3330 27806
rect 3502 27858 3554 27870
rect 3502 27794 3554 27806
rect 4398 27858 4450 27870
rect 7802 27862 7814 27914
rect 7866 27862 7878 27914
rect 8560 27906 8612 27918
rect 10166 27970 10218 27982
rect 10166 27906 10218 27918
rect 10558 27970 10610 27982
rect 24658 27974 24670 28026
rect 24722 27974 24734 28026
rect 28142 28018 28194 28030
rect 29206 28082 29258 28094
rect 29206 28018 29258 28030
rect 30046 28082 30098 28094
rect 30046 28018 30098 28030
rect 27134 27970 27186 27982
rect 37438 27970 37490 27982
rect 16426 27918 16438 27970
rect 16490 27918 16502 27970
rect 30986 27918 30998 27970
rect 31050 27918 31062 27970
rect 10558 27906 10610 27918
rect 20336 27895 20388 27907
rect 4398 27794 4450 27806
rect 8318 27858 8370 27870
rect 10446 27858 10498 27870
rect 9818 27806 9830 27858
rect 9882 27806 9894 27858
rect 8318 27794 8370 27806
rect 10446 27794 10498 27806
rect 10726 27858 10778 27870
rect 10726 27794 10778 27806
rect 10894 27858 10946 27870
rect 10894 27794 10946 27806
rect 11230 27858 11282 27870
rect 11510 27858 11562 27870
rect 11330 27806 11342 27858
rect 11394 27806 11406 27858
rect 11230 27794 11282 27806
rect 11510 27794 11562 27806
rect 14142 27858 14194 27870
rect 14142 27794 14194 27806
rect 15150 27858 15202 27870
rect 15150 27794 15202 27806
rect 16718 27858 16770 27870
rect 16718 27794 16770 27806
rect 16830 27858 16882 27870
rect 16830 27794 16882 27806
rect 17838 27858 17890 27870
rect 17838 27794 17890 27806
rect 17950 27858 18002 27870
rect 17950 27794 18002 27806
rect 18734 27858 18786 27870
rect 19012 27858 19064 27870
rect 18834 27806 18846 27858
rect 18898 27806 18910 27858
rect 18734 27794 18786 27806
rect 19012 27794 19064 27806
rect 20078 27858 20130 27870
rect 20178 27806 20190 27858
rect 20242 27806 20254 27858
rect 23886 27858 23938 27870
rect 25342 27858 25394 27870
rect 25573 27862 25585 27914
rect 25637 27862 25649 27914
rect 20336 27831 20388 27843
rect 21186 27806 21198 27858
rect 21250 27806 21262 27858
rect 21522 27806 21534 27858
rect 21586 27806 21598 27858
rect 24546 27806 24558 27858
rect 24610 27806 24622 27858
rect 20078 27794 20130 27806
rect 23886 27794 23938 27806
rect 25342 27794 25394 27806
rect 26462 27858 26514 27870
rect 26462 27794 26514 27806
rect 26798 27858 26850 27870
rect 26954 27862 26966 27914
rect 27018 27862 27030 27914
rect 27134 27906 27186 27918
rect 26798 27794 26850 27806
rect 27246 27858 27298 27870
rect 27246 27794 27298 27806
rect 27526 27858 27578 27870
rect 27526 27794 27578 27806
rect 27806 27858 27858 27870
rect 30382 27858 30434 27870
rect 28802 27806 28814 27858
rect 28866 27806 28878 27858
rect 27806 27794 27858 27806
rect 30382 27794 30434 27806
rect 30494 27858 30546 27870
rect 30494 27794 30546 27806
rect 30718 27858 30770 27870
rect 30718 27794 30770 27806
rect 31502 27858 31554 27870
rect 31502 27794 31554 27806
rect 31670 27858 31722 27870
rect 31670 27794 31722 27806
rect 32174 27858 32226 27870
rect 32174 27794 32226 27806
rect 32416 27858 32468 27870
rect 32416 27794 32468 27806
rect 33070 27858 33122 27870
rect 33226 27862 33238 27914
rect 33290 27862 33302 27914
rect 37438 27906 37490 27918
rect 33070 27794 33122 27806
rect 33742 27858 33794 27870
rect 33742 27794 33794 27806
rect 34750 27858 34802 27870
rect 34750 27794 34802 27806
rect 38334 27858 38386 27870
rect 38334 27794 38386 27806
rect 11902 27746 11954 27758
rect 11902 27682 11954 27694
rect 19406 27746 19458 27758
rect 19406 27682 19458 27694
rect 20750 27746 20802 27758
rect 29654 27746 29706 27758
rect 20750 27682 20802 27694
rect 21646 27690 21698 27702
rect 5518 27634 5570 27646
rect 5518 27570 5570 27582
rect 17502 27634 17554 27646
rect 21646 27626 21698 27638
rect 28646 27690 28698 27702
rect 35522 27694 35534 27746
rect 35586 27694 35598 27746
rect 29654 27682 29706 27694
rect 28646 27626 28698 27638
rect 33984 27634 34036 27646
rect 17502 27570 17554 27582
rect 33984 27570 34036 27582
rect 37998 27634 38050 27646
rect 37998 27570 38050 27582
rect 1344 27466 38640 27500
rect 1344 27414 5876 27466
rect 5928 27414 5980 27466
rect 6032 27414 6084 27466
rect 6136 27414 15200 27466
rect 15252 27414 15304 27466
rect 15356 27414 15408 27466
rect 15460 27414 24524 27466
rect 24576 27414 24628 27466
rect 24680 27414 24732 27466
rect 24784 27414 33848 27466
rect 33900 27414 33952 27466
rect 34004 27414 34056 27466
rect 34108 27414 38640 27466
rect 1344 27380 38640 27414
rect 8206 27298 8258 27310
rect 8206 27234 8258 27246
rect 14012 27298 14064 27310
rect 14012 27234 14064 27246
rect 17726 27298 17778 27310
rect 24446 27298 24498 27310
rect 30494 27298 30546 27310
rect 34750 27298 34802 27310
rect 18554 27246 18566 27298
rect 18618 27246 18630 27298
rect 17726 27234 17778 27246
rect 21310 27242 21362 27254
rect 4230 27186 4282 27198
rect 12854 27186 12906 27198
rect 9874 27134 9886 27186
rect 9938 27134 9950 27186
rect 11778 27134 11790 27186
rect 11842 27134 11854 27186
rect 4230 27122 4282 27134
rect 12854 27122 12906 27134
rect 13638 27186 13690 27198
rect 19966 27186 20018 27198
rect 13638 27122 13690 27134
rect 14758 27130 14810 27142
rect 8598 27074 8650 27086
rect 8878 27074 8930 27086
rect 8754 27022 8766 27074
rect 8818 27022 8830 27074
rect 8598 27010 8650 27022
rect 8878 27010 8930 27022
rect 9102 27074 9154 27086
rect 14254 27074 14306 27086
rect 12114 27022 12126 27074
rect 12178 27022 12190 27074
rect 26954 27246 26966 27298
rect 27018 27246 27030 27298
rect 32666 27246 32678 27298
rect 32730 27246 32742 27298
rect 24446 27234 24498 27246
rect 30494 27234 30546 27246
rect 34750 27234 34802 27246
rect 21310 27178 21362 27190
rect 27862 27186 27914 27198
rect 19966 27122 20018 27134
rect 27862 27122 27914 27134
rect 29318 27186 29370 27198
rect 29318 27122 29370 27134
rect 31614 27186 31666 27198
rect 31614 27122 31666 27134
rect 37830 27130 37882 27142
rect 14758 27066 14810 27078
rect 15262 27074 15314 27086
rect 9102 27010 9154 27022
rect 14254 27010 14306 27022
rect 15262 27010 15314 27022
rect 15430 27074 15482 27086
rect 15430 27010 15482 27022
rect 15934 27074 15986 27086
rect 15934 27010 15986 27022
rect 16176 27074 16228 27086
rect 16176 27010 16228 27022
rect 17390 27074 17442 27086
rect 17390 27010 17442 27022
rect 18846 27074 18898 27086
rect 18846 27010 18898 27022
rect 19070 27074 19122 27086
rect 19070 27010 19122 27022
rect 19294 27074 19346 27086
rect 19572 27074 19624 27086
rect 19394 27022 19406 27074
rect 19458 27022 19470 27074
rect 19294 27010 19346 27022
rect 19572 27010 19624 27022
rect 20806 27074 20858 27086
rect 23774 27074 23826 27086
rect 24052 27074 24104 27086
rect 21410 27022 21422 27074
rect 21474 27022 21486 27074
rect 21634 27022 21646 27074
rect 21698 27022 21710 27074
rect 23874 27022 23886 27074
rect 23938 27022 23950 27074
rect 20806 27010 20858 27022
rect 23774 27010 23826 27022
rect 24052 27010 24104 27022
rect 25118 27074 25170 27086
rect 26014 27074 26066 27086
rect 25666 27022 25678 27074
rect 25730 27022 25742 27074
rect 25118 27010 25170 27022
rect 14926 26962 14978 26974
rect 25330 26966 25342 27018
rect 25394 26966 25406 27018
rect 26014 27010 26066 27022
rect 26238 27074 26290 27086
rect 27246 27074 27298 27086
rect 26506 27022 26518 27074
rect 26570 27022 26582 27074
rect 26238 27010 26290 27022
rect 27246 27010 27298 27022
rect 27358 27074 27410 27086
rect 27358 27010 27410 27022
rect 30830 27074 30882 27086
rect 30830 27010 30882 27022
rect 31278 27074 31330 27086
rect 32286 27074 32338 27086
rect 31938 27022 31950 27074
rect 32002 27022 32014 27074
rect 31278 27010 31330 27022
rect 31490 26966 31502 27018
rect 31554 26966 31566 27018
rect 32286 27010 32338 27022
rect 32398 27074 32450 27086
rect 36486 27074 36538 27086
rect 32398 27010 32450 27022
rect 33394 26994 33406 27046
rect 33458 26994 33470 27046
rect 36486 27010 36538 27022
rect 37326 27074 37378 27086
rect 37830 27066 37882 27078
rect 37326 27010 37378 27022
rect 14926 26898 14978 26910
rect 37084 26962 37136 26974
rect 25218 26854 25230 26906
rect 25282 26854 25294 26906
rect 37084 26898 37136 26910
rect 37998 26962 38050 26974
rect 37998 26898 38050 26910
rect 28310 26850 28362 26862
rect 28310 26786 28362 26798
rect 1344 26682 38800 26716
rect 1344 26630 10538 26682
rect 10590 26630 10642 26682
rect 10694 26630 10746 26682
rect 10798 26630 19862 26682
rect 19914 26630 19966 26682
rect 20018 26630 20070 26682
rect 20122 26630 29186 26682
rect 29238 26630 29290 26682
rect 29342 26630 29394 26682
rect 29446 26630 38510 26682
rect 38562 26630 38614 26682
rect 38666 26630 38718 26682
rect 38770 26630 38800 26682
rect 1344 26596 38800 26630
rect 11286 26514 11338 26526
rect 11286 26450 11338 26462
rect 13358 26514 13410 26526
rect 13358 26450 13410 26462
rect 16718 26514 16770 26526
rect 16718 26450 16770 26462
rect 26574 26514 26626 26526
rect 7198 26402 7250 26414
rect 2942 26290 2994 26302
rect 3098 26294 3110 26346
rect 3162 26294 3174 26346
rect 7198 26338 7250 26350
rect 20320 26402 20372 26414
rect 21186 26406 21198 26458
rect 21250 26406 21262 26458
rect 26574 26450 26626 26462
rect 27190 26514 27242 26526
rect 27190 26450 27242 26462
rect 33238 26514 33290 26526
rect 33238 26450 33290 26462
rect 35086 26514 35138 26526
rect 35086 26450 35138 26462
rect 2942 26226 2994 26238
rect 3614 26290 3666 26302
rect 3614 26226 3666 26238
rect 4510 26290 4562 26302
rect 5282 26238 5294 26290
rect 5346 26238 5358 26290
rect 10434 26238 10446 26290
rect 10498 26238 10510 26290
rect 10658 26238 10670 26290
rect 10722 26238 10734 26290
rect 12338 26265 12350 26317
rect 12402 26265 12414 26317
rect 16382 26290 16434 26302
rect 4510 26226 4562 26238
rect 16382 26226 16434 26238
rect 17278 26290 17330 26302
rect 17278 26226 17330 26238
rect 19406 26290 19458 26302
rect 19562 26294 19574 26346
rect 19626 26294 19638 26346
rect 20320 26338 20372 26350
rect 25958 26402 26010 26414
rect 30314 26350 30326 26402
rect 30378 26350 30390 26402
rect 25958 26338 26010 26350
rect 21030 26319 21082 26331
rect 19406 26226 19458 26238
rect 20078 26290 20130 26302
rect 24222 26290 24274 26302
rect 21030 26255 21082 26267
rect 21298 26238 21310 26290
rect 21362 26238 21374 26290
rect 20078 26226 20130 26238
rect 24222 26226 24274 26238
rect 25230 26290 25282 26302
rect 25678 26290 25730 26302
rect 25230 26226 25282 26238
rect 25398 26234 25450 26246
rect 25554 26238 25566 26290
rect 25618 26238 25630 26290
rect 7814 26178 7866 26190
rect 14982 26178 15034 26190
rect 7814 26114 7866 26126
rect 10334 26122 10386 26134
rect 3856 26066 3908 26078
rect 14982 26114 15034 26126
rect 24558 26178 24610 26190
rect 25678 26226 25730 26238
rect 26238 26290 26290 26302
rect 26238 26226 26290 26238
rect 28198 26290 28250 26302
rect 28198 26226 28250 26238
rect 30606 26290 30658 26302
rect 30606 26226 30658 26238
rect 30718 26290 30770 26302
rect 31042 26238 31054 26290
rect 31106 26238 31118 26290
rect 31378 26265 31390 26317
rect 31442 26265 31454 26317
rect 31726 26290 31778 26302
rect 30718 26226 30770 26238
rect 31726 26226 31778 26238
rect 33630 26290 33682 26302
rect 35746 26265 35758 26317
rect 35810 26265 35822 26317
rect 33630 26226 33682 26238
rect 25398 26170 25450 26182
rect 31154 26126 31166 26178
rect 31218 26126 31230 26178
rect 36754 26126 36766 26178
rect 36818 26126 36830 26178
rect 24558 26114 24610 26126
rect 10334 26058 10386 26070
rect 17614 26066 17666 26078
rect 3856 26002 3908 26014
rect 17614 26002 17666 26014
rect 1344 25898 38640 25932
rect 1344 25846 5876 25898
rect 5928 25846 5980 25898
rect 6032 25846 6084 25898
rect 6136 25846 15200 25898
rect 15252 25846 15304 25898
rect 15356 25846 15408 25898
rect 15460 25846 24524 25898
rect 24576 25846 24628 25898
rect 24680 25846 24732 25898
rect 24784 25846 33848 25898
rect 33900 25846 33952 25898
rect 34004 25846 34056 25898
rect 34108 25846 38640 25898
rect 1344 25812 38640 25846
rect 10726 25730 10778 25742
rect 4666 25678 4678 25730
rect 4730 25678 4742 25730
rect 10726 25666 10778 25678
rect 13806 25730 13858 25742
rect 20078 25730 20130 25742
rect 13806 25666 13858 25678
rect 15934 25674 15986 25686
rect 10166 25618 10218 25630
rect 20078 25666 20130 25678
rect 20694 25730 20746 25742
rect 25162 25678 25174 25730
rect 25226 25678 25238 25730
rect 20694 25666 20746 25678
rect 15934 25610 15986 25622
rect 18958 25618 19010 25630
rect 10166 25554 10218 25566
rect 32946 25566 32958 25618
rect 33010 25566 33022 25618
rect 18958 25554 19010 25566
rect 37830 25562 37882 25574
rect 3950 25506 4002 25518
rect 3950 25442 4002 25454
rect 4958 25506 5010 25518
rect 4958 25442 5010 25454
rect 5182 25506 5234 25518
rect 5182 25442 5234 25454
rect 5948 25506 6000 25518
rect 5948 25442 6000 25454
rect 6190 25506 6242 25518
rect 6190 25442 6242 25454
rect 6694 25506 6746 25518
rect 11006 25506 11058 25518
rect 15262 25506 15314 25518
rect 19352 25506 19404 25518
rect 19630 25506 19682 25518
rect 7410 25454 7422 25506
rect 7474 25454 7486 25506
rect 6694 25442 6746 25454
rect 9650 25426 9662 25478
rect 9714 25426 9726 25478
rect 10546 25454 10558 25506
rect 10610 25454 10622 25506
rect 12450 25454 12462 25506
rect 12514 25454 12526 25506
rect 15474 25454 15486 25506
rect 15538 25454 15550 25506
rect 15810 25454 15822 25506
rect 15874 25454 15886 25506
rect 18610 25454 18622 25506
rect 18674 25454 18686 25506
rect 19506 25454 19518 25506
rect 19570 25454 19582 25506
rect 11006 25442 11058 25454
rect 15262 25442 15314 25454
rect 19352 25442 19404 25454
rect 19630 25442 19682 25454
rect 20414 25506 20466 25518
rect 24782 25506 24834 25518
rect 20514 25454 20526 25506
rect 20578 25454 20590 25506
rect 24210 25454 24222 25506
rect 24274 25454 24286 25506
rect 20414 25442 20466 25454
rect 24782 25442 24834 25454
rect 25454 25506 25506 25518
rect 25454 25442 25506 25454
rect 25678 25506 25730 25518
rect 25678 25442 25730 25454
rect 26070 25506 26122 25518
rect 28366 25506 28418 25518
rect 30494 25506 30546 25518
rect 27682 25454 27694 25506
rect 27746 25454 27758 25506
rect 29586 25454 29598 25506
rect 29650 25454 29662 25506
rect 29922 25454 29934 25506
rect 29986 25454 29998 25506
rect 26070 25442 26122 25454
rect 28366 25442 28418 25454
rect 30258 25398 30270 25450
rect 30322 25398 30334 25450
rect 30494 25442 30546 25454
rect 31278 25506 31330 25518
rect 32510 25506 32562 25518
rect 34190 25506 34242 25518
rect 37326 25506 37378 25518
rect 31938 25454 31950 25506
rect 32002 25454 32014 25506
rect 33170 25454 33182 25506
rect 33234 25454 33246 25506
rect 33506 25454 33518 25506
rect 33570 25454 33582 25506
rect 31278 25442 31330 25454
rect 31490 25398 31502 25450
rect 31554 25398 31566 25450
rect 32510 25442 32562 25454
rect 32722 25398 32734 25450
rect 32786 25398 32798 25450
rect 33842 25398 33854 25450
rect 33906 25398 33918 25450
rect 34190 25442 34242 25454
rect 35366 25450 35418 25462
rect 35746 25454 35758 25506
rect 35810 25454 35822 25506
rect 37830 25498 37882 25510
rect 35366 25386 35418 25398
rect 35534 25394 35586 25406
rect 35970 25398 35982 25450
rect 36034 25398 36046 25450
rect 37326 25442 37378 25454
rect 29430 25338 29482 25350
rect 2830 25282 2882 25294
rect 2830 25218 2882 25230
rect 4342 25282 4394 25294
rect 6626 25286 6638 25338
rect 6690 25286 6702 25338
rect 4342 25218 4394 25230
rect 18118 25282 18170 25294
rect 18118 25218 18170 25230
rect 18454 25282 18506 25294
rect 18454 25218 18506 25230
rect 21478 25282 21530 25294
rect 24098 25286 24110 25338
rect 24162 25286 24174 25338
rect 21478 25218 21530 25230
rect 26518 25282 26570 25294
rect 27906 25286 27918 25338
rect 27970 25286 27982 25338
rect 30594 25286 30606 25338
rect 30658 25286 30670 25338
rect 31826 25286 31838 25338
rect 31890 25286 31902 25338
rect 33618 25286 33630 25338
rect 33682 25286 33694 25338
rect 35534 25330 35586 25342
rect 37084 25394 37136 25406
rect 37084 25330 37136 25342
rect 37998 25394 38050 25406
rect 37998 25330 38050 25342
rect 29430 25274 29482 25286
rect 26518 25218 26570 25230
rect 1344 25114 38800 25148
rect 1344 25062 10538 25114
rect 10590 25062 10642 25114
rect 10694 25062 10746 25114
rect 10798 25062 19862 25114
rect 19914 25062 19966 25114
rect 20018 25062 20070 25114
rect 20122 25062 29186 25114
rect 29238 25062 29290 25114
rect 29342 25062 29394 25114
rect 29446 25062 38510 25114
rect 38562 25062 38614 25114
rect 38666 25062 38718 25114
rect 38770 25062 38800 25114
rect 1344 25028 38800 25062
rect 13078 24946 13130 24958
rect 15206 24946 15258 24958
rect 14354 24894 14366 24946
rect 14418 24943 14430 24946
rect 14690 24943 14702 24946
rect 14418 24897 14702 24943
rect 14418 24894 14430 24897
rect 14690 24894 14702 24897
rect 14754 24894 14766 24946
rect 13078 24882 13130 24894
rect 15206 24882 15258 24894
rect 24614 24946 24666 24958
rect 24614 24882 24666 24894
rect 30830 24946 30882 24958
rect 30830 24882 30882 24894
rect 32174 24946 32226 24958
rect 32174 24882 32226 24894
rect 33742 24946 33794 24958
rect 33742 24882 33794 24894
rect 4734 24834 4786 24846
rect 23998 24834 24050 24846
rect 5562 24782 5574 24834
rect 5626 24782 5638 24834
rect 4734 24770 4786 24782
rect 18286 24778 18338 24790
rect 19518 24778 19570 24790
rect 2046 24722 2098 24734
rect 5070 24722 5122 24734
rect 2818 24670 2830 24722
rect 2882 24670 2894 24722
rect 2046 24658 2098 24670
rect 5070 24658 5122 24670
rect 5294 24722 5346 24734
rect 5294 24658 5346 24670
rect 7758 24722 7810 24734
rect 7758 24658 7810 24670
rect 8318 24722 8370 24734
rect 8990 24722 9042 24734
rect 8318 24658 8370 24670
rect 8822 24666 8874 24678
rect 6638 24610 6690 24622
rect 8990 24658 9042 24670
rect 12686 24722 12738 24734
rect 15026 24670 15038 24722
rect 15090 24670 15102 24722
rect 17602 24714 17614 24766
rect 17666 24714 17678 24766
rect 17826 24670 17838 24722
rect 17890 24670 17902 24722
rect 18286 24714 18338 24726
rect 18398 24750 18450 24762
rect 18398 24686 18450 24698
rect 18678 24757 18730 24769
rect 18834 24726 18846 24778
rect 18898 24726 18910 24778
rect 19518 24714 19570 24726
rect 19630 24750 19682 24762
rect 18678 24693 18730 24705
rect 19630 24686 19682 24698
rect 19910 24757 19962 24769
rect 20066 24726 20078 24778
rect 20130 24726 20142 24778
rect 23998 24770 24050 24782
rect 30158 24834 30210 24846
rect 34682 24782 34694 24834
rect 34746 24782 34758 24834
rect 30158 24770 30210 24782
rect 19910 24693 19962 24705
rect 20358 24722 20410 24734
rect 12686 24658 12738 24670
rect 20358 24658 20410 24670
rect 20638 24722 20690 24734
rect 20638 24658 20690 24670
rect 21310 24722 21362 24734
rect 29026 24670 29038 24722
rect 29090 24670 29102 24722
rect 29250 24714 29262 24766
rect 29314 24714 29326 24766
rect 29822 24722 29874 24734
rect 21310 24658 21362 24670
rect 29822 24658 29874 24670
rect 30494 24722 30546 24734
rect 31378 24670 31390 24722
rect 31442 24670 31454 24722
rect 31602 24714 31614 24766
rect 31666 24714 31678 24766
rect 32510 24722 32562 24734
rect 30494 24658 30546 24670
rect 32510 24658 32562 24670
rect 33406 24722 33458 24734
rect 33406 24658 33458 24670
rect 34974 24722 35026 24734
rect 34974 24658 35026 24670
rect 35198 24722 35250 24734
rect 35198 24658 35250 24670
rect 37214 24722 37266 24734
rect 37214 24658 37266 24670
rect 37886 24722 37938 24734
rect 37886 24658 37938 24670
rect 8822 24602 8874 24614
rect 20974 24610 21026 24622
rect 37550 24610 37602 24622
rect 17490 24558 17502 24610
rect 17554 24558 17566 24610
rect 22082 24558 22094 24610
rect 22146 24558 22158 24610
rect 29362 24558 29374 24610
rect 29426 24558 29438 24610
rect 31714 24558 31726 24610
rect 31778 24558 31790 24610
rect 6638 24546 6690 24558
rect 20974 24546 21026 24558
rect 37550 24546 37602 24558
rect 38278 24610 38330 24622
rect 38278 24546 38330 24558
rect 8076 24498 8128 24510
rect 8076 24434 8128 24446
rect 12350 24498 12402 24510
rect 12350 24434 12402 24446
rect 19126 24498 19178 24510
rect 36094 24498 36146 24510
rect 25330 24446 25342 24498
rect 25394 24495 25406 24498
rect 26226 24495 26238 24498
rect 25394 24449 26238 24495
rect 25394 24446 25406 24449
rect 26226 24446 26238 24449
rect 26290 24495 26302 24498
rect 26562 24495 26574 24498
rect 26290 24449 26574 24495
rect 26290 24446 26302 24449
rect 26562 24446 26574 24449
rect 26626 24446 26638 24498
rect 27122 24446 27134 24498
rect 27186 24495 27198 24498
rect 27682 24495 27694 24498
rect 27186 24449 27694 24495
rect 27186 24446 27198 24449
rect 27682 24446 27694 24449
rect 27746 24446 27758 24498
rect 19126 24434 19178 24446
rect 36094 24434 36146 24446
rect 1344 24330 38640 24364
rect 1344 24278 5876 24330
rect 5928 24278 5980 24330
rect 6032 24278 6084 24330
rect 6136 24278 15200 24330
rect 15252 24278 15304 24330
rect 15356 24278 15408 24330
rect 15460 24278 24524 24330
rect 24576 24278 24628 24330
rect 24680 24278 24732 24330
rect 24784 24278 33848 24330
rect 33900 24278 33952 24330
rect 34004 24278 34056 24330
rect 34108 24278 38640 24330
rect 1344 24244 38640 24278
rect 3838 24162 3890 24174
rect 3838 24098 3890 24110
rect 5742 24162 5794 24174
rect 5742 24098 5794 24110
rect 18416 24162 18468 24174
rect 18416 24098 18468 24110
rect 19574 24162 19626 24174
rect 25342 24162 25394 24174
rect 20010 24110 20022 24162
rect 20074 24110 20086 24162
rect 32286 24162 32338 24174
rect 19574 24098 19626 24110
rect 25342 24098 25394 24110
rect 28142 24106 28194 24118
rect 10278 24050 10330 24062
rect 7186 23998 7198 24050
rect 7250 23998 7262 24050
rect 10278 23986 10330 23998
rect 11510 24050 11562 24062
rect 24502 24050 24554 24062
rect 11510 23986 11562 23998
rect 12742 23994 12794 24006
rect 4958 23938 5010 23950
rect 4958 23874 5010 23886
rect 6078 23938 6130 23950
rect 9886 23938 9938 23950
rect 9090 23886 9102 23938
rect 9154 23886 9166 23938
rect 6078 23874 6130 23886
rect 9886 23874 9938 23886
rect 12238 23938 12290 23950
rect 13638 23994 13690 24006
rect 12742 23930 12794 23942
rect 12910 23938 12962 23950
rect 12238 23874 12290 23886
rect 17670 23994 17722 24006
rect 13638 23930 13690 23942
rect 14142 23938 14194 23950
rect 12910 23874 12962 23886
rect 14142 23874 14194 23886
rect 14702 23938 14754 23950
rect 14702 23874 14754 23886
rect 16718 23938 16770 23950
rect 16718 23874 16770 23886
rect 17502 23938 17554 23950
rect 19014 23994 19066 24006
rect 23874 23998 23886 24050
rect 23938 23998 23950 24050
rect 17670 23930 17722 23942
rect 18174 23938 18226 23950
rect 17502 23874 17554 23886
rect 18174 23874 18226 23886
rect 18846 23938 18898 23950
rect 24502 23986 24554 23998
rect 26910 24050 26962 24062
rect 28142 24042 28194 24054
rect 29654 24050 29706 24062
rect 26910 23986 26962 23998
rect 29654 23986 29706 23998
rect 30326 24050 30378 24062
rect 30818 24054 30830 24106
rect 30882 24054 30894 24106
rect 32286 24098 32338 24110
rect 30326 23986 30378 23998
rect 34582 24050 34634 24062
rect 34850 23998 34862 24050
rect 34914 23998 34926 24050
rect 34582 23986 34634 23998
rect 35814 23994 35866 24006
rect 19014 23930 19066 23942
rect 19294 23938 19346 23950
rect 19170 23886 19182 23938
rect 19234 23886 19246 23938
rect 18846 23874 18898 23886
rect 19294 23874 19346 23886
rect 20302 23938 20354 23950
rect 20302 23874 20354 23886
rect 20414 23938 20466 23950
rect 20414 23874 20466 23886
rect 21198 23938 21250 23950
rect 25678 23938 25730 23950
rect 27246 23938 27298 23950
rect 21970 23886 21982 23938
rect 22034 23886 22046 23938
rect 26562 23886 26574 23938
rect 26626 23886 26638 23938
rect 21198 23874 21250 23886
rect 25678 23874 25730 23886
rect 11996 23826 12048 23838
rect 11996 23762 12048 23774
rect 14384 23826 14436 23838
rect 27010 23830 27022 23882
rect 27074 23830 27086 23882
rect 27246 23874 27298 23886
rect 27582 23938 27634 23950
rect 31838 23938 31890 23950
rect 28242 23886 28254 23938
rect 28306 23886 28318 23938
rect 28578 23886 28590 23938
rect 28642 23886 28654 23938
rect 30706 23886 30718 23938
rect 30770 23886 30782 23938
rect 30930 23886 30942 23938
rect 30994 23886 31006 23938
rect 27582 23874 27634 23886
rect 31838 23874 31890 23886
rect 31950 23938 32002 23950
rect 35646 23938 35698 23950
rect 31950 23874 32002 23886
rect 34962 23842 34974 23894
rect 35026 23842 35038 23894
rect 35298 23886 35310 23938
rect 35362 23886 35374 23938
rect 37830 23994 37882 24006
rect 35814 23930 35866 23942
rect 36094 23938 36146 23950
rect 35970 23886 35982 23938
rect 36034 23886 36046 23938
rect 35646 23874 35698 23886
rect 36094 23874 36146 23886
rect 36374 23938 36426 23950
rect 36374 23874 36426 23886
rect 37326 23938 37378 23950
rect 37830 23930 37882 23942
rect 37998 23938 38050 23950
rect 37326 23874 37378 23886
rect 37998 23874 38050 23886
rect 6470 23714 6522 23726
rect 6470 23650 6522 23662
rect 10838 23714 10890 23726
rect 13570 23718 13582 23770
rect 13634 23718 13646 23770
rect 14384 23762 14436 23774
rect 37084 23826 37136 23838
rect 37084 23762 37136 23774
rect 10838 23650 10890 23662
rect 15038 23714 15090 23726
rect 15038 23650 15090 23662
rect 17054 23714 17106 23726
rect 17054 23650 17106 23662
rect 31502 23714 31554 23726
rect 31502 23650 31554 23662
rect 1344 23546 38800 23580
rect 1344 23494 10538 23546
rect 10590 23494 10642 23546
rect 10694 23494 10746 23546
rect 10798 23494 19862 23546
rect 19914 23494 19966 23546
rect 20018 23494 20070 23546
rect 20122 23494 29186 23546
rect 29238 23494 29290 23546
rect 29342 23494 29394 23546
rect 29446 23494 38510 23546
rect 38562 23494 38614 23546
rect 38666 23494 38718 23546
rect 38770 23494 38800 23546
rect 1344 23460 38800 23494
rect 4286 23378 4338 23390
rect 4286 23314 4338 23326
rect 8654 23378 8706 23390
rect 8654 23314 8706 23326
rect 11118 23378 11170 23390
rect 11118 23314 11170 23326
rect 15654 23378 15706 23390
rect 15654 23314 15706 23326
rect 16606 23378 16658 23390
rect 16606 23314 16658 23326
rect 20750 23378 20802 23390
rect 20750 23314 20802 23326
rect 28646 23378 28698 23390
rect 28646 23314 28698 23326
rect 37998 23378 38050 23390
rect 37998 23314 38050 23326
rect 6246 23266 6298 23278
rect 6246 23202 6298 23214
rect 10558 23266 10610 23278
rect 10558 23202 10610 23214
rect 14254 23266 14306 23278
rect 20078 23266 20130 23278
rect 18330 23214 18342 23266
rect 18394 23214 18406 23266
rect 18778 23214 18790 23266
rect 18842 23214 18854 23266
rect 14254 23202 14306 23214
rect 20078 23202 20130 23214
rect 36412 23266 36464 23278
rect 4622 23154 4674 23166
rect 6862 23154 6914 23166
rect 6570 23102 6582 23154
rect 6634 23102 6646 23154
rect 4622 23090 4674 23102
rect 6862 23090 6914 23102
rect 7086 23154 7138 23166
rect 7086 23090 7138 23102
rect 7198 23154 7250 23166
rect 7198 23090 7250 23102
rect 9886 23154 9938 23166
rect 10782 23154 10834 23166
rect 9886 23090 9938 23102
rect 10390 23098 10442 23110
rect 5014 23042 5066 23054
rect 10782 23090 10834 23102
rect 11566 23154 11618 23166
rect 14590 23154 14642 23166
rect 12338 23102 12350 23154
rect 12402 23102 12414 23154
rect 11566 23090 11618 23102
rect 14590 23090 14642 23102
rect 14814 23154 14866 23166
rect 14814 23090 14866 23102
rect 16942 23154 16994 23166
rect 16942 23090 16994 23102
rect 17950 23154 18002 23166
rect 17950 23090 18002 23102
rect 18062 23154 18114 23166
rect 18062 23090 18114 23102
rect 19070 23154 19122 23166
rect 19070 23090 19122 23102
rect 19294 23154 19346 23166
rect 19294 23090 19346 23102
rect 19742 23154 19794 23166
rect 19742 23090 19794 23102
rect 20414 23154 20466 23166
rect 27134 23154 27186 23166
rect 22418 23102 22430 23154
rect 22482 23102 22494 23154
rect 22754 23102 22766 23154
rect 22818 23102 22830 23154
rect 25554 23102 25566 23154
rect 25618 23102 25630 23154
rect 26338 23102 26350 23154
rect 26402 23102 26414 23154
rect 20414 23090 20466 23102
rect 27134 23090 27186 23102
rect 27470 23154 27522 23166
rect 27794 23158 27806 23210
rect 27858 23158 27870 23210
rect 36412 23202 36464 23214
rect 37326 23266 37378 23278
rect 28018 23102 28030 23154
rect 28082 23102 28094 23154
rect 29026 23102 29038 23154
rect 29090 23102 29102 23154
rect 29250 23102 29262 23154
rect 29314 23102 29326 23154
rect 29810 23146 29822 23198
rect 29874 23146 29886 23198
rect 30494 23154 30546 23166
rect 31614 23154 31666 23166
rect 34526 23154 34578 23166
rect 30146 23102 30158 23154
rect 30210 23102 30222 23154
rect 31042 23102 31054 23154
rect 31106 23102 31118 23154
rect 32274 23102 32286 23154
rect 32338 23102 32350 23154
rect 27470 23090 27522 23102
rect 30494 23090 30546 23102
rect 31614 23090 31666 23102
rect 34526 23090 34578 23102
rect 35422 23154 35474 23166
rect 35422 23090 35474 23102
rect 35758 23154 35810 23166
rect 35758 23090 35810 23102
rect 36654 23154 36706 23166
rect 37146 23158 37158 23210
rect 37210 23158 37222 23210
rect 37326 23202 37378 23214
rect 36654 23090 36706 23102
rect 38334 23154 38386 23166
rect 38334 23090 38386 23102
rect 10390 23034 10442 23046
rect 16102 23042 16154 23054
rect 5014 22978 5066 22990
rect 25342 23042 25394 23054
rect 16102 22978 16154 22990
rect 22318 22986 22370 22998
rect 9644 22930 9696 22942
rect 27906 22990 27918 23042
rect 27970 22990 27982 23042
rect 29698 22990 29710 23042
rect 29762 22990 29774 23042
rect 25342 22978 25394 22990
rect 29026 22934 29038 22986
rect 29090 22934 29102 22986
rect 31266 22934 31278 22986
rect 31330 22934 31342 22986
rect 32386 22934 32398 22986
rect 32450 22934 32462 22986
rect 15082 22878 15094 22930
rect 15146 22878 15158 22930
rect 22318 22922 22370 22934
rect 34862 22930 34914 22942
rect 9644 22866 9696 22878
rect 34862 22866 34914 22878
rect 1344 22762 38640 22796
rect 1344 22710 5876 22762
rect 5928 22710 5980 22762
rect 6032 22710 6084 22762
rect 6136 22710 15200 22762
rect 15252 22710 15304 22762
rect 15356 22710 15408 22762
rect 15460 22710 24524 22762
rect 24576 22710 24628 22762
rect 24680 22710 24732 22762
rect 24784 22710 33848 22762
rect 33900 22710 33952 22762
rect 34004 22710 34056 22762
rect 34108 22710 38640 22762
rect 1344 22676 38640 22710
rect 19966 22594 20018 22606
rect 12394 22542 12406 22594
rect 12458 22542 12470 22594
rect 19966 22530 20018 22542
rect 29150 22538 29202 22550
rect 19462 22482 19514 22494
rect 10994 22430 11006 22482
rect 11058 22430 11070 22482
rect 18722 22430 18734 22482
rect 18786 22430 18798 22482
rect 19462 22418 19514 22430
rect 26014 22482 26066 22494
rect 27906 22430 27918 22482
rect 27970 22430 27982 22482
rect 29150 22474 29202 22486
rect 31502 22538 31554 22550
rect 31502 22474 31554 22486
rect 32174 22482 32226 22494
rect 26014 22418 26066 22430
rect 32174 22418 32226 22430
rect 38278 22482 38330 22494
rect 38278 22418 38330 22430
rect 2942 22370 2994 22382
rect 2942 22306 2994 22318
rect 3166 22370 3218 22382
rect 3166 22306 3218 22318
rect 5182 22370 5234 22382
rect 5182 22306 5234 22318
rect 7982 22370 8034 22382
rect 7982 22306 8034 22318
rect 8206 22370 8258 22382
rect 8206 22306 8258 22318
rect 8318 22370 8370 22382
rect 11902 22370 11954 22382
rect 9090 22318 9102 22370
rect 9154 22318 9166 22370
rect 8318 22306 8370 22318
rect 11902 22306 11954 22318
rect 12126 22370 12178 22382
rect 12126 22306 12178 22318
rect 14030 22370 14082 22382
rect 16046 22370 16098 22382
rect 19630 22370 19682 22382
rect 15474 22318 15486 22370
rect 15538 22318 15550 22370
rect 16818 22318 16830 22370
rect 16882 22318 16894 22370
rect 14030 22306 14082 22318
rect 16046 22306 16098 22318
rect 19630 22306 19682 22318
rect 23214 22370 23266 22382
rect 23214 22306 23266 22318
rect 23438 22370 23490 22382
rect 26350 22370 26402 22382
rect 28142 22370 28194 22382
rect 30494 22370 30546 22382
rect 32510 22370 32562 22382
rect 23706 22318 23718 22370
rect 23770 22318 23782 22370
rect 25666 22318 25678 22370
rect 25730 22318 25742 22370
rect 27570 22318 27582 22370
rect 27634 22318 27646 22370
rect 29250 22318 29262 22370
rect 29314 22318 29326 22370
rect 29474 22318 29486 22370
rect 29538 22318 29550 22370
rect 23438 22306 23490 22318
rect 4062 22258 4114 22270
rect 26114 22262 26126 22314
rect 26178 22262 26190 22314
rect 26350 22306 26402 22318
rect 28142 22306 28194 22318
rect 30494 22306 30546 22318
rect 30702 22280 30714 22332
rect 30766 22280 30778 22332
rect 31378 22318 31390 22370
rect 31442 22318 31454 22370
rect 31826 22318 31838 22370
rect 31890 22318 31902 22370
rect 32162 22262 32174 22314
rect 32226 22262 32238 22314
rect 32510 22306 32562 22318
rect 32846 22370 32898 22382
rect 32846 22306 32898 22318
rect 33406 22370 33458 22382
rect 33406 22306 33458 22318
rect 34078 22370 34130 22382
rect 33562 22262 33574 22314
rect 33626 22262 33638 22314
rect 34078 22306 34130 22318
rect 34638 22370 34690 22382
rect 34638 22306 34690 22318
rect 34862 22370 34914 22382
rect 34862 22306 34914 22318
rect 34320 22258 34372 22270
rect 2650 22206 2662 22258
rect 2714 22206 2726 22258
rect 7690 22206 7702 22258
rect 7754 22206 7766 22258
rect 35130 22206 35142 22258
rect 35194 22206 35206 22258
rect 4062 22194 4114 22206
rect 34320 22194 34372 22206
rect 5798 22146 5850 22158
rect 5798 22082 5850 22094
rect 7366 22146 7418 22158
rect 7366 22082 7418 22094
rect 30158 22146 30210 22158
rect 30158 22082 30210 22094
rect 1344 21978 38800 22012
rect 1344 21926 10538 21978
rect 10590 21926 10642 21978
rect 10694 21926 10746 21978
rect 10798 21926 19862 21978
rect 19914 21926 19966 21978
rect 20018 21926 20070 21978
rect 20122 21926 29186 21978
rect 29238 21926 29290 21978
rect 29342 21926 29394 21978
rect 29446 21926 38510 21978
rect 38562 21926 38614 21978
rect 38666 21926 38718 21978
rect 38770 21926 38800 21978
rect 1344 21892 38800 21926
rect 6694 21810 6746 21822
rect 6694 21746 6746 21758
rect 15878 21810 15930 21822
rect 15878 21746 15930 21758
rect 18342 21810 18394 21822
rect 18342 21746 18394 21758
rect 19070 21810 19122 21822
rect 19070 21746 19122 21758
rect 5276 21698 5328 21710
rect 5276 21634 5328 21646
rect 6190 21698 6242 21710
rect 2046 21586 2098 21598
rect 2046 21522 2098 21534
rect 5518 21586 5570 21598
rect 6010 21590 6022 21642
rect 6074 21590 6086 21642
rect 6190 21634 6242 21646
rect 12686 21698 12738 21710
rect 33338 21646 33350 21698
rect 33402 21646 33414 21698
rect 12686 21634 12738 21646
rect 25510 21615 25562 21627
rect 5518 21522 5570 21534
rect 11566 21586 11618 21598
rect 11566 21522 11618 21534
rect 11790 21586 11842 21598
rect 11790 21522 11842 21534
rect 13806 21586 13858 21598
rect 13806 21522 13858 21534
rect 14478 21586 14530 21598
rect 19406 21586 19458 21598
rect 18162 21534 18174 21586
rect 18226 21534 18238 21586
rect 14478 21522 14530 21534
rect 19406 21522 19458 21534
rect 19798 21586 19850 21598
rect 19798 21522 19850 21534
rect 21646 21586 21698 21598
rect 25218 21534 25230 21586
rect 25282 21534 25294 21586
rect 26574 21625 26626 21637
rect 25510 21551 25562 21563
rect 26114 21534 26126 21586
rect 26178 21534 26190 21586
rect 26574 21561 26626 21573
rect 26798 21586 26850 21598
rect 21646 21522 21698 21534
rect 26798 21522 26850 21534
rect 27134 21586 27186 21598
rect 27134 21522 27186 21534
rect 27582 21586 27634 21598
rect 27582 21522 27634 21534
rect 27806 21586 27858 21598
rect 30158 21586 30210 21598
rect 30370 21590 30382 21642
rect 30434 21590 30446 21642
rect 31938 21590 31950 21642
rect 32002 21590 32014 21642
rect 32286 21586 32338 21598
rect 28578 21534 28590 21586
rect 28642 21534 28654 21586
rect 28914 21534 28926 21586
rect 28978 21534 28990 21586
rect 30706 21534 30718 21586
rect 30770 21534 30782 21586
rect 31602 21534 31614 21586
rect 31666 21534 31678 21586
rect 27806 21522 27858 21534
rect 30158 21522 30210 21534
rect 32286 21522 32338 21534
rect 33630 21586 33682 21598
rect 33630 21522 33682 21534
rect 33742 21586 33794 21598
rect 33742 21522 33794 21534
rect 33966 21586 34018 21598
rect 33966 21522 34018 21534
rect 35982 21586 36034 21598
rect 35982 21522 36034 21534
rect 8374 21474 8426 21486
rect 2818 21422 2830 21474
rect 2882 21422 2894 21474
rect 4722 21422 4734 21474
rect 4786 21422 4798 21474
rect 8374 21410 8426 21422
rect 24054 21474 24106 21486
rect 31334 21474 31386 21486
rect 25666 21422 25678 21474
rect 25730 21422 25742 21474
rect 26226 21422 26238 21474
rect 26290 21422 26302 21474
rect 28074 21422 28086 21474
rect 28138 21422 28150 21474
rect 24054 21410 24106 21422
rect 28478 21418 28530 21430
rect 30594 21422 30606 21474
rect 30658 21422 30670 21474
rect 14142 21362 14194 21374
rect 11274 21310 11286 21362
rect 11338 21310 11350 21362
rect 14142 21298 14194 21310
rect 21982 21362 22034 21374
rect 31334 21410 31386 21422
rect 31950 21474 32002 21486
rect 31950 21410 32002 21422
rect 28478 21354 28530 21366
rect 35422 21362 35474 21374
rect 21982 21298 22034 21310
rect 35422 21298 35474 21310
rect 37438 21362 37490 21374
rect 37438 21298 37490 21310
rect 1344 21194 38640 21228
rect 1344 21142 5876 21194
rect 5928 21142 5980 21194
rect 6032 21142 6084 21194
rect 6136 21142 15200 21194
rect 15252 21142 15304 21194
rect 15356 21142 15408 21194
rect 15460 21142 24524 21194
rect 24576 21142 24628 21194
rect 24680 21142 24732 21194
rect 24784 21142 33848 21194
rect 33900 21142 33952 21194
rect 34004 21142 34056 21194
rect 34108 21142 38640 21194
rect 1344 21108 38640 21142
rect 3166 21026 3218 21038
rect 3166 20962 3218 20974
rect 9326 21026 9378 21038
rect 9326 20962 9378 20974
rect 13564 21026 13616 21038
rect 13564 20962 13616 20974
rect 19406 21026 19458 21038
rect 19406 20962 19458 20974
rect 22094 21026 22146 21038
rect 22094 20962 22146 20974
rect 24838 21026 24890 21038
rect 24838 20962 24890 20974
rect 37904 21026 37956 21038
rect 20190 20914 20242 20926
rect 25666 20918 25678 20970
rect 25730 20918 25742 20970
rect 37904 20962 37956 20974
rect 6470 20858 6522 20870
rect 2046 20802 2098 20814
rect 2046 20738 2098 20750
rect 4958 20802 5010 20814
rect 4958 20738 5010 20750
rect 5182 20802 5234 20814
rect 5182 20738 5234 20750
rect 5724 20802 5776 20814
rect 5724 20738 5776 20750
rect 5966 20802 6018 20814
rect 35746 20862 35758 20914
rect 35810 20862 35822 20914
rect 20190 20850 20242 20862
rect 6470 20794 6522 20806
rect 6638 20802 6690 20814
rect 5966 20738 6018 20750
rect 6638 20738 6690 20750
rect 7310 20802 7362 20814
rect 7310 20738 7362 20750
rect 7814 20802 7866 20814
rect 7814 20738 7866 20750
rect 8206 20802 8258 20814
rect 8206 20738 8258 20750
rect 11118 20802 11170 20814
rect 11118 20738 11170 20750
rect 13806 20802 13858 20814
rect 13806 20738 13858 20750
rect 14478 20802 14530 20814
rect 7068 20690 7120 20702
rect 4666 20638 4678 20690
rect 4730 20638 4742 20690
rect 7068 20626 7120 20638
rect 7982 20690 8034 20702
rect 14298 20694 14310 20746
rect 14362 20694 14374 20746
rect 14478 20738 14530 20750
rect 19070 20802 19122 20814
rect 20526 20802 20578 20814
rect 19842 20750 19854 20802
rect 19906 20750 19918 20802
rect 24110 20802 24162 20814
rect 19070 20738 19122 20750
rect 20290 20694 20302 20746
rect 20354 20694 20366 20746
rect 20526 20738 20578 20750
rect 23762 20722 23774 20774
rect 23826 20722 23838 20774
rect 24110 20738 24162 20750
rect 24558 20802 24610 20814
rect 26126 20802 26178 20814
rect 25554 20750 25566 20802
rect 25618 20750 25630 20802
rect 25778 20750 25790 20802
rect 25842 20750 25854 20802
rect 24266 20694 24278 20746
rect 24330 20694 24342 20746
rect 24558 20738 24610 20750
rect 26126 20738 26178 20750
rect 30326 20802 30378 20814
rect 32062 20802 32114 20814
rect 31378 20750 31390 20802
rect 31442 20750 31454 20802
rect 30326 20738 30378 20750
rect 32062 20738 32114 20750
rect 32286 20802 32338 20814
rect 32286 20738 32338 20750
rect 33854 20802 33906 20814
rect 33854 20738 33906 20750
rect 36542 20802 36594 20814
rect 36542 20738 36594 20750
rect 36990 20802 37042 20814
rect 36990 20738 37042 20750
rect 37158 20802 37210 20814
rect 37158 20738 37210 20750
rect 37662 20802 37714 20814
rect 37662 20738 37714 20750
rect 7982 20626 8034 20638
rect 24446 20690 24498 20702
rect 24446 20626 24498 20638
rect 31726 20690 31778 20702
rect 32554 20638 32566 20690
rect 32618 20638 32630 20690
rect 31726 20626 31778 20638
rect 12574 20578 12626 20590
rect 12574 20514 12626 20526
rect 14982 20578 15034 20590
rect 26462 20578 26514 20590
rect 15306 20526 15318 20578
rect 15370 20575 15382 20578
rect 15922 20575 15934 20578
rect 15370 20529 15934 20575
rect 15370 20526 15382 20529
rect 15922 20526 15934 20529
rect 15986 20526 15998 20578
rect 14982 20514 15034 20526
rect 26462 20514 26514 20526
rect 27078 20578 27130 20590
rect 27078 20514 27130 20526
rect 1344 20410 38800 20444
rect 1344 20358 10538 20410
rect 10590 20358 10642 20410
rect 10694 20358 10746 20410
rect 10798 20358 19862 20410
rect 19914 20358 19966 20410
rect 20018 20358 20070 20410
rect 20122 20358 29186 20410
rect 29238 20358 29290 20410
rect 29342 20358 29394 20410
rect 29446 20358 38510 20410
rect 38562 20358 38614 20410
rect 38666 20358 38718 20410
rect 38770 20358 38800 20410
rect 1344 20324 38800 20358
rect 15318 20242 15370 20254
rect 9606 20186 9658 20198
rect 6862 20130 6914 20142
rect 6862 20066 6914 20078
rect 7310 20130 7362 20142
rect 25846 20242 25898 20254
rect 15318 20178 15370 20190
rect 19910 20186 19962 20198
rect 9606 20122 9658 20134
rect 14702 20130 14754 20142
rect 7310 20066 7362 20078
rect 25846 20178 25898 20190
rect 19910 20122 19962 20134
rect 33294 20130 33346 20142
rect 3838 20018 3890 20030
rect 3838 19954 3890 19966
rect 4062 20018 4114 20030
rect 4062 19954 4114 19966
rect 4174 20018 4226 20030
rect 7466 20022 7478 20074
rect 7530 20022 7542 20074
rect 14702 20066 14754 20078
rect 20302 20053 20354 20065
rect 4174 19954 4226 19966
rect 7982 20018 8034 20030
rect 12014 20018 12066 20030
rect 9426 19966 9438 20018
rect 9490 19966 9502 20018
rect 12786 19966 12798 20018
rect 12850 19966 12862 20018
rect 20066 19966 20078 20018
rect 20130 19966 20142 20018
rect 20302 19989 20354 20001
rect 20414 20046 20466 20058
rect 20414 19982 20466 19994
rect 20638 20046 20690 20058
rect 20638 19982 20690 19994
rect 20912 20046 20964 20058
rect 20912 19982 20964 19994
rect 21422 20018 21474 20030
rect 23438 20018 23490 20030
rect 22866 19966 22878 20018
rect 22930 19966 22942 20018
rect 7982 19954 8034 19966
rect 12014 19954 12066 19966
rect 21422 19954 21474 19966
rect 23438 19954 23490 19966
rect 24110 20018 24162 20030
rect 29038 20018 29090 20030
rect 25442 19966 25454 20018
rect 25506 19966 25518 20018
rect 24110 19954 24162 19966
rect 29038 19954 29090 19966
rect 29262 20018 29314 20030
rect 30258 20022 30270 20074
rect 30322 20022 30334 20074
rect 33294 20066 33346 20078
rect 34208 20130 34260 20142
rect 30606 20018 30658 20030
rect 29530 19966 29542 20018
rect 29594 19966 29606 20018
rect 29922 19966 29934 20018
rect 29986 19966 29998 20018
rect 29262 19954 29314 19966
rect 30606 19954 30658 19966
rect 30942 20018 30994 20030
rect 30942 19954 30994 19966
rect 31390 20018 31442 20030
rect 31390 19954 31442 19966
rect 31614 20018 31666 20030
rect 33450 20022 33462 20074
rect 33514 20022 33526 20074
rect 34208 20066 34260 20078
rect 35646 20130 35698 20142
rect 35646 20066 35698 20078
rect 31614 19954 31666 19966
rect 33966 20018 34018 20030
rect 38334 20018 38386 20030
rect 37538 19966 37550 20018
rect 37602 19966 37614 20018
rect 33966 19954 34018 19966
rect 38334 19954 38386 19966
rect 15766 19906 15818 19918
rect 4946 19854 4958 19906
rect 5010 19854 5022 19906
rect 15766 19842 15818 19854
rect 30270 19906 30322 19918
rect 35254 19906 35306 19918
rect 31882 19854 31894 19906
rect 31946 19854 31958 19906
rect 30270 19842 30322 19854
rect 35254 19842 35306 19854
rect 8224 19794 8276 19806
rect 3546 19742 3558 19794
rect 3610 19742 3622 19794
rect 8224 19730 8276 19742
rect 21142 19794 21194 19806
rect 21142 19730 21194 19742
rect 23774 19794 23826 19806
rect 23774 19730 23826 19742
rect 24446 19794 24498 19806
rect 24446 19730 24498 19742
rect 25286 19794 25338 19806
rect 25286 19730 25338 19742
rect 1344 19626 38640 19660
rect 1344 19574 5876 19626
rect 5928 19574 5980 19626
rect 6032 19574 6084 19626
rect 6136 19574 15200 19626
rect 15252 19574 15304 19626
rect 15356 19574 15408 19626
rect 15460 19574 24524 19626
rect 24576 19574 24628 19626
rect 24680 19574 24732 19626
rect 24784 19574 33848 19626
rect 33900 19574 33952 19626
rect 34004 19574 34056 19626
rect 34108 19574 38640 19626
rect 1344 19540 38640 19574
rect 4734 19458 4786 19470
rect 4734 19394 4786 19406
rect 21366 19458 21418 19470
rect 21366 19394 21418 19406
rect 21814 19458 21866 19470
rect 21814 19394 21866 19406
rect 29486 19458 29538 19470
rect 29486 19394 29538 19406
rect 29990 19458 30042 19470
rect 29990 19394 30042 19406
rect 37998 19458 38050 19470
rect 37998 19394 38050 19406
rect 23102 19346 23154 19358
rect 10658 19294 10670 19346
rect 10722 19294 10734 19346
rect 13414 19290 13466 19302
rect 17154 19294 17166 19346
rect 17218 19294 17230 19346
rect 3278 19234 3330 19246
rect 3278 19170 3330 19182
rect 5518 19234 5570 19246
rect 5518 19170 5570 19182
rect 7982 19234 8034 19246
rect 11902 19234 11954 19246
rect 8754 19182 8766 19234
rect 8818 19182 8830 19234
rect 7982 19170 8034 19182
rect 11902 19170 11954 19182
rect 12574 19234 12626 19246
rect 23102 19282 23154 19294
rect 25006 19346 25058 19358
rect 32342 19346 32394 19358
rect 25006 19282 25058 19294
rect 31894 19290 31946 19302
rect 13414 19226 13466 19238
rect 14478 19234 14530 19246
rect 17782 19234 17834 19246
rect 13794 19182 13806 19234
rect 13858 19182 13870 19234
rect 14142 19196 14194 19208
rect 12058 19126 12070 19178
rect 12122 19126 12134 19178
rect 12574 19170 12626 19182
rect 15250 19182 15262 19234
rect 15314 19182 15326 19234
rect 14478 19170 14530 19182
rect 17782 19170 17834 19182
rect 18846 19234 18898 19246
rect 20526 19234 20578 19246
rect 22430 19234 22482 19246
rect 19506 19182 19518 19234
rect 19570 19182 19582 19234
rect 19954 19182 19966 19234
rect 20018 19182 20030 19234
rect 21522 19182 21534 19234
rect 21586 19182 21598 19234
rect 21970 19182 21982 19234
rect 22034 19182 22046 19234
rect 18846 19170 18898 19182
rect 12816 19122 12868 19134
rect 12816 19058 12868 19070
rect 13582 19122 13634 19134
rect 14142 19132 14194 19144
rect 19058 19126 19070 19178
rect 19122 19126 19134 19178
rect 20178 19126 20190 19178
rect 20242 19126 20254 19178
rect 20526 19170 20578 19182
rect 22430 19170 22482 19182
rect 22766 19234 22818 19246
rect 23774 19234 23826 19246
rect 22766 19170 22818 19182
rect 22990 19195 23042 19207
rect 23426 19182 23438 19234
rect 23490 19182 23502 19234
rect 23774 19170 23826 19182
rect 23998 19234 24050 19246
rect 25342 19234 25394 19246
rect 26574 19234 26626 19246
rect 24770 19182 24782 19234
rect 24834 19182 24846 19234
rect 25890 19182 25902 19234
rect 25954 19182 25966 19234
rect 23998 19170 24050 19182
rect 22990 19131 23042 19143
rect 24994 19126 25006 19178
rect 25058 19126 25070 19178
rect 25342 19170 25394 19182
rect 26338 19126 26350 19178
rect 26402 19126 26414 19178
rect 26574 19170 26626 19182
rect 27022 19234 27074 19246
rect 27022 19170 27074 19182
rect 27246 19234 27298 19246
rect 27246 19170 27298 19182
rect 29150 19234 29202 19246
rect 29150 19170 29202 19182
rect 30270 19234 30322 19246
rect 30550 19234 30602 19246
rect 30370 19182 30382 19234
rect 30434 19182 30446 19234
rect 30270 19170 30322 19182
rect 30550 19170 30602 19182
rect 30718 19234 30770 19246
rect 31042 19238 31054 19290
rect 31106 19238 31118 19290
rect 32342 19282 32394 19294
rect 37158 19346 37210 19358
rect 37158 19282 37210 19294
rect 31894 19226 31946 19238
rect 37606 19234 37658 19246
rect 30718 19170 30770 19182
rect 31166 19196 31218 19208
rect 37606 19170 37658 19182
rect 38334 19234 38386 19246
rect 38334 19170 38386 19182
rect 31166 19132 31218 19144
rect 31726 19122 31778 19134
rect 24266 19070 24278 19122
rect 24330 19070 24342 19122
rect 27514 19070 27526 19122
rect 27578 19070 27590 19122
rect 13582 19058 13634 19070
rect 6638 19010 6690 19022
rect 6638 18946 6690 18958
rect 7814 19010 7866 19022
rect 7814 18946 7866 18958
rect 11286 19010 11338 19022
rect 19394 19014 19406 19066
rect 19458 19014 19470 19066
rect 20626 19014 20638 19066
rect 20690 19014 20702 19066
rect 26674 19014 26686 19066
rect 26738 19014 26750 19066
rect 31726 19058 31778 19070
rect 11286 18946 11338 18958
rect 1344 18842 38800 18876
rect 1344 18790 10538 18842
rect 10590 18790 10642 18842
rect 10694 18790 10746 18842
rect 10798 18790 19862 18842
rect 19914 18790 19966 18842
rect 20018 18790 20070 18842
rect 20122 18790 29186 18842
rect 29238 18790 29290 18842
rect 29342 18790 29394 18842
rect 29446 18790 38510 18842
rect 38562 18790 38614 18842
rect 38666 18790 38718 18842
rect 38770 18790 38800 18842
rect 1344 18756 38800 18790
rect 15262 18674 15314 18686
rect 15262 18610 15314 18622
rect 8430 18562 8482 18574
rect 8430 18498 8482 18510
rect 12462 18562 12514 18574
rect 5742 18450 5794 18462
rect 9046 18450 9098 18462
rect 6514 18398 6526 18450
rect 6578 18398 6590 18450
rect 5742 18386 5794 18398
rect 9046 18386 9098 18398
rect 9438 18450 9490 18462
rect 9438 18386 9490 18398
rect 9662 18450 9714 18462
rect 9662 18386 9714 18398
rect 11006 18450 11058 18462
rect 11006 18386 11058 18398
rect 11118 18450 11170 18462
rect 11118 18386 11170 18398
rect 11790 18450 11842 18462
rect 12282 18454 12294 18506
rect 12346 18454 12358 18506
rect 12462 18498 12514 18510
rect 19966 18562 20018 18574
rect 29486 18562 29538 18574
rect 19966 18498 20018 18510
rect 21982 18506 22034 18518
rect 23370 18510 23382 18562
rect 23434 18510 23446 18562
rect 11790 18386 11842 18398
rect 12910 18450 12962 18462
rect 12910 18386 12962 18398
rect 13134 18450 13186 18462
rect 13806 18450 13858 18462
rect 13402 18398 13414 18450
rect 13466 18398 13478 18450
rect 13134 18386 13186 18398
rect 13806 18386 13858 18398
rect 17278 18450 17330 18462
rect 20402 18398 20414 18450
rect 20466 18398 20478 18450
rect 20738 18398 20750 18450
rect 20802 18398 20814 18450
rect 21186 18398 21198 18450
rect 21250 18398 21262 18450
rect 21522 18398 21534 18450
rect 21586 18398 21598 18450
rect 21982 18442 22034 18454
rect 22094 18478 22146 18490
rect 22094 18414 22146 18426
rect 22318 18478 22370 18490
rect 22318 18414 22370 18426
rect 22542 18478 22594 18490
rect 22542 18414 22594 18426
rect 23662 18450 23714 18462
rect 17278 18386 17330 18398
rect 23662 18386 23714 18398
rect 23774 18450 23826 18462
rect 23774 18386 23826 18398
rect 24110 18450 24162 18462
rect 24110 18386 24162 18398
rect 24334 18450 24386 18462
rect 25890 18454 25902 18506
rect 25954 18454 25966 18506
rect 29486 18498 29538 18510
rect 26238 18450 26290 18462
rect 24602 18398 24614 18450
rect 24666 18398 24678 18450
rect 25554 18398 25566 18450
rect 25618 18398 25630 18450
rect 24334 18386 24386 18398
rect 26238 18386 26290 18398
rect 26686 18450 26738 18462
rect 26686 18386 26738 18398
rect 26910 18450 26962 18462
rect 26910 18386 26962 18398
rect 28030 18450 28082 18462
rect 28030 18386 28082 18398
rect 29374 18450 29426 18462
rect 29822 18450 29874 18462
rect 29374 18386 29426 18398
rect 29654 18394 29706 18406
rect 20302 18338 20354 18350
rect 18050 18286 18062 18338
rect 18114 18286 18126 18338
rect 20302 18274 20354 18286
rect 22822 18338 22874 18350
rect 22822 18274 22874 18286
rect 25902 18338 25954 18350
rect 25902 18274 25954 18286
rect 27694 18338 27746 18350
rect 30258 18398 30270 18450
rect 30322 18398 30334 18450
rect 30998 18436 31010 18488
rect 31062 18436 31074 18488
rect 33966 18450 34018 18462
rect 31154 18398 31166 18450
rect 31218 18398 31230 18450
rect 29822 18386 29874 18398
rect 33966 18386 34018 18398
rect 34190 18450 34242 18462
rect 34750 18450 34802 18462
rect 34458 18398 34470 18450
rect 34522 18398 34534 18450
rect 35746 18398 35758 18450
rect 35810 18398 35822 18450
rect 34190 18386 34242 18398
rect 34750 18386 34802 18398
rect 29654 18330 29706 18342
rect 33798 18338 33850 18350
rect 27694 18274 27746 18286
rect 30158 18282 30210 18294
rect 11548 18226 11600 18238
rect 29094 18226 29146 18238
rect 9930 18174 9942 18226
rect 9994 18174 10006 18226
rect 10714 18174 10726 18226
rect 10778 18174 10790 18226
rect 27178 18174 27190 18226
rect 27242 18174 27254 18226
rect 30158 18218 30210 18230
rect 31334 18282 31386 18294
rect 33798 18274 33850 18286
rect 35926 18282 35978 18294
rect 31334 18218 31386 18230
rect 35086 18226 35138 18238
rect 11548 18162 11600 18174
rect 29094 18162 29146 18174
rect 35926 18218 35978 18230
rect 35086 18162 35138 18174
rect 1344 18058 38640 18092
rect 1344 18006 5876 18058
rect 5928 18006 5980 18058
rect 6032 18006 6084 18058
rect 6136 18006 15200 18058
rect 15252 18006 15304 18058
rect 15356 18006 15408 18058
rect 15460 18006 24524 18058
rect 24576 18006 24628 18058
rect 24680 18006 24732 18058
rect 24784 18006 33848 18058
rect 33900 18006 33952 18058
rect 34004 18006 34056 18058
rect 34108 18006 38640 18058
rect 1344 17972 38640 18006
rect 8542 17890 8594 17902
rect 8542 17826 8594 17838
rect 17838 17890 17890 17902
rect 17838 17826 17890 17838
rect 24334 17834 24386 17846
rect 12674 17726 12686 17778
rect 12738 17726 12750 17778
rect 24334 17770 24386 17782
rect 28646 17778 28698 17790
rect 27078 17722 27130 17734
rect 9662 17666 9714 17678
rect 9662 17602 9714 17614
rect 9998 17666 10050 17678
rect 13358 17666 13410 17678
rect 10770 17614 10782 17666
rect 10834 17614 10846 17666
rect 9998 17602 10050 17614
rect 13358 17602 13410 17614
rect 13582 17666 13634 17678
rect 13582 17602 13634 17614
rect 14142 17666 14194 17678
rect 14142 17602 14194 17614
rect 15094 17666 15146 17678
rect 15094 17602 15146 17614
rect 18174 17666 18226 17678
rect 18174 17602 18226 17614
rect 20750 17666 20802 17678
rect 25174 17666 25226 17678
rect 23874 17614 23886 17666
rect 23938 17614 23950 17666
rect 24210 17614 24222 17666
rect 24274 17614 24286 17666
rect 20750 17602 20802 17614
rect 25174 17602 25226 17614
rect 25454 17666 25506 17678
rect 25902 17666 25954 17678
rect 28646 17714 28698 17726
rect 30494 17778 30546 17790
rect 30494 17714 30546 17726
rect 31110 17778 31162 17790
rect 37158 17778 37210 17790
rect 34402 17726 34414 17778
rect 34466 17726 34478 17778
rect 31110 17714 31162 17726
rect 37158 17714 37210 17726
rect 25554 17614 25566 17666
rect 25618 17614 25630 17666
rect 25454 17602 25506 17614
rect 20022 17554 20074 17566
rect 25722 17558 25734 17610
rect 25786 17558 25798 17610
rect 25902 17602 25954 17614
rect 26450 17586 26462 17638
rect 26514 17586 26526 17638
rect 26674 17614 26686 17666
rect 26738 17614 26750 17666
rect 27078 17658 27130 17670
rect 29822 17666 29874 17678
rect 38334 17666 38386 17678
rect 29362 17614 29374 17666
rect 29426 17614 29438 17666
rect 29922 17614 29934 17666
rect 29986 17614 29998 17666
rect 29822 17602 29874 17614
rect 13850 17502 13862 17554
rect 13914 17502 13926 17554
rect 20022 17490 20074 17502
rect 26910 17554 26962 17566
rect 30088 17558 30100 17610
rect 30152 17558 30164 17610
rect 33674 17588 33686 17640
rect 33738 17588 33750 17640
rect 38334 17602 38386 17614
rect 26910 17490 26962 17502
rect 36318 17554 36370 17566
rect 36318 17490 36370 17502
rect 14478 17442 14530 17454
rect 14478 17378 14530 17390
rect 20414 17442 20466 17454
rect 29206 17442 29258 17454
rect 27458 17390 27470 17442
rect 27522 17439 27534 17442
rect 27794 17439 27806 17442
rect 27522 17393 27806 17439
rect 27522 17390 27534 17393
rect 27794 17390 27806 17393
rect 27858 17390 27870 17442
rect 20414 17378 20466 17390
rect 29206 17378 29258 17390
rect 37606 17442 37658 17454
rect 37606 17378 37658 17390
rect 37998 17442 38050 17454
rect 37998 17378 38050 17390
rect 1344 17274 38800 17308
rect 1344 17222 10538 17274
rect 10590 17222 10642 17274
rect 10694 17222 10746 17274
rect 10798 17222 19862 17274
rect 19914 17222 19966 17274
rect 20018 17222 20070 17274
rect 20122 17222 29186 17274
rect 29238 17222 29290 17274
rect 29342 17222 29394 17274
rect 29446 17222 38510 17274
rect 38562 17222 38614 17274
rect 38666 17222 38718 17274
rect 38770 17222 38800 17274
rect 1344 17188 38800 17222
rect 9718 17106 9770 17118
rect 9718 17042 9770 17054
rect 11006 17106 11058 17118
rect 11006 17042 11058 17054
rect 17558 17106 17610 17118
rect 23046 17106 23098 17118
rect 17558 17042 17610 17054
rect 22486 17050 22538 17062
rect 12350 16994 12402 17006
rect 12350 16930 12402 16942
rect 13264 16994 13316 17006
rect 8654 16882 8706 16894
rect 8654 16818 8706 16830
rect 8990 16882 9042 16894
rect 8990 16818 9042 16830
rect 9886 16882 9938 16894
rect 12506 16886 12518 16938
rect 12570 16886 12582 16938
rect 13264 16930 13316 16942
rect 16382 16994 16434 17006
rect 20066 16998 20078 17050
rect 20130 16998 20142 17050
rect 23046 17042 23098 17054
rect 28142 17106 28194 17118
rect 28142 17042 28194 17054
rect 31110 17106 31162 17118
rect 31110 17042 31162 17054
rect 33686 17106 33738 17118
rect 33686 17042 33738 17054
rect 22486 16986 22538 16998
rect 25902 16994 25954 17006
rect 16382 16930 16434 16942
rect 20414 16938 20466 16950
rect 9886 16818 9938 16830
rect 13022 16882 13074 16894
rect 13022 16818 13074 16830
rect 13694 16882 13746 16894
rect 13694 16818 13746 16830
rect 18790 16882 18842 16894
rect 18790 16818 18842 16830
rect 19294 16882 19346 16894
rect 19954 16830 19966 16882
rect 20018 16830 20030 16882
rect 20414 16874 20466 16886
rect 20526 16910 20578 16922
rect 20738 16886 20750 16938
rect 20802 16886 20814 16938
rect 20962 16886 20974 16938
rect 21026 16886 21038 16938
rect 20526 16846 20578 16858
rect 21254 16882 21306 16894
rect 21746 16874 21758 16926
rect 21810 16874 21822 16926
rect 23550 16882 23602 16894
rect 21970 16830 21982 16882
rect 22034 16830 22046 16882
rect 22306 16830 22318 16882
rect 22370 16830 22382 16882
rect 19294 16818 19346 16830
rect 21254 16818 21306 16830
rect 23550 16818 23602 16830
rect 23662 16882 23714 16894
rect 23662 16818 23714 16830
rect 25566 16882 25618 16894
rect 25722 16886 25734 16938
rect 25786 16886 25798 16938
rect 25902 16930 25954 16942
rect 25566 16818 25618 16830
rect 26014 16882 26066 16894
rect 26014 16818 26066 16830
rect 26294 16882 26346 16894
rect 26294 16818 26346 16830
rect 27806 16882 27858 16894
rect 28578 16830 28590 16882
rect 28642 16830 28654 16882
rect 28914 16830 28926 16882
rect 28978 16830 28990 16882
rect 29542 16870 29554 16922
rect 29606 16870 29618 16922
rect 29698 16866 29710 16918
rect 29762 16866 29774 16918
rect 30146 16866 30158 16918
rect 30210 16866 30222 16918
rect 30482 16886 30494 16938
rect 30546 16886 30558 16938
rect 34414 16882 34466 16894
rect 27806 16818 27858 16830
rect 34414 16818 34466 16830
rect 34526 16882 34578 16894
rect 34526 16818 34578 16830
rect 34078 16770 34130 16782
rect 14466 16718 14478 16770
rect 14530 16718 14542 16770
rect 21634 16718 21646 16770
rect 21698 16718 21710 16770
rect 29038 16714 29090 16726
rect 29474 16718 29486 16770
rect 29538 16718 29550 16770
rect 35298 16718 35310 16770
rect 35362 16718 35374 16770
rect 37202 16718 37214 16770
rect 37266 16718 37278 16770
rect 34078 16706 34130 16718
rect 23930 16606 23942 16658
rect 23994 16606 24006 16658
rect 29038 16650 29090 16662
rect 1344 16490 38640 16524
rect 1344 16438 5876 16490
rect 5928 16438 5980 16490
rect 6032 16438 6084 16490
rect 6136 16438 15200 16490
rect 15252 16438 15304 16490
rect 15356 16438 15408 16490
rect 15460 16438 24524 16490
rect 24576 16438 24628 16490
rect 24680 16438 24732 16490
rect 24784 16438 33848 16490
rect 33900 16438 33952 16490
rect 34004 16438 34056 16490
rect 34108 16438 38640 16490
rect 1344 16404 38640 16438
rect 14478 16322 14530 16334
rect 14478 16258 14530 16270
rect 18398 16322 18450 16334
rect 18398 16258 18450 16270
rect 22224 16322 22276 16334
rect 19618 16214 19630 16266
rect 19682 16214 19694 16266
rect 22224 16258 22276 16270
rect 22766 16322 22818 16334
rect 22766 16258 22818 16270
rect 35068 16322 35120 16334
rect 37370 16270 37382 16322
rect 37434 16270 37446 16322
rect 35068 16258 35120 16270
rect 20638 16210 20690 16222
rect 20638 16146 20690 16158
rect 27414 16210 27466 16222
rect 31390 16210 31442 16222
rect 28354 16158 28366 16210
rect 28418 16158 28430 16210
rect 27414 16146 27466 16158
rect 31390 16146 31442 16158
rect 32006 16210 32058 16222
rect 32006 16146 32058 16158
rect 33798 16210 33850 16222
rect 33798 16146 33850 16158
rect 36486 16210 36538 16222
rect 36486 16146 36538 16158
rect 11342 16098 11394 16110
rect 11342 16034 11394 16046
rect 11734 16098 11786 16110
rect 11734 16034 11786 16046
rect 13358 16098 13410 16110
rect 13358 16034 13410 16046
rect 15374 16098 15426 16110
rect 15374 16034 15426 16046
rect 18062 16098 18114 16110
rect 18062 16034 18114 16046
rect 18846 16098 18898 16110
rect 21310 16098 21362 16110
rect 19506 16046 19518 16098
rect 19570 16046 19582 16098
rect 20402 16046 20414 16098
rect 20466 16046 20478 16098
rect 18846 16034 18898 16046
rect 20806 16042 20858 16054
rect 11006 15986 11058 15998
rect 20234 15990 20246 16042
rect 20298 15990 20310 16042
rect 21310 16034 21362 16046
rect 21982 16098 22034 16110
rect 21466 15990 21478 16042
rect 21530 15990 21542 16042
rect 21982 16034 22034 16046
rect 23102 16098 23154 16110
rect 25454 16098 25506 16110
rect 24565 16046 24577 16098
rect 24629 16046 24641 16098
rect 23102 16034 23154 16046
rect 25454 16034 25506 16046
rect 27918 16098 27970 16110
rect 30718 16098 30770 16110
rect 30996 16098 31048 16110
rect 28578 16046 28590 16098
rect 28642 16046 28654 16098
rect 27918 16034 27970 16046
rect 20806 15978 20858 15990
rect 24334 15986 24386 15998
rect 28242 15990 28254 16042
rect 28306 15990 28318 16042
rect 29318 16013 29330 16065
rect 29382 16013 29394 16065
rect 29474 16009 29486 16061
rect 29538 16009 29550 16061
rect 29922 16009 29934 16061
rect 29986 16009 29998 16061
rect 30370 16013 30382 16065
rect 30434 16013 30446 16065
rect 30818 16046 30830 16098
rect 30882 16046 30894 16098
rect 30718 16034 30770 16046
rect 30996 16034 31048 16046
rect 32846 16098 32898 16110
rect 32846 16034 32898 16046
rect 34526 16098 34578 16110
rect 34526 16034 34578 16046
rect 35310 16098 35362 16110
rect 35310 16034 35362 16046
rect 36878 16098 36930 16110
rect 11006 15922 11058 15934
rect 24334 15922 24386 15934
rect 29150 15986 29202 15998
rect 35802 15990 35814 16042
rect 35866 15990 35878 16042
rect 36878 16034 36930 16046
rect 37102 16098 37154 16110
rect 37102 16034 37154 16046
rect 29150 15922 29202 15934
rect 35982 15986 36034 15998
rect 35982 15922 36034 15934
rect 15710 15874 15762 15886
rect 15710 15810 15762 15822
rect 23494 15874 23546 15886
rect 23494 15810 23546 15822
rect 33182 15874 33234 15886
rect 33182 15810 33234 15822
rect 34190 15874 34242 15886
rect 34190 15810 34242 15822
rect 1344 15706 38800 15740
rect 1344 15654 10538 15706
rect 10590 15654 10642 15706
rect 10694 15654 10746 15706
rect 10798 15654 19862 15706
rect 19914 15654 19966 15706
rect 20018 15654 20070 15706
rect 20122 15654 29186 15706
rect 29238 15654 29290 15706
rect 29342 15654 29394 15706
rect 29446 15654 38510 15706
rect 38562 15654 38614 15706
rect 38666 15654 38718 15706
rect 38770 15654 38800 15706
rect 1344 15620 38800 15654
rect 12126 15538 12178 15550
rect 12126 15474 12178 15486
rect 15206 15538 15258 15550
rect 15206 15474 15258 15486
rect 23326 15538 23378 15550
rect 23326 15474 23378 15486
rect 23942 15538 23994 15550
rect 23942 15474 23994 15486
rect 25510 15538 25562 15550
rect 26002 15486 26014 15538
rect 26066 15535 26078 15538
rect 26338 15535 26350 15538
rect 26066 15489 26350 15535
rect 26066 15486 26078 15489
rect 26338 15486 26350 15489
rect 26402 15486 26414 15538
rect 25510 15474 25562 15486
rect 19966 15426 20018 15438
rect 19966 15362 20018 15374
rect 21758 15426 21810 15438
rect 21124 15352 21176 15364
rect 21758 15362 21810 15374
rect 22672 15426 22724 15438
rect 22672 15362 22724 15374
rect 27470 15426 27522 15438
rect 27470 15362 27522 15374
rect 31502 15426 31554 15438
rect 31502 15362 31554 15374
rect 33854 15426 33906 15438
rect 33854 15362 33906 15374
rect 35292 15426 35344 15438
rect 35292 15362 35344 15374
rect 36206 15426 36258 15438
rect 36206 15362 36258 15374
rect 12462 15314 12514 15326
rect 12462 15250 12514 15262
rect 17278 15314 17330 15326
rect 18050 15262 18062 15314
rect 18114 15262 18126 15314
rect 21422 15314 21474 15326
rect 21124 15288 21176 15300
rect 21298 15262 21310 15314
rect 21362 15262 21374 15314
rect 22430 15314 22482 15326
rect 17278 15250 17330 15262
rect 21422 15250 21474 15262
rect 21926 15258 21978 15270
rect 20750 15202 20802 15214
rect 22430 15250 22482 15262
rect 22990 15314 23042 15326
rect 28142 15314 28194 15326
rect 25330 15262 25342 15314
rect 25394 15262 25406 15314
rect 22990 15250 23042 15262
rect 27638 15258 27690 15270
rect 21926 15194 21978 15206
rect 24390 15202 24442 15214
rect 20750 15138 20802 15150
rect 28142 15250 28194 15262
rect 28814 15314 28866 15326
rect 34526 15314 34578 15326
rect 29586 15262 29598 15314
rect 29650 15262 29662 15314
rect 32946 15262 32958 15314
rect 33010 15262 33022 15314
rect 28814 15250 28866 15262
rect 34022 15258 34074 15270
rect 27638 15194 27690 15206
rect 32342 15202 32394 15214
rect 24390 15138 24442 15150
rect 34526 15250 34578 15262
rect 35534 15314 35586 15326
rect 35534 15250 35586 15262
rect 36038 15258 36090 15270
rect 34022 15194 34074 15206
rect 36038 15194 36090 15206
rect 32342 15138 32394 15150
rect 28384 15090 28436 15102
rect 28384 15026 28436 15038
rect 34768 15090 34820 15102
rect 34768 15026 34820 15038
rect 1344 14922 38640 14956
rect 1344 14870 5876 14922
rect 5928 14870 5980 14922
rect 6032 14870 6084 14922
rect 6136 14870 15200 14922
rect 15252 14870 15304 14922
rect 15356 14870 15408 14922
rect 15460 14870 24524 14922
rect 24576 14870 24628 14922
rect 24680 14870 24732 14922
rect 24784 14870 33848 14922
rect 33900 14870 33952 14922
rect 34004 14870 34056 14922
rect 34108 14870 38640 14922
rect 1344 14836 38640 14870
rect 13582 14754 13634 14766
rect 36336 14754 36388 14766
rect 11498 14702 11510 14754
rect 11562 14702 11574 14754
rect 20570 14702 20582 14754
rect 20634 14702 20646 14754
rect 13582 14690 13634 14702
rect 36336 14690 36388 14702
rect 12070 14642 12122 14654
rect 24502 14642 24554 14654
rect 17714 14590 17726 14642
rect 17778 14590 17790 14642
rect 19618 14590 19630 14642
rect 19682 14590 19694 14642
rect 12070 14578 12122 14590
rect 24502 14578 24554 14590
rect 27078 14642 27130 14654
rect 27078 14578 27130 14590
rect 29318 14642 29370 14654
rect 37158 14642 37210 14654
rect 33618 14590 33630 14642
rect 33682 14590 33694 14642
rect 29318 14578 29370 14590
rect 37158 14578 37210 14590
rect 7086 14530 7138 14542
rect 10894 14530 10946 14542
rect 7858 14478 7870 14530
rect 7922 14478 7934 14530
rect 7086 14466 7138 14478
rect 10894 14466 10946 14478
rect 11006 14530 11058 14542
rect 11006 14466 11058 14478
rect 11230 14530 11282 14542
rect 11230 14466 11282 14478
rect 13918 14530 13970 14542
rect 13918 14466 13970 14478
rect 16942 14530 16994 14542
rect 16942 14466 16994 14478
rect 20078 14530 20130 14542
rect 20078 14466 20130 14478
rect 20302 14530 20354 14542
rect 20302 14466 20354 14478
rect 21310 14530 21362 14542
rect 21310 14466 21362 14478
rect 21982 14530 22034 14542
rect 9774 14418 9826 14430
rect 21466 14422 21478 14474
rect 21530 14422 21542 14474
rect 21982 14466 22034 14478
rect 22224 14530 22276 14542
rect 23326 14530 23378 14542
rect 22642 14478 22654 14530
rect 22706 14478 22718 14530
rect 22224 14466 22276 14478
rect 23090 14422 23102 14474
rect 23154 14422 23166 14474
rect 23326 14466 23378 14478
rect 25118 14530 25170 14542
rect 25118 14466 25170 14478
rect 25342 14530 25394 14542
rect 25342 14466 25394 14478
rect 25902 14530 25954 14542
rect 25902 14466 25954 14478
rect 26574 14530 26626 14542
rect 25660 14418 25712 14430
rect 26394 14422 26406 14474
rect 26458 14422 26470 14474
rect 26574 14466 26626 14478
rect 28590 14530 28642 14542
rect 28590 14466 28642 14478
rect 31502 14530 31554 14542
rect 36094 14530 36146 14542
rect 31502 14466 31554 14478
rect 32610 14450 32622 14502
rect 32674 14450 32686 14502
rect 24826 14366 24838 14418
rect 24890 14366 24902 14418
rect 9774 14354 9826 14366
rect 10558 14306 10610 14318
rect 10558 14242 10610 14254
rect 14310 14306 14362 14318
rect 22754 14310 22766 14362
rect 22818 14310 22830 14362
rect 25660 14354 25712 14366
rect 35422 14418 35474 14430
rect 35578 14422 35590 14474
rect 35642 14422 35654 14474
rect 36094 14466 36146 14478
rect 38334 14530 38386 14542
rect 38334 14466 38386 14478
rect 35422 14354 35474 14366
rect 37998 14418 38050 14430
rect 37998 14354 38050 14366
rect 14310 14242 14362 14254
rect 24054 14306 24106 14318
rect 24054 14242 24106 14254
rect 28254 14306 28306 14318
rect 28254 14242 28306 14254
rect 31838 14306 31890 14318
rect 31838 14242 31890 14254
rect 37606 14306 37658 14318
rect 37606 14242 37658 14254
rect 1344 14138 38800 14172
rect 1344 14086 10538 14138
rect 10590 14086 10642 14138
rect 10694 14086 10746 14138
rect 10798 14086 19862 14138
rect 19914 14086 19966 14138
rect 20018 14086 20070 14138
rect 20122 14086 29186 14138
rect 29238 14086 29290 14138
rect 29342 14086 29394 14138
rect 29446 14086 38510 14138
rect 38562 14086 38614 14138
rect 38666 14086 38718 14138
rect 38770 14086 38800 14138
rect 1344 14052 38800 14086
rect 7982 13970 8034 13982
rect 7982 13906 8034 13918
rect 15094 13970 15146 13982
rect 15094 13906 15146 13918
rect 18006 13970 18058 13982
rect 18006 13906 18058 13918
rect 23942 13970 23994 13982
rect 23942 13906 23994 13918
rect 19630 13858 19682 13870
rect 19630 13794 19682 13806
rect 21310 13858 21362 13870
rect 21310 13794 21362 13806
rect 22318 13858 22370 13870
rect 22318 13794 22370 13806
rect 29934 13858 29986 13870
rect 29934 13794 29986 13806
rect 36300 13858 36352 13870
rect 36300 13794 36352 13806
rect 9102 13746 9154 13758
rect 9102 13682 9154 13694
rect 9998 13746 10050 13758
rect 10670 13746 10722 13758
rect 9998 13682 10050 13694
rect 10502 13690 10554 13702
rect 10670 13682 10722 13694
rect 14142 13746 14194 13758
rect 14142 13682 14194 13694
rect 16494 13746 16546 13758
rect 16494 13682 16546 13694
rect 18174 13746 18226 13758
rect 18174 13682 18226 13694
rect 20190 13746 20242 13758
rect 22990 13746 23042 13758
rect 20190 13682 20242 13694
rect 22486 13690 22538 13702
rect 10502 13626 10554 13638
rect 14534 13634 14586 13646
rect 11442 13582 11454 13634
rect 11506 13582 11518 13634
rect 13346 13582 13358 13634
rect 13410 13582 13422 13634
rect 22990 13682 23042 13694
rect 23232 13746 23284 13758
rect 25678 13746 25730 13758
rect 23762 13694 23774 13746
rect 23826 13694 23838 13746
rect 23232 13682 23284 13694
rect 25678 13682 25730 13694
rect 25790 13746 25842 13758
rect 25790 13682 25842 13694
rect 27246 13746 27298 13758
rect 31278 13746 31330 13758
rect 28018 13694 28030 13746
rect 28082 13694 28094 13746
rect 27246 13682 27298 13694
rect 31278 13682 31330 13694
rect 31390 13746 31442 13758
rect 31390 13682 31442 13694
rect 32174 13746 32226 13758
rect 32174 13682 32226 13694
rect 33070 13746 33122 13758
rect 35758 13746 35810 13758
rect 33842 13694 33854 13746
rect 33906 13694 33918 13746
rect 33070 13682 33122 13694
rect 35758 13682 35810 13694
rect 36542 13746 36594 13758
rect 37034 13750 37046 13802
rect 37098 13750 37110 13802
rect 36542 13682 36594 13694
rect 37214 13746 37266 13758
rect 37214 13682 37266 13694
rect 37438 13746 37490 13758
rect 37438 13682 37490 13694
rect 22486 13626 22538 13638
rect 24502 13634 24554 13646
rect 14534 13570 14586 13582
rect 24502 13570 24554 13582
rect 30662 13634 30714 13646
rect 30662 13570 30714 13582
rect 9756 13522 9808 13534
rect 9756 13458 9808 13470
rect 16158 13522 16210 13534
rect 16158 13458 16210 13470
rect 25342 13522 25394 13534
rect 25342 13458 25394 13470
rect 26126 13522 26178 13534
rect 31838 13522 31890 13534
rect 30986 13470 30998 13522
rect 31050 13470 31062 13522
rect 26126 13458 26178 13470
rect 31838 13458 31890 13470
rect 37774 13522 37826 13534
rect 37774 13458 37826 13470
rect 1344 13354 38640 13388
rect 1344 13302 5876 13354
rect 5928 13302 5980 13354
rect 6032 13302 6084 13354
rect 6136 13302 15200 13354
rect 15252 13302 15304 13354
rect 15356 13302 15408 13354
rect 15460 13302 24524 13354
rect 24576 13302 24628 13354
rect 24680 13302 24732 13354
rect 24784 13302 33848 13354
rect 33900 13302 33952 13354
rect 34004 13302 34056 13354
rect 34108 13302 38640 13354
rect 1344 13268 38640 13302
rect 12574 13186 12626 13198
rect 8586 13134 8598 13186
rect 8650 13134 8662 13186
rect 10490 13134 10502 13186
rect 10554 13134 10566 13186
rect 12574 13122 12626 13134
rect 19406 13186 19458 13198
rect 19406 13122 19458 13134
rect 22430 13186 22482 13198
rect 36362 13134 36374 13186
rect 36426 13134 36438 13186
rect 22430 13122 22482 13134
rect 13638 13074 13690 13086
rect 13638 13010 13690 13022
rect 14198 13074 14250 13086
rect 15810 13022 15822 13074
rect 15874 13022 15886 13074
rect 22866 13022 22878 13074
rect 22930 13022 22942 13074
rect 24322 13022 24334 13074
rect 24386 13022 24398 13074
rect 26226 13022 26238 13074
rect 26290 13022 26302 13074
rect 14198 13010 14250 13022
rect 8878 12962 8930 12974
rect 8878 12898 8930 12910
rect 9102 12962 9154 12974
rect 9102 12898 9154 12910
rect 10222 12962 10274 12974
rect 10222 12898 10274 12910
rect 10782 12962 10834 12974
rect 10782 12898 10834 12910
rect 11006 12962 11058 12974
rect 11006 12898 11058 12910
rect 11118 12962 11170 12974
rect 11118 12898 11170 12910
rect 14366 12962 14418 12974
rect 14366 12898 14418 12910
rect 15038 12962 15090 12974
rect 15038 12898 15090 12910
rect 17726 12962 17778 12974
rect 17726 12898 17778 12910
rect 20862 12962 20914 12974
rect 20862 12898 20914 12910
rect 21310 12962 21362 12974
rect 23550 12962 23602 12974
rect 29598 12962 29650 12974
rect 21310 12898 21362 12910
rect 18342 12850 18394 12862
rect 22174 12854 22186 12906
rect 22238 12854 22250 12906
rect 22978 12895 22990 12947
rect 23042 12895 23054 12947
rect 23202 12910 23214 12962
rect 23266 12910 23278 12962
rect 28690 12910 28702 12962
rect 28754 12910 28766 12962
rect 23550 12898 23602 12910
rect 29598 12898 29650 12910
rect 29934 12962 29986 12974
rect 29934 12898 29986 12910
rect 30046 12962 30098 12974
rect 33182 12962 33234 12974
rect 30818 12910 30830 12962
rect 30882 12910 30894 12962
rect 30046 12898 30098 12910
rect 33182 12898 33234 12910
rect 33854 12962 33906 12974
rect 18342 12786 18394 12798
rect 32734 12850 32786 12862
rect 33338 12854 33350 12906
rect 33402 12854 33414 12906
rect 33854 12898 33906 12910
rect 34638 12962 34690 12974
rect 34638 12898 34690 12910
rect 35310 12962 35362 12974
rect 32734 12786 32786 12798
rect 34096 12850 34148 12862
rect 34794 12854 34806 12906
rect 34858 12854 34870 12906
rect 35310 12898 35362 12910
rect 35552 12962 35604 12974
rect 35552 12898 35604 12910
rect 35870 12962 35922 12974
rect 35870 12898 35922 12910
rect 36094 12962 36146 12974
rect 36094 12898 36146 12910
rect 36990 12962 37042 12974
rect 36990 12898 37042 12910
rect 37158 12962 37210 12974
rect 37158 12898 37210 12910
rect 37662 12962 37714 12974
rect 37662 12898 37714 12910
rect 34096 12786 34148 12798
rect 37904 12850 37956 12862
rect 37904 12786 37956 12798
rect 7814 12738 7866 12750
rect 7814 12674 7866 12686
rect 9550 12738 9602 12750
rect 9550 12674 9602 12686
rect 14702 12738 14754 12750
rect 14702 12674 14754 12686
rect 1344 12570 38800 12604
rect 1344 12518 10538 12570
rect 10590 12518 10642 12570
rect 10694 12518 10746 12570
rect 10798 12518 19862 12570
rect 19914 12518 19966 12570
rect 20018 12518 20070 12570
rect 20122 12518 29186 12570
rect 29238 12518 29290 12570
rect 29342 12518 29394 12570
rect 29446 12518 38510 12570
rect 38562 12518 38614 12570
rect 38666 12518 38718 12570
rect 38770 12518 38800 12570
rect 1344 12484 38800 12518
rect 7310 12402 7362 12414
rect 7310 12338 7362 12350
rect 15094 12402 15146 12414
rect 10670 12290 10722 12302
rect 11890 12294 11902 12346
rect 11954 12294 11966 12346
rect 15094 12338 15146 12350
rect 22934 12402 22986 12414
rect 22934 12338 22986 12350
rect 23382 12402 23434 12414
rect 23382 12338 23434 12350
rect 33910 12402 33962 12414
rect 33910 12338 33962 12350
rect 35254 12402 35306 12414
rect 35254 12338 35306 12350
rect 18062 12290 18114 12302
rect 16202 12238 16214 12290
rect 16266 12238 16278 12290
rect 10670 12226 10722 12238
rect 18062 12226 18114 12238
rect 22318 12290 22370 12302
rect 22318 12226 22370 12238
rect 27806 12290 27858 12302
rect 27806 12226 27858 12238
rect 31166 12290 31218 12302
rect 31166 12226 31218 12238
rect 32080 12290 32132 12302
rect 35646 12290 35698 12302
rect 34234 12238 34246 12290
rect 34298 12238 34310 12290
rect 32080 12226 32132 12238
rect 35646 12226 35698 12238
rect 7646 12178 7698 12190
rect 7646 12114 7698 12126
rect 7870 12178 7922 12190
rect 7870 12114 7922 12126
rect 8038 12178 8090 12190
rect 8038 12114 8090 12126
rect 8542 12178 8594 12190
rect 9886 12178 9938 12190
rect 9594 12126 9606 12178
rect 9658 12126 9670 12178
rect 8542 12114 8594 12126
rect 9886 12114 9938 12126
rect 9998 12178 10050 12190
rect 9998 12114 10050 12126
rect 11006 12178 11058 12190
rect 11006 12114 11058 12126
rect 11566 12178 11618 12190
rect 11566 12114 11618 12126
rect 12070 12178 12122 12190
rect 12070 12114 12122 12126
rect 13806 12178 13858 12190
rect 14366 12178 14418 12190
rect 14074 12126 14086 12178
rect 14138 12126 14150 12178
rect 13806 12114 13858 12126
rect 14366 12114 14418 12126
rect 14590 12178 14642 12190
rect 16494 12178 16546 12190
rect 15250 12126 15262 12178
rect 15314 12126 15326 12178
rect 14590 12114 14642 12126
rect 16494 12114 16546 12126
rect 16718 12178 16770 12190
rect 16718 12114 16770 12126
rect 19182 12178 19234 12190
rect 19182 12114 19234 12126
rect 19630 12178 19682 12190
rect 25118 12178 25170 12190
rect 20402 12126 20414 12178
rect 20466 12126 20478 12178
rect 25890 12126 25902 12178
rect 25954 12126 25966 12178
rect 28578 12153 28590 12205
rect 28642 12153 28654 12205
rect 31838 12178 31890 12190
rect 19630 12114 19682 12126
rect 25118 12114 25170 12126
rect 31334 12122 31386 12134
rect 11324 12066 11376 12078
rect 11324 12002 11376 12014
rect 12742 12066 12794 12078
rect 12742 12002 12794 12014
rect 13134 12066 13186 12078
rect 31838 12114 31890 12126
rect 34526 12178 34578 12190
rect 34526 12114 34578 12126
rect 34638 12178 34690 12190
rect 38334 12178 38386 12190
rect 37538 12126 37550 12178
rect 37602 12126 37614 12178
rect 34638 12114 34690 12126
rect 38334 12114 38386 12126
rect 31334 12058 31386 12070
rect 13134 12002 13186 12014
rect 8784 11954 8836 11966
rect 8784 11890 8836 11902
rect 29374 11954 29426 11966
rect 29374 11890 29426 11902
rect 1344 11786 38640 11820
rect 1344 11734 5876 11786
rect 5928 11734 5980 11786
rect 6032 11734 6084 11786
rect 6136 11734 15200 11786
rect 15252 11734 15304 11786
rect 15356 11734 15408 11786
rect 15460 11734 24524 11786
rect 24576 11734 24628 11786
rect 24680 11734 24732 11786
rect 24784 11734 33848 11786
rect 33900 11734 33952 11786
rect 34004 11734 34056 11786
rect 34108 11734 38640 11786
rect 1344 11700 38640 11734
rect 22430 11618 22482 11630
rect 22430 11554 22482 11566
rect 37998 11618 38050 11630
rect 37998 11554 38050 11566
rect 17670 11506 17722 11518
rect 14578 11454 14590 11506
rect 14642 11454 14654 11506
rect 17670 11442 17722 11454
rect 23046 11506 23098 11518
rect 23046 11442 23098 11454
rect 28086 11506 28138 11518
rect 28086 11442 28138 11454
rect 5854 11394 5906 11406
rect 9326 11394 9378 11406
rect 6626 11342 6638 11394
rect 6690 11342 6702 11394
rect 5854 11330 5906 11342
rect 9326 11330 9378 11342
rect 9438 11394 9490 11406
rect 9438 11330 9490 11342
rect 9998 11394 10050 11406
rect 9998 11330 10050 11342
rect 10110 11394 10162 11406
rect 11902 11394 11954 11406
rect 10378 11342 10390 11394
rect 10442 11342 10454 11394
rect 10658 11342 10670 11394
rect 10722 11342 10734 11394
rect 10110 11330 10162 11342
rect 11902 11330 11954 11342
rect 12070 11394 12122 11406
rect 12070 11330 12122 11342
rect 12574 11394 12626 11406
rect 12574 11330 12626 11342
rect 12816 11394 12868 11406
rect 12816 11330 12868 11342
rect 14030 11394 14082 11406
rect 14030 11330 14082 11342
rect 14142 11394 14194 11406
rect 17278 11394 17330 11406
rect 16482 11342 16494 11394
rect 16546 11342 16558 11394
rect 14142 11330 14194 11342
rect 17278 11330 17330 11342
rect 17950 11394 18002 11406
rect 20638 11394 20690 11406
rect 18722 11342 18734 11394
rect 18786 11342 18798 11394
rect 17950 11330 18002 11342
rect 20638 11330 20690 11342
rect 21310 11394 21362 11406
rect 26350 11394 26402 11406
rect 22174 11342 22186 11394
rect 22238 11342 22250 11394
rect 21310 11330 21362 11342
rect 26350 11330 26402 11342
rect 26574 11394 26626 11406
rect 26574 11330 26626 11342
rect 27246 11394 27298 11406
rect 27246 11330 27298 11342
rect 30046 11394 30098 11406
rect 30046 11330 30098 11342
rect 30158 11394 30210 11406
rect 30158 11330 30210 11342
rect 38334 11394 38386 11406
rect 38334 11330 38386 11342
rect 8542 11282 8594 11294
rect 37606 11282 37658 11294
rect 9034 11230 9046 11282
rect 9098 11230 9110 11282
rect 13738 11230 13750 11282
rect 13802 11230 13814 11282
rect 26058 11230 26070 11282
rect 26122 11230 26134 11282
rect 8542 11218 8594 11230
rect 37606 11218 37658 11230
rect 26910 11170 26962 11182
rect 26910 11106 26962 11118
rect 29710 11170 29762 11182
rect 29710 11106 29762 11118
rect 30494 11170 30546 11182
rect 30494 11106 30546 11118
rect 35254 11170 35306 11182
rect 35254 11106 35306 11118
rect 1344 11002 38800 11036
rect 1344 10950 10538 11002
rect 10590 10950 10642 11002
rect 10694 10950 10746 11002
rect 10798 10950 19862 11002
rect 19914 10950 19966 11002
rect 20018 10950 20070 11002
rect 20122 10950 29186 11002
rect 29238 10950 29290 11002
rect 29342 10950 29394 11002
rect 29446 10950 38510 11002
rect 38562 10950 38614 11002
rect 38666 10950 38718 11002
rect 38770 10950 38800 11002
rect 1344 10916 38800 10950
rect 6526 10834 6578 10846
rect 6526 10770 6578 10782
rect 12238 10834 12290 10846
rect 12238 10770 12290 10782
rect 15822 10834 15874 10846
rect 15822 10770 15874 10782
rect 17558 10834 17610 10846
rect 17558 10770 17610 10782
rect 18902 10834 18954 10846
rect 18902 10770 18954 10782
rect 21030 10834 21082 10846
rect 21030 10770 21082 10782
rect 37270 10834 37322 10846
rect 37270 10770 37322 10782
rect 9550 10722 9602 10734
rect 30848 10722 30900 10734
rect 29530 10670 29542 10722
rect 29594 10670 29606 10722
rect 9550 10658 9602 10670
rect 30848 10658 30900 10670
rect 36654 10722 36706 10734
rect 36654 10658 36706 10670
rect 7982 10610 8034 10622
rect 7982 10546 8034 10558
rect 8430 10610 8482 10622
rect 8430 10546 8482 10558
rect 8654 10610 8706 10622
rect 10222 10610 10274 10622
rect 8654 10546 8706 10558
rect 9718 10554 9770 10566
rect 11218 10585 11230 10637
rect 11282 10585 11294 10637
rect 14254 10610 14306 10622
rect 10222 10546 10274 10558
rect 14254 10546 14306 10558
rect 14366 10610 14418 10622
rect 14366 10546 14418 10558
rect 19294 10610 19346 10622
rect 19294 10546 19346 10558
rect 19630 10610 19682 10622
rect 19630 10546 19682 10558
rect 19742 10610 19794 10622
rect 19742 10546 19794 10558
rect 23886 10610 23938 10622
rect 23886 10546 23938 10558
rect 25118 10610 25170 10622
rect 28702 10610 28754 10622
rect 25890 10558 25902 10610
rect 25954 10558 25966 10610
rect 25118 10546 25170 10558
rect 28702 10546 28754 10558
rect 29150 10610 29202 10622
rect 29150 10546 29202 10558
rect 29262 10610 29314 10622
rect 29262 10546 29314 10558
rect 29934 10610 29986 10622
rect 30606 10610 30658 10622
rect 29934 10546 29986 10558
rect 30102 10554 30154 10566
rect 9718 10490 9770 10502
rect 30606 10546 30658 10558
rect 33966 10610 34018 10622
rect 33966 10546 34018 10558
rect 27794 10446 27806 10498
rect 27858 10446 27870 10498
rect 30102 10490 30154 10502
rect 34738 10446 34750 10498
rect 34802 10446 34814 10498
rect 10464 10386 10516 10398
rect 8922 10334 8934 10386
rect 8986 10334 8998 10386
rect 10464 10322 10516 10334
rect 13918 10386 13970 10398
rect 13918 10322 13970 10334
rect 20078 10386 20130 10398
rect 20078 10322 20130 10334
rect 23550 10386 23602 10398
rect 23550 10322 23602 10334
rect 28366 10386 28418 10398
rect 28366 10322 28418 10334
rect 1344 10218 38640 10252
rect 1344 10166 5876 10218
rect 5928 10166 5980 10218
rect 6032 10166 6084 10218
rect 6136 10166 15200 10218
rect 15252 10166 15304 10218
rect 15356 10166 15408 10218
rect 15460 10166 24524 10218
rect 24576 10166 24628 10218
rect 24680 10166 24732 10218
rect 24784 10166 33848 10218
rect 33900 10166 33952 10218
rect 34004 10166 34056 10218
rect 34108 10166 38640 10218
rect 1344 10132 38640 10166
rect 34862 10050 34914 10062
rect 34862 9986 34914 9998
rect 10166 9938 10218 9950
rect 10166 9874 10218 9886
rect 12966 9938 13018 9950
rect 12966 9874 13018 9886
rect 14422 9938 14474 9950
rect 14422 9874 14474 9886
rect 14870 9938 14922 9950
rect 14870 9874 14922 9886
rect 20470 9938 20522 9950
rect 23202 9886 23214 9938
rect 23266 9886 23278 9938
rect 20470 9874 20522 9886
rect 26630 9882 26682 9894
rect 5518 9826 5570 9838
rect 8990 9826 9042 9838
rect 6290 9774 6302 9826
rect 6354 9774 6366 9826
rect 5518 9762 5570 9774
rect 8990 9762 9042 9774
rect 9662 9826 9714 9838
rect 8206 9714 8258 9726
rect 8206 9650 8258 9662
rect 8748 9714 8800 9726
rect 9482 9718 9494 9770
rect 9546 9718 9558 9770
rect 9662 9762 9714 9774
rect 10446 9826 10498 9838
rect 10446 9762 10498 9774
rect 13806 9826 13858 9838
rect 13806 9762 13858 9774
rect 13918 9826 13970 9838
rect 17502 9826 17554 9838
rect 13918 9762 13970 9774
rect 15474 9746 15486 9798
rect 15538 9746 15550 9798
rect 17502 9762 17554 9774
rect 20078 9826 20130 9838
rect 20078 9762 20130 9774
rect 22430 9826 22482 9838
rect 22430 9762 22482 9774
rect 25118 9826 25170 9838
rect 25118 9762 25170 9774
rect 26126 9826 26178 9838
rect 26630 9818 26682 9830
rect 27302 9882 27354 9894
rect 29250 9886 29262 9938
rect 29314 9886 29326 9938
rect 31154 9886 31166 9938
rect 31218 9886 31230 9938
rect 27302 9818 27354 9830
rect 27806 9826 27858 9838
rect 26126 9762 26178 9774
rect 27806 9762 27858 9774
rect 31950 9826 32002 9838
rect 31950 9762 32002 9774
rect 32622 9826 32674 9838
rect 32622 9762 32674 9774
rect 32846 9826 32898 9838
rect 33406 9826 33458 9838
rect 33114 9774 33126 9826
rect 33178 9774 33190 9826
rect 32846 9762 32898 9774
rect 33406 9762 33458 9774
rect 37662 9826 37714 9838
rect 25884 9714 25936 9726
rect 13514 9662 13526 9714
rect 13578 9662 13590 9714
rect 8748 9650 8800 9662
rect 25884 9650 25936 9662
rect 26798 9714 26850 9726
rect 26798 9650 26850 9662
rect 27134 9714 27186 9726
rect 27134 9650 27186 9662
rect 28048 9714 28100 9726
rect 37146 9718 37158 9770
rect 37210 9718 37222 9770
rect 37662 9762 37714 9774
rect 37904 9826 37956 9838
rect 37904 9762 37956 9774
rect 28048 9650 28100 9662
rect 11566 9602 11618 9614
rect 11566 9538 11618 9550
rect 18958 9602 19010 9614
rect 18958 9538 19010 9550
rect 32342 9602 32394 9614
rect 37314 9606 37326 9658
rect 37378 9606 37390 9658
rect 32342 9538 32394 9550
rect 1344 9434 38800 9468
rect 1344 9382 10538 9434
rect 10590 9382 10642 9434
rect 10694 9382 10746 9434
rect 10798 9382 19862 9434
rect 19914 9382 19966 9434
rect 20018 9382 20070 9434
rect 20122 9382 29186 9434
rect 29238 9382 29290 9434
rect 29342 9382 29394 9434
rect 29446 9382 38510 9434
rect 38562 9382 38614 9434
rect 38666 9382 38718 9434
rect 38770 9382 38800 9434
rect 1344 9348 38800 9382
rect 5966 9266 6018 9278
rect 5966 9202 6018 9214
rect 17558 9266 17610 9278
rect 17558 9202 17610 9214
rect 18230 9266 18282 9278
rect 18230 9202 18282 9214
rect 35254 9266 35306 9278
rect 9774 9154 9826 9166
rect 26562 9158 26574 9210
rect 26626 9158 26638 9210
rect 35254 9202 35306 9214
rect 29038 9154 29090 9166
rect 8922 9102 8934 9154
rect 8986 9102 8998 9154
rect 27290 9102 27302 9154
rect 27354 9102 27366 9154
rect 9774 9090 9826 9102
rect 29038 9090 29090 9102
rect 29468 9154 29520 9166
rect 29468 9090 29520 9102
rect 30382 9154 30434 9166
rect 30382 9090 30434 9102
rect 7086 9042 7138 9054
rect 8094 9042 8146 9054
rect 7802 8990 7814 9042
rect 7866 8990 7878 9042
rect 7086 8978 7138 8990
rect 8094 8978 8146 8990
rect 8318 9042 8370 9054
rect 8318 8978 8370 8990
rect 8430 9042 8482 9054
rect 8430 8978 8482 8990
rect 8654 9042 8706 9054
rect 12462 9042 12514 9054
rect 11666 8990 11678 9042
rect 11730 8990 11742 9042
rect 8654 8978 8706 8990
rect 12462 8978 12514 8990
rect 12798 9042 12850 9054
rect 12798 8978 12850 8990
rect 16942 9042 16994 9054
rect 16942 8978 16994 8990
rect 20638 9042 20690 9054
rect 20638 8978 20690 8990
rect 26238 9042 26290 9054
rect 27582 9042 27634 9054
rect 26238 8978 26290 8990
rect 26742 8986 26794 8998
rect 27582 8978 27634 8990
rect 27806 9042 27858 9054
rect 27806 8978 27858 8990
rect 28124 9042 28176 9054
rect 28124 8978 28176 8990
rect 28366 9042 28418 9054
rect 29710 9042 29762 9054
rect 28366 8978 28418 8990
rect 28870 8986 28922 8998
rect 26742 8922 26794 8934
rect 29710 8978 29762 8990
rect 30214 9042 30266 9054
rect 30214 8978 30266 8990
rect 30718 9042 30770 9054
rect 30718 8978 30770 8990
rect 38334 9042 38386 9054
rect 38334 8978 38386 8990
rect 28870 8922 28922 8934
rect 35634 8878 35646 8930
rect 35698 8878 35710 8930
rect 37538 8878 37550 8930
rect 37602 8878 37614 8930
rect 14254 8818 14306 8830
rect 14254 8754 14306 8766
rect 15822 8818 15874 8830
rect 15822 8754 15874 8766
rect 19182 8818 19234 8830
rect 19182 8754 19234 8766
rect 25996 8818 26048 8830
rect 25996 8754 26048 8766
rect 32174 8818 32226 8830
rect 32174 8754 32226 8766
rect 1344 8650 38640 8684
rect 1344 8598 5876 8650
rect 5928 8598 5980 8650
rect 6032 8598 6084 8650
rect 6136 8598 15200 8650
rect 15252 8598 15304 8650
rect 15356 8598 15408 8650
rect 15460 8598 24524 8650
rect 24576 8598 24628 8650
rect 24680 8598 24732 8650
rect 24784 8598 33848 8650
rect 33900 8598 33952 8650
rect 34004 8598 34056 8650
rect 34108 8598 38640 8650
rect 1344 8564 38640 8598
rect 13564 8482 13616 8494
rect 11498 8430 11510 8482
rect 11562 8430 11574 8482
rect 13564 8418 13616 8430
rect 8560 8370 8612 8382
rect 14982 8370 15034 8382
rect 36000 8370 36052 8382
rect 8560 8306 8612 8318
rect 14310 8314 14362 8326
rect 7646 8258 7698 8270
rect 7646 8194 7698 8206
rect 8318 8258 8370 8270
rect 7802 8150 7814 8202
rect 7866 8150 7878 8202
rect 8318 8194 8370 8206
rect 9326 8258 9378 8270
rect 9326 8194 9378 8206
rect 9438 8258 9490 8270
rect 9438 8194 9490 8206
rect 11790 8258 11842 8270
rect 11790 8194 11842 8206
rect 12014 8258 12066 8270
rect 12014 8194 12066 8206
rect 13806 8258 13858 8270
rect 18722 8318 18734 8370
rect 18786 8318 18798 8370
rect 26058 8318 26070 8370
rect 26122 8318 26134 8370
rect 14982 8306 15034 8318
rect 36000 8306 36052 8318
rect 37904 8370 37956 8382
rect 37904 8306 37956 8318
rect 14310 8250 14362 8262
rect 17950 8258 18002 8270
rect 13806 8194 13858 8206
rect 17950 8194 18002 8206
rect 22206 8258 22258 8270
rect 22206 8194 22258 8206
rect 23326 8258 23378 8270
rect 23326 8194 23378 8206
rect 23550 8258 23602 8270
rect 23550 8194 23602 8206
rect 26350 8258 26402 8270
rect 26350 8194 26402 8206
rect 26462 8258 26514 8270
rect 26462 8194 26514 8206
rect 27134 8258 27186 8270
rect 27134 8194 27186 8206
rect 27246 8258 27298 8270
rect 27246 8194 27298 8206
rect 29038 8258 29090 8270
rect 29038 8194 29090 8206
rect 32062 8258 32114 8270
rect 32062 8194 32114 8206
rect 32174 8258 32226 8270
rect 32174 8194 32226 8206
rect 34190 8258 34242 8270
rect 34190 8194 34242 8206
rect 34414 8258 34466 8270
rect 34414 8194 34466 8206
rect 35758 8258 35810 8270
rect 14478 8146 14530 8158
rect 9034 8094 9046 8146
rect 9098 8094 9110 8146
rect 14478 8082 14530 8094
rect 20638 8146 20690 8158
rect 35086 8146 35138 8158
rect 35242 8150 35254 8202
rect 35306 8150 35318 8202
rect 35758 8194 35810 8206
rect 37662 8258 37714 8270
rect 23034 8094 23046 8146
rect 23098 8094 23110 8146
rect 26842 8094 26854 8146
rect 26906 8094 26918 8146
rect 34682 8094 34694 8146
rect 34746 8094 34758 8146
rect 20638 8082 20690 8094
rect 35086 8082 35138 8094
rect 36990 8146 37042 8158
rect 37146 8150 37158 8202
rect 37210 8150 37222 8202
rect 37662 8194 37714 8206
rect 36990 8082 37042 8094
rect 9942 8034 9994 8046
rect 9942 7970 9994 7982
rect 17110 8034 17162 8046
rect 17110 7970 17162 7982
rect 17782 8034 17834 8046
rect 17782 7970 17834 7982
rect 22542 8034 22594 8046
rect 22542 7970 22594 7982
rect 29374 8034 29426 8046
rect 29374 7970 29426 7982
rect 30606 8034 30658 8046
rect 30606 7970 30658 7982
rect 32510 8034 32562 8046
rect 32510 7970 32562 7982
rect 1344 7866 38800 7900
rect 1344 7814 10538 7866
rect 10590 7814 10642 7866
rect 10694 7814 10746 7866
rect 10798 7814 19862 7866
rect 19914 7814 19966 7866
rect 20018 7814 20070 7866
rect 20122 7814 29186 7866
rect 29238 7814 29290 7866
rect 29342 7814 29394 7866
rect 29446 7814 38510 7866
rect 38562 7814 38614 7866
rect 38666 7814 38718 7866
rect 38770 7814 38800 7866
rect 1344 7780 38800 7814
rect 11062 7698 11114 7710
rect 11062 7634 11114 7646
rect 36654 7698 36706 7710
rect 7982 7586 8034 7598
rect 7578 7534 7590 7586
rect 7642 7534 7654 7586
rect 7982 7522 8034 7534
rect 12462 7586 12514 7598
rect 12462 7522 12514 7534
rect 25436 7586 25488 7598
rect 25436 7522 25488 7534
rect 26350 7586 26402 7598
rect 27010 7590 27022 7642
rect 27074 7590 27086 7642
rect 36654 7634 36706 7646
rect 37998 7698 38050 7710
rect 37998 7634 38050 7646
rect 7086 7474 7138 7486
rect 7086 7410 7138 7422
rect 7310 7474 7362 7486
rect 7310 7410 7362 7422
rect 8150 7474 8202 7486
rect 8150 7410 8202 7422
rect 8654 7474 8706 7486
rect 8654 7410 8706 7422
rect 9438 7474 9490 7486
rect 9438 7410 9490 7422
rect 9662 7474 9714 7486
rect 11902 7474 11954 7486
rect 9930 7422 9942 7474
rect 9994 7422 10006 7474
rect 9662 7410 9714 7422
rect 11902 7410 11954 7422
rect 12126 7474 12178 7486
rect 15150 7474 15202 7486
rect 14354 7422 14366 7474
rect 14418 7422 14430 7474
rect 12126 7410 12178 7422
rect 15150 7410 15202 7422
rect 16718 7474 16770 7486
rect 16718 7410 16770 7422
rect 16942 7474 16994 7486
rect 16942 7410 16994 7422
rect 17278 7474 17330 7486
rect 17278 7410 17330 7422
rect 20750 7474 20802 7486
rect 21422 7474 21474 7486
rect 20750 7410 20802 7422
rect 21254 7418 21306 7430
rect 15542 7362 15594 7374
rect 21422 7410 21474 7422
rect 21870 7474 21922 7486
rect 21870 7410 21922 7422
rect 24558 7474 24610 7486
rect 24558 7410 24610 7422
rect 25678 7474 25730 7486
rect 26170 7478 26182 7530
rect 26234 7478 26246 7530
rect 26350 7522 26402 7534
rect 29038 7586 29090 7598
rect 29038 7522 29090 7534
rect 35216 7586 35268 7598
rect 35216 7522 35268 7534
rect 27358 7474 27410 7486
rect 25678 7410 25730 7422
rect 26854 7418 26906 7430
rect 18050 7310 18062 7362
rect 18114 7310 18126 7362
rect 19954 7310 19966 7362
rect 20018 7310 20030 7362
rect 21254 7354 21306 7366
rect 27358 7410 27410 7422
rect 28366 7474 28418 7486
rect 30942 7474 30994 7486
rect 28366 7410 28418 7422
rect 28870 7418 28922 7430
rect 22642 7310 22654 7362
rect 22706 7310 22718 7362
rect 26854 7354 26906 7366
rect 30942 7410 30994 7422
rect 34302 7474 34354 7486
rect 34974 7474 35026 7486
rect 34302 7410 34354 7422
rect 34470 7418 34522 7430
rect 28870 7354 28922 7366
rect 34974 7410 35026 7422
rect 35534 7474 35586 7486
rect 35534 7410 35586 7422
rect 38334 7474 38386 7486
rect 38334 7410 38386 7422
rect 34470 7354 34522 7366
rect 15542 7298 15594 7310
rect 8896 7250 8948 7262
rect 20508 7250 20560 7262
rect 11610 7198 11622 7250
rect 11674 7198 11686 7250
rect 16426 7198 16438 7250
rect 16490 7198 16502 7250
rect 8896 7186 8948 7198
rect 20508 7186 20560 7198
rect 27600 7250 27652 7262
rect 27600 7186 27652 7198
rect 28124 7250 28176 7262
rect 28124 7186 28176 7198
rect 30606 7250 30658 7262
rect 30606 7186 30658 7198
rect 1344 7082 38640 7116
rect 1344 7030 5876 7082
rect 5928 7030 5980 7082
rect 6032 7030 6084 7082
rect 6136 7030 15200 7082
rect 15252 7030 15304 7082
rect 15356 7030 15408 7082
rect 15460 7030 24524 7082
rect 24576 7030 24628 7082
rect 24680 7030 24732 7082
rect 24784 7030 33848 7082
rect 33900 7030 33952 7082
rect 34004 7030 34056 7082
rect 34108 7030 38640 7082
rect 1344 6996 38640 7030
rect 15356 6914 15408 6926
rect 15356 6850 15408 6862
rect 17950 6914 18002 6926
rect 17950 6850 18002 6862
rect 22542 6914 22594 6926
rect 22542 6850 22594 6862
rect 19014 6746 19066 6758
rect 8094 6690 8146 6702
rect 8094 6626 8146 6638
rect 10110 6690 10162 6702
rect 10670 6690 10722 6702
rect 10378 6638 10390 6690
rect 10442 6638 10454 6690
rect 10110 6626 10162 6638
rect 10670 6626 10722 6638
rect 10782 6690 10834 6702
rect 10782 6626 10834 6638
rect 11118 6690 11170 6702
rect 11118 6626 11170 6638
rect 13806 6690 13858 6702
rect 13806 6626 13858 6638
rect 15598 6690 15650 6702
rect 13564 6578 13616 6590
rect 14298 6582 14310 6634
rect 14362 6582 14374 6634
rect 15598 6626 15650 6638
rect 16270 6690 16322 6702
rect 13564 6514 13616 6526
rect 14478 6578 14530 6590
rect 16090 6582 16102 6634
rect 16154 6582 16166 6634
rect 16270 6626 16322 6638
rect 16494 6690 16546 6702
rect 16494 6626 16546 6638
rect 18846 6690 18898 6702
rect 19014 6682 19066 6694
rect 19518 6690 19570 6702
rect 18846 6626 18898 6638
rect 19518 6626 19570 6638
rect 19760 6690 19812 6702
rect 19760 6626 19812 6638
rect 20078 6690 20130 6702
rect 20078 6626 20130 6638
rect 20302 6690 20354 6702
rect 21758 6690 21810 6702
rect 20570 6638 20582 6690
rect 20634 6638 20646 6690
rect 20302 6626 20354 6638
rect 21758 6626 21810 6638
rect 23998 6690 24050 6702
rect 23998 6626 24050 6638
rect 24670 6690 24722 6702
rect 24670 6626 24722 6638
rect 26686 6690 26738 6702
rect 26686 6626 26738 6638
rect 29486 6690 29538 6702
rect 29486 6626 29538 6638
rect 29654 6690 29706 6702
rect 29654 6626 29706 6638
rect 30158 6690 30210 6702
rect 30158 6626 30210 6638
rect 30718 6690 30770 6702
rect 30718 6626 30770 6638
rect 30942 6690 30994 6702
rect 30942 6626 30994 6638
rect 33294 6690 33346 6702
rect 33294 6626 33346 6638
rect 33966 6690 34018 6702
rect 14478 6514 14530 6526
rect 30400 6578 30452 6590
rect 33450 6582 33462 6634
rect 33514 6582 33526 6634
rect 33966 6626 34018 6638
rect 34638 6690 34690 6702
rect 34638 6626 34690 6638
rect 36990 6690 37042 6702
rect 36990 6626 37042 6638
rect 37662 6690 37714 6702
rect 34208 6578 34260 6590
rect 37146 6582 37158 6634
rect 37210 6582 37222 6634
rect 37662 6626 37714 6638
rect 31210 6526 31222 6578
rect 31274 6526 31286 6578
rect 30400 6514 30452 6526
rect 34208 6514 34260 6526
rect 37904 6578 37956 6590
rect 37904 6514 37956 6526
rect 6638 6466 6690 6478
rect 6638 6402 6690 6414
rect 8990 6466 9042 6478
rect 8990 6402 9042 6414
rect 12238 6466 12290 6478
rect 12238 6402 12290 6414
rect 21422 6466 21474 6478
rect 21422 6402 21474 6414
rect 25790 6466 25842 6478
rect 25790 6402 25842 6414
rect 27806 6466 27858 6478
rect 27806 6402 27858 6414
rect 36094 6466 36146 6478
rect 36094 6402 36146 6414
rect 1344 6298 38800 6332
rect 1344 6246 10538 6298
rect 10590 6246 10642 6298
rect 10694 6246 10746 6298
rect 10798 6246 19862 6298
rect 19914 6246 19966 6298
rect 20018 6246 20070 6298
rect 20122 6246 29186 6298
rect 29238 6246 29290 6298
rect 29342 6246 29394 6298
rect 29446 6246 38510 6298
rect 38562 6246 38614 6298
rect 38666 6246 38718 6298
rect 38770 6246 38800 6298
rect 1344 6212 38800 6246
rect 8542 6018 8594 6030
rect 9986 6022 9998 6074
rect 10050 6022 10062 6074
rect 8542 5954 8594 5966
rect 10688 6018 10740 6030
rect 10688 5954 10740 5966
rect 13694 6018 13746 6030
rect 13694 5954 13746 5966
rect 21422 6018 21474 6030
rect 29468 6018 29520 6030
rect 30034 6022 30046 6074
rect 30098 6022 30110 6074
rect 24602 5966 24614 6018
rect 24666 5966 24678 6018
rect 21422 5954 21474 5966
rect 5854 5906 5906 5918
rect 9942 5906 9994 5918
rect 6626 5854 6638 5906
rect 6690 5854 6702 5906
rect 5854 5842 5906 5854
rect 9942 5842 9994 5854
rect 10446 5906 10498 5918
rect 10446 5842 10498 5854
rect 11006 5906 11058 5918
rect 11778 5854 11790 5906
rect 11842 5854 11854 5906
rect 14130 5881 14142 5933
rect 14194 5881 14206 5933
rect 17490 5881 17502 5933
rect 17554 5881 17566 5933
rect 20302 5906 20354 5918
rect 11006 5842 11058 5854
rect 20302 5842 20354 5854
rect 20414 5906 20466 5918
rect 20414 5842 20466 5854
rect 21590 5906 21642 5918
rect 21590 5842 21642 5854
rect 22094 5906 22146 5918
rect 22094 5842 22146 5854
rect 22766 5906 22818 5918
rect 22766 5842 22818 5854
rect 22878 5906 22930 5918
rect 22878 5842 22930 5854
rect 24110 5906 24162 5918
rect 24110 5842 24162 5854
rect 24334 5906 24386 5918
rect 25218 5881 25230 5933
rect 25282 5881 25294 5933
rect 28124 5906 28176 5918
rect 24334 5842 24386 5854
rect 28124 5842 28176 5854
rect 28366 5906 28418 5918
rect 28858 5910 28870 5962
rect 28922 5910 28934 5962
rect 29468 5954 29520 5966
rect 30718 6018 30770 6030
rect 28366 5842 28418 5854
rect 29038 5906 29090 5918
rect 29038 5842 29090 5854
rect 29710 5906 29762 5918
rect 30202 5910 30214 5962
rect 30266 5910 30278 5962
rect 30718 5954 30770 5966
rect 31632 6018 31684 6030
rect 30874 5910 30886 5962
rect 30938 5910 30950 5962
rect 31632 5954 31684 5966
rect 33164 6018 33216 6030
rect 38110 6018 38162 6030
rect 35130 5966 35142 6018
rect 35194 5966 35206 6018
rect 33164 5954 33216 5966
rect 29710 5842 29762 5854
rect 31390 5906 31442 5918
rect 31390 5842 31442 5854
rect 31950 5906 32002 5918
rect 31950 5842 32002 5854
rect 32174 5906 32226 5918
rect 32174 5842 32226 5854
rect 33406 5906 33458 5918
rect 33898 5910 33910 5962
rect 33962 5910 33974 5962
rect 38110 5954 38162 5966
rect 33406 5842 33458 5854
rect 34078 5906 34130 5918
rect 34078 5842 34130 5854
rect 34638 5906 34690 5918
rect 34638 5842 34690 5854
rect 34862 5906 34914 5918
rect 34862 5842 34914 5854
rect 35422 5906 35474 5918
rect 36194 5854 36206 5906
rect 36258 5854 36270 5906
rect 35422 5842 35474 5854
rect 20962 5742 20974 5794
rect 21026 5791 21038 5794
rect 21186 5791 21198 5794
rect 21026 5745 21198 5791
rect 21026 5742 21038 5745
rect 21186 5742 21198 5745
rect 21250 5742 21262 5794
rect 15150 5682 15202 5694
rect 15150 5618 15202 5630
rect 18510 5682 18562 5694
rect 22336 5682 22388 5694
rect 26238 5682 26290 5694
rect 20682 5630 20694 5682
rect 20746 5630 20758 5682
rect 23146 5630 23158 5682
rect 23210 5630 23222 5682
rect 32442 5630 32454 5682
rect 32506 5630 32518 5682
rect 18510 5618 18562 5630
rect 22336 5618 22388 5630
rect 26238 5618 26290 5630
rect 1344 5514 38640 5548
rect 1344 5462 5876 5514
rect 5928 5462 5980 5514
rect 6032 5462 6084 5514
rect 6136 5462 15200 5514
rect 15252 5462 15304 5514
rect 15356 5462 15408 5514
rect 15460 5462 24524 5514
rect 24576 5462 24628 5514
rect 24680 5462 24732 5514
rect 24784 5462 33848 5514
rect 33900 5462 33952 5514
rect 34004 5462 34056 5514
rect 34108 5462 38640 5514
rect 1344 5428 38640 5462
rect 37998 5346 38050 5358
rect 37998 5282 38050 5294
rect 14254 5234 14306 5246
rect 36262 5234 36314 5246
rect 8306 5182 8318 5234
rect 8370 5182 8382 5234
rect 10210 5182 10222 5234
rect 10274 5182 10286 5234
rect 16258 5182 16270 5234
rect 16322 5182 16334 5234
rect 18162 5182 18174 5234
rect 18226 5182 18238 5234
rect 25554 5182 25566 5234
rect 25618 5182 25630 5234
rect 27458 5182 27470 5234
rect 27522 5182 27534 5234
rect 32610 5182 32622 5234
rect 32674 5182 32686 5234
rect 35634 5182 35646 5234
rect 35698 5182 35710 5234
rect 14254 5170 14306 5182
rect 36262 5170 36314 5182
rect 37158 5234 37210 5246
rect 37158 5170 37210 5182
rect 6638 5122 6690 5134
rect 1922 5070 1934 5122
rect 1986 5070 1998 5122
rect 4162 5042 4174 5094
rect 4226 5042 4238 5094
rect 6638 5058 6690 5070
rect 7310 5122 7362 5134
rect 7310 5058 7362 5070
rect 7982 5122 8034 5134
rect 7982 5058 8034 5070
rect 11006 5122 11058 5134
rect 11006 5058 11058 5070
rect 13022 5122 13074 5134
rect 13022 5058 13074 5070
rect 15374 5122 15426 5134
rect 15374 5058 15426 5070
rect 15486 5122 15538 5134
rect 15486 5058 15538 5070
rect 20862 5122 20914 5134
rect 20862 5058 20914 5070
rect 23662 5122 23714 5134
rect 23662 5058 23714 5070
rect 24782 5122 24834 5134
rect 24782 5058 24834 5070
rect 29934 5122 29986 5134
rect 32958 5122 33010 5134
rect 38334 5122 38386 5134
rect 30706 5070 30718 5122
rect 30770 5070 30782 5122
rect 33730 5070 33742 5122
rect 33794 5070 33806 5122
rect 29934 5058 29986 5070
rect 32958 5058 33010 5070
rect 38334 5058 38386 5070
rect 6302 4898 6354 4910
rect 6302 4834 6354 4846
rect 6974 4898 7026 4910
rect 6974 4834 7026 4846
rect 7646 4898 7698 4910
rect 7646 4834 7698 4846
rect 11902 4898 11954 4910
rect 11902 4834 11954 4846
rect 18790 4898 18842 4910
rect 18790 4834 18842 4846
rect 19406 4898 19458 4910
rect 19406 4834 19458 4846
rect 22542 4898 22594 4910
rect 22542 4834 22594 4846
rect 37606 4898 37658 4910
rect 37606 4834 37658 4846
rect 1344 4730 38800 4764
rect 1344 4678 10538 4730
rect 10590 4678 10642 4730
rect 10694 4678 10746 4730
rect 10798 4678 19862 4730
rect 19914 4678 19966 4730
rect 20018 4678 20070 4730
rect 20122 4678 29186 4730
rect 29238 4678 29290 4730
rect 29342 4678 29394 4730
rect 29446 4678 38510 4730
rect 38562 4678 38614 4730
rect 38666 4678 38718 4730
rect 38770 4678 38800 4730
rect 1344 4644 38800 4678
rect 2774 4562 2826 4574
rect 2774 4498 2826 4510
rect 30718 4562 30770 4574
rect 30718 4498 30770 4510
rect 34078 4562 34130 4574
rect 34078 4498 34130 4510
rect 38278 4562 38330 4574
rect 38278 4498 38330 4510
rect 15822 4450 15874 4462
rect 21758 4450 21810 4462
rect 29598 4450 29650 4462
rect 17434 4398 17446 4450
rect 17498 4398 17510 4450
rect 26506 4398 26518 4450
rect 26570 4398 26582 4450
rect 15822 4386 15874 4398
rect 21758 4386 21810 4398
rect 29598 4386 29650 4398
rect 35086 4450 35138 4462
rect 35086 4386 35138 4398
rect 36000 4450 36052 4462
rect 3502 4338 3554 4350
rect 5842 4313 5854 4365
rect 5906 4313 5918 4365
rect 6514 4313 6526 4365
rect 6578 4313 6590 4365
rect 10098 4313 10110 4365
rect 10162 4313 10174 4365
rect 12574 4338 12626 4350
rect 15262 4338 15314 4350
rect 3502 4274 3554 4286
rect 13346 4286 13358 4338
rect 13410 4286 13422 4338
rect 12574 4274 12626 4286
rect 15262 4274 15314 4286
rect 15990 4338 16042 4350
rect 15990 4274 16042 4286
rect 16494 4338 16546 4350
rect 16494 4274 16546 4286
rect 16736 4338 16788 4350
rect 16736 4274 16788 4286
rect 17726 4338 17778 4350
rect 17726 4274 17778 4286
rect 17950 4338 18002 4350
rect 17950 4274 18002 4286
rect 18342 4338 18394 4350
rect 18342 4274 18394 4286
rect 18510 4338 18562 4350
rect 24446 4338 24498 4350
rect 19282 4286 19294 4338
rect 19346 4286 19358 4338
rect 23650 4286 23662 4338
rect 23714 4286 23726 4338
rect 18510 4274 18562 4286
rect 24446 4274 24498 4286
rect 26014 4338 26066 4350
rect 26014 4274 26066 4286
rect 26238 4338 26290 4350
rect 26238 4274 26290 4286
rect 26910 4338 26962 4350
rect 31838 4338 31890 4350
rect 27682 4286 27694 4338
rect 27746 4286 27758 4338
rect 26910 4274 26962 4286
rect 31838 4274 31890 4286
rect 32958 4338 33010 4350
rect 35242 4342 35254 4394
rect 35306 4342 35318 4394
rect 36000 4386 36052 4398
rect 32958 4274 33010 4286
rect 35758 4338 35810 4350
rect 35758 4274 35810 4286
rect 37830 4226 37882 4238
rect 21186 4174 21198 4226
rect 21250 4174 21262 4226
rect 37830 4162 37882 4174
rect 3166 4114 3218 4126
rect 3166 4050 3218 4062
rect 4846 4114 4898 4126
rect 4846 4050 4898 4062
rect 7534 4114 7586 4126
rect 7534 4050 7586 4062
rect 10894 4114 10946 4126
rect 10894 4050 10946 4062
rect 1344 3946 38640 3980
rect 1344 3894 5876 3946
rect 5928 3894 5980 3946
rect 6032 3894 6084 3946
rect 6136 3894 15200 3946
rect 15252 3894 15304 3946
rect 15356 3894 15408 3946
rect 15460 3894 24524 3946
rect 24576 3894 24628 3946
rect 24680 3894 24732 3946
rect 24784 3894 33848 3946
rect 33900 3894 33952 3946
rect 34004 3894 34056 3946
rect 34108 3894 38640 3946
rect 1344 3860 38640 3894
rect 5742 3778 5794 3790
rect 5742 3714 5794 3726
rect 9550 3778 9602 3790
rect 27470 3778 27522 3790
rect 13178 3726 13190 3778
rect 13242 3726 13254 3778
rect 9550 3714 9602 3726
rect 27470 3714 27522 3726
rect 28478 3778 28530 3790
rect 28478 3714 28530 3726
rect 30158 3778 30210 3790
rect 30158 3714 30210 3726
rect 32398 3778 32450 3790
rect 32398 3714 32450 3726
rect 33854 3778 33906 3790
rect 33854 3714 33906 3726
rect 36206 3778 36258 3790
rect 36206 3714 36258 3726
rect 37438 3778 37490 3790
rect 37438 3714 37490 3726
rect 3490 3614 3502 3666
rect 3554 3614 3566 3666
rect 22082 3614 22094 3666
rect 22146 3614 22158 3666
rect 25554 3614 25566 3666
rect 25618 3614 25630 3666
rect 6078 3554 6130 3566
rect 2818 3474 2830 3526
rect 2882 3474 2894 3526
rect 8318 3554 8370 3566
rect 6078 3490 6130 3502
rect 6626 3474 6638 3526
rect 6690 3474 6702 3526
rect 8318 3490 8370 3502
rect 9886 3554 9938 3566
rect 13470 3554 13522 3566
rect 9886 3490 9938 3502
rect 10210 3474 10222 3526
rect 10274 3474 10286 3526
rect 13470 3490 13522 3502
rect 13582 3554 13634 3566
rect 27806 3554 27858 3566
rect 13582 3490 13634 3502
rect 13906 3474 13918 3526
rect 13970 3474 13982 3526
rect 18050 3474 18062 3526
rect 18114 3474 18126 3526
rect 21074 3474 21086 3526
rect 21138 3474 21150 3526
rect 24546 3474 24558 3526
rect 24610 3474 24622 3526
rect 27806 3490 27858 3502
rect 28814 3554 28866 3566
rect 28814 3490 28866 3502
rect 29654 3554 29706 3566
rect 29654 3490 29706 3502
rect 30494 3554 30546 3566
rect 30494 3490 30546 3502
rect 30886 3554 30938 3566
rect 30886 3490 30938 3502
rect 31670 3554 31722 3566
rect 31670 3490 31722 3502
rect 32062 3554 32114 3566
rect 32062 3490 32114 3502
rect 33518 3554 33570 3566
rect 33518 3490 33570 3502
rect 35870 3554 35922 3566
rect 35870 3490 35922 3502
rect 37102 3554 37154 3566
rect 37102 3490 37154 3502
rect 37998 3554 38050 3566
rect 37998 3490 38050 3502
rect 38334 3554 38386 3566
rect 38334 3490 38386 3502
rect 29206 3442 29258 3454
rect 29206 3378 29258 3390
rect 33350 3442 33402 3454
rect 33350 3378 33402 3390
rect 35478 3442 35530 3454
rect 35478 3378 35530 3390
rect 36934 3442 36986 3454
rect 36934 3378 36986 3390
rect 11790 3330 11842 3342
rect 11790 3266 11842 3278
rect 15598 3330 15650 3342
rect 15598 3266 15650 3278
rect 19070 3330 19122 3342
rect 19070 3266 19122 3278
rect 1344 3162 38800 3196
rect 1344 3110 10538 3162
rect 10590 3110 10642 3162
rect 10694 3110 10746 3162
rect 10798 3110 19862 3162
rect 19914 3110 19966 3162
rect 20018 3110 20070 3162
rect 20122 3110 29186 3162
rect 29238 3110 29290 3162
rect 29342 3110 29394 3162
rect 29446 3110 38510 3162
rect 38562 3110 38614 3162
rect 38666 3110 38718 3162
rect 38770 3110 38800 3162
rect 1344 3076 38800 3110
<< via1 >>
rect 5876 36822 5928 36874
rect 5980 36822 6032 36874
rect 6084 36822 6136 36874
rect 15200 36822 15252 36874
rect 15304 36822 15356 36874
rect 15408 36822 15460 36874
rect 24524 36822 24576 36874
rect 24628 36822 24680 36874
rect 24732 36822 24784 36874
rect 33848 36822 33900 36874
rect 33952 36822 34004 36874
rect 34056 36822 34108 36874
rect 19182 36654 19234 36706
rect 33182 36542 33234 36594
rect 37606 36542 37658 36594
rect 10222 36402 10274 36454
rect 12350 36430 12402 36482
rect 13694 36430 13746 36482
rect 13918 36402 13970 36454
rect 16158 36430 16210 36482
rect 17390 36430 17442 36482
rect 19854 36402 19906 36454
rect 22766 36430 22818 36482
rect 23550 36430 23602 36482
rect 24558 36402 24610 36454
rect 27246 36430 27298 36482
rect 28590 36430 28642 36482
rect 30718 36402 30770 36454
rect 31054 36430 31106 36482
rect 32510 36402 32562 36454
rect 35422 36430 35474 36482
rect 38334 36430 38386 36482
rect 3446 36262 3498 36314
rect 4566 36262 4618 36314
rect 5686 36262 5738 36314
rect 6806 36262 6858 36314
rect 7926 36262 7978 36314
rect 8710 36262 8762 36314
rect 9718 36262 9770 36314
rect 20862 36318 20914 36370
rect 36150 36318 36202 36370
rect 13358 36206 13410 36258
rect 17054 36206 17106 36258
rect 23942 36206 23994 36258
rect 25902 36206 25954 36258
rect 27582 36206 27634 36258
rect 31390 36206 31442 36258
rect 35086 36206 35138 36258
rect 37998 36206 38050 36258
rect 10538 36038 10590 36090
rect 10642 36038 10694 36090
rect 10746 36038 10798 36090
rect 19862 36038 19914 36090
rect 19966 36038 20018 36090
rect 20070 36038 20122 36090
rect 29186 36038 29238 36090
rect 29290 36038 29342 36090
rect 29394 36038 29446 36090
rect 38510 36038 38562 36090
rect 38614 36038 38666 36090
rect 38718 36038 38770 36090
rect 11286 35870 11338 35922
rect 30942 35870 30994 35922
rect 8878 35758 8930 35810
rect 20974 35758 21026 35810
rect 2494 35646 2546 35698
rect 5798 35646 5850 35698
rect 6190 35646 6242 35698
rect 12238 35646 12290 35698
rect 12350 35646 12402 35698
rect 15710 35646 15762 35698
rect 16046 35646 16098 35698
rect 16270 35685 16322 35737
rect 16606 35646 16658 35698
rect 17278 35646 17330 35698
rect 23662 35646 23714 35698
rect 24782 35646 24834 35698
rect 25230 35673 25282 35725
rect 28030 35673 28082 35725
rect 31278 35646 31330 35698
rect 31726 35646 31778 35698
rect 33070 35673 33122 35725
rect 35758 35646 35810 35698
rect 36430 35646 36482 35698
rect 3278 35534 3330 35586
rect 5182 35534 5234 35586
rect 6974 35534 7026 35586
rect 9718 35534 9770 35586
rect 10950 35534 11002 35586
rect 13134 35534 13186 35586
rect 15038 35534 15090 35586
rect 16494 35534 16546 35586
rect 18062 35534 18114 35586
rect 19966 35534 20018 35586
rect 20582 35534 20634 35586
rect 22878 35534 22930 35586
rect 24054 35534 24106 35586
rect 11902 35422 11954 35474
rect 24446 35422 24498 35474
rect 26238 35422 26290 35474
rect 29038 35422 29090 35474
rect 32062 35422 32114 35474
rect 34414 35422 34466 35474
rect 36094 35422 36146 35474
rect 36766 35422 36818 35474
rect 5876 35254 5928 35306
rect 5980 35254 6032 35306
rect 6084 35254 6136 35306
rect 15200 35254 15252 35306
rect 15304 35254 15356 35306
rect 15408 35254 15460 35306
rect 24524 35254 24576 35306
rect 24628 35254 24680 35306
rect 24732 35254 24784 35306
rect 33848 35254 33900 35306
rect 33952 35254 34004 35306
rect 34056 35254 34108 35306
rect 2942 35086 2994 35138
rect 8766 35086 8818 35138
rect 15374 35086 15426 35138
rect 22318 35086 22370 35138
rect 24334 35086 24386 35138
rect 9494 34974 9546 35026
rect 9942 34974 9994 35026
rect 12798 34974 12850 35026
rect 16718 34974 16770 35026
rect 19966 34974 20018 35026
rect 20806 34974 20858 35026
rect 25790 34974 25842 35026
rect 4062 34862 4114 34914
rect 5518 34862 5570 34914
rect 6302 34862 6354 34914
rect 9102 34862 9154 34914
rect 10110 34862 10162 34914
rect 10894 34862 10946 34914
rect 13750 34862 13802 34914
rect 13918 34862 13970 34914
rect 15934 34862 15986 34914
rect 19630 34862 19682 34914
rect 20302 34862 20354 34914
rect 8206 34750 8258 34802
rect 19966 34806 20018 34858
rect 21534 34834 21586 34886
rect 23998 34862 24050 34914
rect 25006 34862 25058 34914
rect 28030 34862 28082 34914
rect 28254 34862 28306 34914
rect 28534 34862 28586 34914
rect 29038 34862 29090 34914
rect 30494 34862 30546 34914
rect 31054 34862 31106 34914
rect 31838 34862 31890 34914
rect 34638 34862 34690 34914
rect 35310 34862 35362 34914
rect 35422 34862 35474 34914
rect 18622 34750 18674 34802
rect 27694 34750 27746 34802
rect 33742 34750 33794 34802
rect 36374 34750 36426 34802
rect 34302 34638 34354 34690
rect 34974 34638 35026 34690
rect 35758 34638 35810 34690
rect 37830 34638 37882 34690
rect 38278 34638 38330 34690
rect 10538 34470 10590 34522
rect 10642 34470 10694 34522
rect 10746 34470 10798 34522
rect 19862 34470 19914 34522
rect 19966 34470 20018 34522
rect 20070 34470 20122 34522
rect 29186 34470 29238 34522
rect 29290 34470 29342 34522
rect 29394 34470 29446 34522
rect 38510 34470 38562 34522
rect 38614 34470 38666 34522
rect 38718 34470 38770 34522
rect 5966 34302 6018 34354
rect 10894 34302 10946 34354
rect 15710 34302 15762 34354
rect 17950 34246 18002 34298
rect 18790 34302 18842 34354
rect 20414 34302 20466 34354
rect 28926 34190 28978 34242
rect 7086 34078 7138 34130
rect 8598 34078 8650 34130
rect 8878 34078 8930 34130
rect 8990 34078 9042 34130
rect 9438 34078 9490 34130
rect 11790 34105 11842 34157
rect 14366 34105 14418 34157
rect 17614 34078 17666 34130
rect 17838 34117 17890 34169
rect 18174 34078 18226 34130
rect 19070 34105 19122 34157
rect 21870 34078 21922 34130
rect 27470 34078 27522 34130
rect 28254 34078 28306 34130
rect 31614 34078 31666 34130
rect 31726 34078 31778 34130
rect 32958 34078 33010 34130
rect 33742 34078 33794 34130
rect 36262 34078 36314 34130
rect 37662 34078 37714 34130
rect 38334 34078 38386 34130
rect 12574 33966 12626 34018
rect 22654 33966 22706 34018
rect 24558 33966 24610 34018
rect 25566 33966 25618 34018
rect 30830 33966 30882 34018
rect 32062 33966 32114 34018
rect 35646 33966 35698 34018
rect 36710 33966 36762 34018
rect 37326 33966 37378 34018
rect 7422 33854 7474 33906
rect 7758 33854 7810 33906
rect 37998 33854 38050 33906
rect 5876 33686 5928 33738
rect 5980 33686 6032 33738
rect 6084 33686 6136 33738
rect 15200 33686 15252 33738
rect 15304 33686 15356 33738
rect 15408 33686 15460 33738
rect 24524 33686 24576 33738
rect 24628 33686 24680 33738
rect 24732 33686 24784 33738
rect 33848 33686 33900 33738
rect 33952 33686 34004 33738
rect 34056 33686 34108 33738
rect 9046 33518 9098 33570
rect 14758 33518 14810 33570
rect 16158 33518 16210 33570
rect 18958 33518 19010 33570
rect 22654 33518 22706 33570
rect 25678 33518 25730 33570
rect 10446 33406 10498 33458
rect 12350 33406 12402 33458
rect 30588 33406 30640 33458
rect 32510 33406 32562 33458
rect 8766 33294 8818 33346
rect 9326 33294 9378 33346
rect 9438 33294 9490 33346
rect 10054 33294 10106 33346
rect 10782 33294 10834 33346
rect 11454 33294 11506 33346
rect 11902 33294 11954 33346
rect 12462 33294 12514 33346
rect 13806 33294 13858 33346
rect 12238 33238 12290 33290
rect 13918 33294 13970 33346
rect 14254 33294 14306 33346
rect 14478 33294 14530 33346
rect 15486 33266 15538 33318
rect 17950 33266 18002 33318
rect 21310 33238 21362 33290
rect 13526 33182 13578 33234
rect 21422 33238 21474 33290
rect 22150 33294 22202 33346
rect 22318 33294 22370 33346
rect 22990 33294 23042 33346
rect 25006 33294 25058 33346
rect 25118 33294 25170 33346
rect 25284 33294 25336 33346
rect 26462 33266 26514 33318
rect 27806 33294 27858 33346
rect 29822 33294 29874 33346
rect 21982 33182 22034 33234
rect 24278 33182 24330 33234
rect 29318 33238 29370 33290
rect 30830 33294 30882 33346
rect 31334 33350 31386 33402
rect 31726 33294 31778 33346
rect 35534 33350 35586 33402
rect 37662 33294 37714 33346
rect 29150 33182 29202 33234
rect 30064 33182 30116 33234
rect 31502 33182 31554 33234
rect 34414 33182 34466 33234
rect 35030 33238 35082 33290
rect 34862 33182 34914 33234
rect 35776 33182 35828 33234
rect 37158 33238 37210 33290
rect 36990 33182 37042 33234
rect 37904 33182 37956 33234
rect 8430 33070 8482 33122
rect 11118 33070 11170 33122
rect 23326 33070 23378 33122
rect 24726 33070 24778 33122
rect 36374 33070 36426 33122
rect 10538 32902 10590 32954
rect 10642 32902 10694 32954
rect 10746 32902 10798 32954
rect 19862 32902 19914 32954
rect 19966 32902 20018 32954
rect 20070 32902 20122 32954
rect 29186 32902 29238 32954
rect 29290 32902 29342 32954
rect 29394 32902 29446 32954
rect 38510 32902 38562 32954
rect 38614 32902 38666 32954
rect 38718 32902 38770 32954
rect 5686 32734 5738 32786
rect 13022 32734 13074 32786
rect 24278 32734 24330 32786
rect 9606 32622 9658 32674
rect 18846 32678 18898 32730
rect 17502 32622 17554 32674
rect 2382 32510 2434 32562
rect 7198 32510 7250 32562
rect 7758 32510 7810 32562
rect 8094 32525 8146 32577
rect 8430 32510 8482 32562
rect 9886 32566 9938 32618
rect 19630 32622 19682 32674
rect 8654 32510 8706 32562
rect 10110 32538 10162 32590
rect 10334 32538 10386 32590
rect 10502 32526 10554 32578
rect 10894 32510 10946 32562
rect 11118 32510 11170 32562
rect 11678 32510 11730 32562
rect 11902 32525 11954 32577
rect 14142 32510 14194 32562
rect 14366 32510 14418 32562
rect 14702 32510 14754 32562
rect 15710 32510 15762 32562
rect 15934 32525 15986 32577
rect 16494 32525 16546 32577
rect 16718 32510 16770 32562
rect 17838 32510 17890 32562
rect 18062 32510 18114 32562
rect 18398 32537 18450 32589
rect 18734 32510 18786 32562
rect 19462 32566 19514 32618
rect 22990 32622 23042 32674
rect 24614 32678 24666 32730
rect 29710 32734 29762 32786
rect 19294 32510 19346 32562
rect 19742 32510 19794 32562
rect 20022 32510 20074 32562
rect 20414 32510 20466 32562
rect 20526 32510 20578 32562
rect 20672 32548 20724 32600
rect 21422 32510 21474 32562
rect 22598 32566 22650 32618
rect 23158 32566 23210 32618
rect 31446 32622 31498 32674
rect 21646 32510 21698 32562
rect 22766 32510 22818 32562
rect 23662 32510 23714 32562
rect 24782 32510 24834 32562
rect 25678 32538 25730 32590
rect 26294 32566 26346 32618
rect 25902 32510 25954 32562
rect 26574 32510 26626 32562
rect 26686 32510 26738 32562
rect 26844 32560 26896 32612
rect 28030 32537 28082 32589
rect 30942 32510 30994 32562
rect 31166 32510 31218 32562
rect 31950 32510 32002 32562
rect 32174 32510 32226 32562
rect 35198 32510 35250 32562
rect 35310 32510 35362 32562
rect 3166 32398 3218 32450
rect 5070 32398 5122 32450
rect 8206 32398 8258 32450
rect 7366 32342 7418 32394
rect 12014 32398 12066 32450
rect 15318 32398 15370 32450
rect 16046 32398 16098 32450
rect 16382 32398 16434 32450
rect 21086 32398 21138 32450
rect 11230 32342 11282 32394
rect 14702 32342 14754 32394
rect 26126 32398 26178 32450
rect 27246 32398 27298 32450
rect 34078 32398 34130 32450
rect 36094 32398 36146 32450
rect 37998 32398 38050 32450
rect 8934 32286 8986 32338
rect 21926 32286 21978 32338
rect 23494 32286 23546 32338
rect 32454 32286 32506 32338
rect 5876 32118 5928 32170
rect 5980 32118 6032 32170
rect 6084 32118 6136 32170
rect 15200 32118 15252 32170
rect 15304 32118 15356 32170
rect 15408 32118 15460 32170
rect 24524 32118 24576 32170
rect 24628 32118 24680 32170
rect 24732 32118 24784 32170
rect 33848 32118 33900 32170
rect 33952 32118 34004 32170
rect 34056 32118 34108 32170
rect 3166 31950 3218 32002
rect 11118 31950 11170 32002
rect 14310 31950 14362 32002
rect 22766 31950 22818 32002
rect 25230 31950 25282 32002
rect 4286 31726 4338 31778
rect 4398 31726 4450 31778
rect 4622 31726 4674 31778
rect 7758 31726 7810 31778
rect 7254 31670 7306 31722
rect 8000 31726 8052 31778
rect 8598 31782 8650 31834
rect 9344 31838 9396 31890
rect 9830 31838 9882 31890
rect 16718 31838 16770 31890
rect 19966 31838 20018 31890
rect 24222 31838 24274 31890
rect 29150 31838 29202 31890
rect 31502 31838 31554 31890
rect 34190 31838 34242 31890
rect 35926 31838 35978 31890
rect 9102 31726 9154 31778
rect 10110 31698 10162 31750
rect 4902 31614 4954 31666
rect 7086 31614 7138 31666
rect 10334 31670 10386 31722
rect 10558 31698 10610 31750
rect 10726 31710 10778 31762
rect 11678 31726 11730 31778
rect 11790 31726 11842 31778
rect 11510 31670 11562 31722
rect 12126 31726 12178 31778
rect 12686 31726 12738 31778
rect 13470 31670 13522 31722
rect 13582 31670 13634 31722
rect 13806 31670 13858 31722
rect 14030 31698 14082 31750
rect 14590 31726 14642 31778
rect 14814 31726 14866 31778
rect 15822 31726 15874 31778
rect 15934 31726 15986 31778
rect 16270 31726 16322 31778
rect 16606 31682 16658 31734
rect 17278 31726 17330 31778
rect 18062 31726 18114 31778
rect 20302 31726 20354 31778
rect 22094 31726 22146 31778
rect 22206 31726 22258 31778
rect 22374 31726 22426 31778
rect 23438 31726 23490 31778
rect 23774 31726 23826 31778
rect 24334 31726 24386 31778
rect 25566 31726 25618 31778
rect 24110 31670 24162 31722
rect 26014 31698 26066 31750
rect 29262 31711 29314 31763
rect 29486 31726 29538 31778
rect 32286 31698 32338 31750
rect 32846 31698 32898 31750
rect 36206 31726 36258 31778
rect 36318 31726 36370 31778
rect 37158 31726 37210 31778
rect 37662 31726 37714 31778
rect 8430 31614 8482 31666
rect 15094 31614 15146 31666
rect 15542 31614 15594 31666
rect 36990 31614 37042 31666
rect 12574 31558 12626 31610
rect 37904 31614 37956 31666
rect 20638 31502 20690 31554
rect 10538 31334 10590 31386
rect 10642 31334 10694 31386
rect 10746 31334 10798 31386
rect 19862 31334 19914 31386
rect 19966 31334 20018 31386
rect 20070 31334 20122 31386
rect 29186 31334 29238 31386
rect 29290 31334 29342 31386
rect 29394 31334 29446 31386
rect 38510 31334 38562 31386
rect 38614 31334 38666 31386
rect 38718 31334 38770 31386
rect 7422 31110 7474 31162
rect 5742 31054 5794 31106
rect 6582 31054 6634 31106
rect 8038 31054 8090 31106
rect 11660 31054 11712 31106
rect 1990 30998 2042 31050
rect 15206 31054 15258 31106
rect 1822 30942 1874 30994
rect 2494 30942 2546 30994
rect 3054 30942 3106 30994
rect 6078 30942 6130 30994
rect 6302 30942 6354 30994
rect 7310 30957 7362 31009
rect 7646 30942 7698 30994
rect 8318 30942 8370 30994
rect 8542 30942 8594 30994
rect 12406 30998 12458 31050
rect 10054 30942 10106 30994
rect 10222 30942 10274 30994
rect 2736 30830 2788 30882
rect 3838 30830 3890 30882
rect 9662 30830 9714 30882
rect 10334 30886 10386 30938
rect 11902 30942 11954 30994
rect 12574 30942 12626 30994
rect 13246 30942 13298 30994
rect 13358 30942 13410 30994
rect 13526 30942 13578 30994
rect 14366 30998 14418 31050
rect 14478 30998 14530 31050
rect 14702 30970 14754 31022
rect 14926 30970 14978 31022
rect 15710 30998 15762 31050
rect 16270 31054 16322 31106
rect 21702 31054 21754 31106
rect 33164 31054 33216 31106
rect 16046 30942 16098 30994
rect 16942 30942 16994 30994
rect 17502 30942 17554 30994
rect 17838 30942 17890 30994
rect 19518 30942 19570 30994
rect 13918 30830 13970 30882
rect 16438 30886 16490 30938
rect 19854 30942 19906 30994
rect 19966 30942 20018 30994
rect 20190 30942 20242 30994
rect 21198 30942 21250 30994
rect 21422 30942 21474 30994
rect 22318 30942 22370 30994
rect 22654 30942 22706 30994
rect 22878 30981 22930 31033
rect 23326 30942 23378 30994
rect 23774 30942 23826 30994
rect 24110 30942 24162 30994
rect 25454 30942 25506 30994
rect 25678 30942 25730 30994
rect 26014 30942 26066 30994
rect 26798 30942 26850 30994
rect 29038 30942 29090 30994
rect 29262 30942 29314 30994
rect 30382 30969 30434 31021
rect 33406 30942 33458 30994
rect 21030 30830 21082 30882
rect 17726 30774 17778 30826
rect 22990 30830 23042 30882
rect 33910 30886 33962 30938
rect 34078 30942 34130 30994
rect 34302 30942 34354 30994
rect 36990 30942 37042 30994
rect 37326 30942 37378 30994
rect 24726 30830 24778 30882
rect 28702 30830 28754 30882
rect 29542 30830 29594 30882
rect 35086 30830 35138 30882
rect 37662 30830 37714 30882
rect 25790 30774 25842 30826
rect 16774 30718 16826 30770
rect 20470 30718 20522 30770
rect 5876 30550 5928 30602
rect 5980 30550 6032 30602
rect 6084 30550 6136 30602
rect 15200 30550 15252 30602
rect 15304 30550 15356 30602
rect 15408 30550 15460 30602
rect 24524 30550 24576 30602
rect 24628 30550 24680 30602
rect 24732 30550 24784 30602
rect 33848 30550 33900 30602
rect 33952 30550 34004 30602
rect 34056 30550 34108 30602
rect 3726 30382 3778 30434
rect 8262 30382 8314 30434
rect 12798 30382 12850 30434
rect 9550 30270 9602 30322
rect 13526 30326 13578 30378
rect 17950 30382 18002 30434
rect 22150 30382 22202 30434
rect 31726 30382 31778 30434
rect 1878 30158 1930 30210
rect 2382 30158 2434 30210
rect 2624 30158 2676 30210
rect 4846 30158 4898 30210
rect 6134 30158 6186 30210
rect 6862 30158 6914 30210
rect 7534 30158 7586 30210
rect 7030 30102 7082 30154
rect 7776 30158 7828 30210
rect 8542 30102 8594 30154
rect 8766 30102 8818 30154
rect 8990 30130 9042 30182
rect 10110 30158 10162 30210
rect 10222 30158 10274 30210
rect 9102 30102 9154 30154
rect 9944 30102 9996 30154
rect 14198 30214 14250 30266
rect 14944 30270 14996 30322
rect 17110 30270 17162 30322
rect 36038 30270 36090 30322
rect 10446 30158 10498 30210
rect 12238 30158 12290 30210
rect 13694 30158 13746 30210
rect 14702 30158 14754 30210
rect 12126 30102 12178 30154
rect 12406 30102 12458 30154
rect 15542 30158 15594 30210
rect 16046 30158 16098 30210
rect 16288 30158 16340 30210
rect 17614 30158 17666 30210
rect 19630 30158 19682 30210
rect 20190 30158 20242 30210
rect 20302 30158 20354 30210
rect 21310 30158 21362 30210
rect 21422 30158 21474 30210
rect 21702 30158 21754 30210
rect 22430 30158 22482 30210
rect 22542 30158 22594 30210
rect 22878 30158 22930 30210
rect 1710 30046 1762 30098
rect 14030 30046 14082 30098
rect 22710 30102 22762 30154
rect 23774 30158 23826 30210
rect 24558 30158 24610 30210
rect 26462 30158 26514 30210
rect 27078 30158 27130 30210
rect 27694 30158 27746 30210
rect 28030 30158 28082 30210
rect 28142 30158 28194 30210
rect 29486 30158 29538 30210
rect 29598 30158 29650 30210
rect 29878 30158 29930 30210
rect 32398 30130 32450 30182
rect 35310 30130 35362 30182
rect 37158 30158 37210 30210
rect 37662 30158 37714 30210
rect 15374 30046 15426 30098
rect 19910 30046 19962 30098
rect 36990 30046 37042 30098
rect 37904 30046 37956 30098
rect 10782 29934 10834 29986
rect 11398 29934 11450 29986
rect 11846 29934 11898 29986
rect 19294 29934 19346 29986
rect 28478 29934 28530 29986
rect 34190 29934 34242 29986
rect 10538 29766 10590 29818
rect 10642 29766 10694 29818
rect 10746 29766 10798 29818
rect 19862 29766 19914 29818
rect 19966 29766 20018 29818
rect 20070 29766 20122 29818
rect 29186 29766 29238 29818
rect 29290 29766 29342 29818
rect 29394 29766 29446 29818
rect 38510 29766 38562 29818
rect 38614 29766 38666 29818
rect 38718 29766 38770 29818
rect 11230 29598 11282 29650
rect 12126 29598 12178 29650
rect 14534 29598 14586 29650
rect 23774 29598 23826 29650
rect 14926 29542 14978 29594
rect 29094 29598 29146 29650
rect 33238 29598 33290 29650
rect 8150 29486 8202 29538
rect 13936 29486 13988 29538
rect 2494 29374 2546 29426
rect 5462 29430 5514 29482
rect 4958 29374 5010 29426
rect 5630 29374 5682 29426
rect 7310 29389 7362 29441
rect 7646 29374 7698 29426
rect 8430 29374 8482 29426
rect 8654 29374 8706 29426
rect 9550 29374 9602 29426
rect 9886 29374 9938 29426
rect 10782 29374 10834 29426
rect 10894 29374 10946 29426
rect 12462 29374 12514 29426
rect 13190 29430 13242 29482
rect 19910 29486 19962 29538
rect 13022 29374 13074 29426
rect 13694 29374 13746 29426
rect 15262 29430 15314 29482
rect 19350 29430 19402 29482
rect 25510 29486 25562 29538
rect 15038 29374 15090 29426
rect 15598 29374 15650 29426
rect 19182 29374 19234 29426
rect 19518 29374 19570 29426
rect 19630 29374 19682 29426
rect 20750 29430 20802 29482
rect 20526 29374 20578 29426
rect 21198 29374 21250 29426
rect 21646 29374 21698 29426
rect 22318 29374 22370 29426
rect 22878 29374 22930 29426
rect 23438 29374 23490 29426
rect 26126 29401 26178 29453
rect 29262 29430 29314 29482
rect 32062 29486 32114 29538
rect 29374 29374 29426 29426
rect 33854 29374 33906 29426
rect 36094 29401 36146 29453
rect 38222 29374 38274 29426
rect 7198 29262 7250 29314
rect 17558 29262 17610 29314
rect 3614 29150 3666 29202
rect 9662 29206 9714 29258
rect 18230 29262 18282 29314
rect 18678 29262 18730 29314
rect 20862 29262 20914 29314
rect 4716 29150 4768 29202
rect 21534 29206 21586 29258
rect 22710 29206 22762 29258
rect 24726 29262 24778 29314
rect 28758 29262 28810 29314
rect 30158 29262 30210 29314
rect 10446 29150 10498 29202
rect 26798 29150 26850 29202
rect 36766 29150 36818 29202
rect 5876 28982 5928 29034
rect 5980 28982 6032 29034
rect 6084 28982 6136 29034
rect 15200 28982 15252 29034
rect 15304 28982 15356 29034
rect 15408 28982 15460 29034
rect 24524 28982 24576 29034
rect 24628 28982 24680 29034
rect 24732 28982 24784 29034
rect 33848 28982 33900 29034
rect 33952 28982 34004 29034
rect 34056 28982 34108 29034
rect 7086 28814 7138 28866
rect 8374 28814 8426 28866
rect 11342 28814 11394 28866
rect 12126 28814 12178 28866
rect 16886 28814 16938 28866
rect 19872 28814 19924 28866
rect 22262 28814 22314 28866
rect 3054 28702 3106 28754
rect 4958 28702 5010 28754
rect 5798 28702 5850 28754
rect 6582 28702 6634 28754
rect 10222 28702 10274 28754
rect 12742 28702 12794 28754
rect 13638 28702 13690 28754
rect 20526 28758 20578 28810
rect 25454 28814 25506 28866
rect 30960 28814 31012 28866
rect 34750 28814 34802 28866
rect 2270 28590 2322 28642
rect 6750 28590 6802 28642
rect 7646 28575 7698 28627
rect 7982 28590 8034 28642
rect 8654 28562 8706 28614
rect 8878 28562 8930 28614
rect 9046 28534 9098 28586
rect 9214 28555 9266 28607
rect 10446 28590 10498 28642
rect 10054 28534 10106 28586
rect 10782 28534 10834 28586
rect 11678 28590 11730 28642
rect 11790 28590 11842 28642
rect 16158 28590 16210 28642
rect 16326 28646 16378 28698
rect 17390 28702 17442 28754
rect 19126 28646 19178 28698
rect 16606 28590 16658 28642
rect 17950 28590 18002 28642
rect 18062 28590 18114 28642
rect 18734 28590 18786 28642
rect 19630 28590 19682 28642
rect 20414 28590 20466 28642
rect 20638 28590 20690 28642
rect 21534 28590 21586 28642
rect 21702 28646 21754 28698
rect 22766 28702 22818 28754
rect 24502 28702 24554 28754
rect 28478 28702 28530 28754
rect 17784 28534 17836 28586
rect 21982 28590 22034 28642
rect 23102 28590 23154 28642
rect 24782 28590 24834 28642
rect 24894 28590 24946 28642
rect 25060 28590 25112 28642
rect 25790 28590 25842 28642
rect 26574 28590 26626 28642
rect 29262 28590 29314 28642
rect 29598 28590 29650 28642
rect 30214 28590 30266 28642
rect 30718 28590 30770 28642
rect 32062 28590 32114 28642
rect 7646 28422 7698 28474
rect 16494 28478 16546 28530
rect 18958 28478 19010 28530
rect 21870 28478 21922 28530
rect 31558 28534 31610 28586
rect 32846 28590 32898 28642
rect 33070 28590 33122 28642
rect 37158 28646 37210 28698
rect 36430 28562 36482 28614
rect 37662 28590 37714 28642
rect 31390 28478 31442 28530
rect 18566 28366 18618 28418
rect 30270 28422 30322 28474
rect 32304 28478 32356 28530
rect 33350 28478 33402 28530
rect 36990 28478 37042 28530
rect 37904 28478 37956 28530
rect 23494 28366 23546 28418
rect 10538 28198 10590 28250
rect 10642 28198 10694 28250
rect 10746 28198 10798 28250
rect 19862 28198 19914 28250
rect 19966 28198 20018 28250
rect 20070 28198 20122 28250
rect 29186 28198 29238 28250
rect 29290 28198 29342 28250
rect 29394 28198 29446 28250
rect 38510 28198 38562 28250
rect 38614 28198 38666 28250
rect 38718 28198 38770 28250
rect 9718 28030 9770 28082
rect 13022 28030 13074 28082
rect 14814 28030 14866 28082
rect 18286 28030 18338 28082
rect 22150 28030 22202 28082
rect 28142 28030 28194 28082
rect 2998 27918 3050 27970
rect 7646 27918 7698 27970
rect 8560 27918 8612 27970
rect 3278 27806 3330 27858
rect 3502 27806 3554 27858
rect 7814 27862 7866 27914
rect 10166 27918 10218 27970
rect 24670 27974 24722 28026
rect 29206 28030 29258 28082
rect 30046 28030 30098 28082
rect 10558 27918 10610 27970
rect 16438 27918 16490 27970
rect 27134 27918 27186 27970
rect 30998 27918 31050 27970
rect 37438 27918 37490 27970
rect 4398 27806 4450 27858
rect 8318 27806 8370 27858
rect 9830 27806 9882 27858
rect 10446 27806 10498 27858
rect 10726 27806 10778 27858
rect 10894 27806 10946 27858
rect 11230 27806 11282 27858
rect 11342 27806 11394 27858
rect 11510 27806 11562 27858
rect 14142 27806 14194 27858
rect 15150 27806 15202 27858
rect 16718 27806 16770 27858
rect 16830 27806 16882 27858
rect 17838 27806 17890 27858
rect 17950 27806 18002 27858
rect 18734 27806 18786 27858
rect 18846 27806 18898 27858
rect 19012 27806 19064 27858
rect 20078 27806 20130 27858
rect 20190 27806 20242 27858
rect 20336 27843 20388 27895
rect 25585 27862 25637 27914
rect 21198 27806 21250 27858
rect 21534 27806 21586 27858
rect 23886 27806 23938 27858
rect 24558 27806 24610 27858
rect 25342 27806 25394 27858
rect 26462 27806 26514 27858
rect 26966 27862 27018 27914
rect 26798 27806 26850 27858
rect 27246 27806 27298 27858
rect 27526 27806 27578 27858
rect 27806 27806 27858 27858
rect 28814 27806 28866 27858
rect 30382 27806 30434 27858
rect 30494 27806 30546 27858
rect 30718 27806 30770 27858
rect 31502 27806 31554 27858
rect 31670 27806 31722 27858
rect 32174 27806 32226 27858
rect 32416 27806 32468 27858
rect 33238 27862 33290 27914
rect 33070 27806 33122 27858
rect 33742 27806 33794 27858
rect 34750 27806 34802 27858
rect 38334 27806 38386 27858
rect 11902 27694 11954 27746
rect 19406 27694 19458 27746
rect 20750 27694 20802 27746
rect 5518 27582 5570 27634
rect 17502 27582 17554 27634
rect 21646 27638 21698 27690
rect 28646 27638 28698 27690
rect 29654 27694 29706 27746
rect 35534 27694 35586 27746
rect 33984 27582 34036 27634
rect 37998 27582 38050 27634
rect 5876 27414 5928 27466
rect 5980 27414 6032 27466
rect 6084 27414 6136 27466
rect 15200 27414 15252 27466
rect 15304 27414 15356 27466
rect 15408 27414 15460 27466
rect 24524 27414 24576 27466
rect 24628 27414 24680 27466
rect 24732 27414 24784 27466
rect 33848 27414 33900 27466
rect 33952 27414 34004 27466
rect 34056 27414 34108 27466
rect 8206 27246 8258 27298
rect 14012 27246 14064 27298
rect 17726 27246 17778 27298
rect 18566 27246 18618 27298
rect 4230 27134 4282 27186
rect 9886 27134 9938 27186
rect 11790 27134 11842 27186
rect 12854 27134 12906 27186
rect 13638 27134 13690 27186
rect 8598 27022 8650 27074
rect 8766 27022 8818 27074
rect 8878 27022 8930 27074
rect 9102 27022 9154 27074
rect 12126 27022 12178 27074
rect 14254 27022 14306 27074
rect 14758 27078 14810 27130
rect 19966 27134 20018 27186
rect 21310 27190 21362 27242
rect 24446 27246 24498 27298
rect 26966 27246 27018 27298
rect 30494 27246 30546 27298
rect 32678 27246 32730 27298
rect 34750 27246 34802 27298
rect 27862 27134 27914 27186
rect 29318 27134 29370 27186
rect 31614 27134 31666 27186
rect 15262 27022 15314 27074
rect 15430 27022 15482 27074
rect 15934 27022 15986 27074
rect 16176 27022 16228 27074
rect 17390 27022 17442 27074
rect 18846 27022 18898 27074
rect 19070 27022 19122 27074
rect 19294 27022 19346 27074
rect 19406 27022 19458 27074
rect 19572 27022 19624 27074
rect 20806 27022 20858 27074
rect 21422 27022 21474 27074
rect 21646 27022 21698 27074
rect 23774 27022 23826 27074
rect 23886 27022 23938 27074
rect 24052 27022 24104 27074
rect 25118 27022 25170 27074
rect 25678 27022 25730 27074
rect 26014 27022 26066 27074
rect 25342 26966 25394 27018
rect 26238 27022 26290 27074
rect 26518 27022 26570 27074
rect 27246 27022 27298 27074
rect 27358 27022 27410 27074
rect 30830 27022 30882 27074
rect 31278 27022 31330 27074
rect 31950 27022 32002 27074
rect 32286 27022 32338 27074
rect 31502 26966 31554 27018
rect 32398 27022 32450 27074
rect 33406 26994 33458 27046
rect 36486 27022 36538 27074
rect 37326 27022 37378 27074
rect 37830 27078 37882 27130
rect 14926 26910 14978 26962
rect 37084 26910 37136 26962
rect 25230 26854 25282 26906
rect 37998 26910 38050 26962
rect 28310 26798 28362 26850
rect 10538 26630 10590 26682
rect 10642 26630 10694 26682
rect 10746 26630 10798 26682
rect 19862 26630 19914 26682
rect 19966 26630 20018 26682
rect 20070 26630 20122 26682
rect 29186 26630 29238 26682
rect 29290 26630 29342 26682
rect 29394 26630 29446 26682
rect 38510 26630 38562 26682
rect 38614 26630 38666 26682
rect 38718 26630 38770 26682
rect 11286 26462 11338 26514
rect 13358 26462 13410 26514
rect 16718 26462 16770 26514
rect 26574 26462 26626 26514
rect 7198 26350 7250 26402
rect 3110 26294 3162 26346
rect 21198 26406 21250 26458
rect 27190 26462 27242 26514
rect 33238 26462 33290 26514
rect 35086 26462 35138 26514
rect 20320 26350 20372 26402
rect 2942 26238 2994 26290
rect 3614 26238 3666 26290
rect 4510 26238 4562 26290
rect 5294 26238 5346 26290
rect 10446 26238 10498 26290
rect 10670 26238 10722 26290
rect 12350 26265 12402 26317
rect 16382 26238 16434 26290
rect 17278 26238 17330 26290
rect 19574 26294 19626 26346
rect 25958 26350 26010 26402
rect 30326 26350 30378 26402
rect 19406 26238 19458 26290
rect 20078 26238 20130 26290
rect 21030 26267 21082 26319
rect 21310 26238 21362 26290
rect 24222 26238 24274 26290
rect 25230 26238 25282 26290
rect 25566 26238 25618 26290
rect 25678 26238 25730 26290
rect 7814 26126 7866 26178
rect 3856 26014 3908 26066
rect 10334 26070 10386 26122
rect 14982 26126 15034 26178
rect 24558 26126 24610 26178
rect 25398 26182 25450 26234
rect 26238 26238 26290 26290
rect 28198 26238 28250 26290
rect 30606 26238 30658 26290
rect 30718 26238 30770 26290
rect 31054 26238 31106 26290
rect 31390 26265 31442 26317
rect 31726 26238 31778 26290
rect 33630 26238 33682 26290
rect 35758 26265 35810 26317
rect 31166 26126 31218 26178
rect 36766 26126 36818 26178
rect 17614 26014 17666 26066
rect 5876 25846 5928 25898
rect 5980 25846 6032 25898
rect 6084 25846 6136 25898
rect 15200 25846 15252 25898
rect 15304 25846 15356 25898
rect 15408 25846 15460 25898
rect 24524 25846 24576 25898
rect 24628 25846 24680 25898
rect 24732 25846 24784 25898
rect 33848 25846 33900 25898
rect 33952 25846 34004 25898
rect 34056 25846 34108 25898
rect 4678 25678 4730 25730
rect 10726 25678 10778 25730
rect 13806 25678 13858 25730
rect 10166 25566 10218 25618
rect 15934 25622 15986 25674
rect 20078 25678 20130 25730
rect 20694 25678 20746 25730
rect 25174 25678 25226 25730
rect 18958 25566 19010 25618
rect 32958 25566 33010 25618
rect 3950 25454 4002 25506
rect 4958 25454 5010 25506
rect 5182 25454 5234 25506
rect 5948 25454 6000 25506
rect 6190 25454 6242 25506
rect 6694 25454 6746 25506
rect 7422 25454 7474 25506
rect 9662 25426 9714 25478
rect 10558 25454 10610 25506
rect 11006 25454 11058 25506
rect 12462 25454 12514 25506
rect 15262 25454 15314 25506
rect 15486 25454 15538 25506
rect 15822 25454 15874 25506
rect 18622 25454 18674 25506
rect 19352 25454 19404 25506
rect 19518 25454 19570 25506
rect 19630 25454 19682 25506
rect 20414 25454 20466 25506
rect 20526 25454 20578 25506
rect 24222 25454 24274 25506
rect 24782 25454 24834 25506
rect 25454 25454 25506 25506
rect 25678 25454 25730 25506
rect 26070 25454 26122 25506
rect 27694 25454 27746 25506
rect 28366 25454 28418 25506
rect 29598 25454 29650 25506
rect 29934 25454 29986 25506
rect 30494 25454 30546 25506
rect 30270 25398 30322 25450
rect 31278 25454 31330 25506
rect 31950 25454 32002 25506
rect 32510 25454 32562 25506
rect 33182 25454 33234 25506
rect 33518 25454 33570 25506
rect 34190 25454 34242 25506
rect 31502 25398 31554 25450
rect 32734 25398 32786 25450
rect 33854 25398 33906 25450
rect 35758 25454 35810 25506
rect 37326 25454 37378 25506
rect 37830 25510 37882 25562
rect 35366 25398 35418 25450
rect 35982 25398 36034 25450
rect 35534 25342 35586 25394
rect 2830 25230 2882 25282
rect 6638 25286 6690 25338
rect 4342 25230 4394 25282
rect 18118 25230 18170 25282
rect 18454 25230 18506 25282
rect 24110 25286 24162 25338
rect 21478 25230 21530 25282
rect 27918 25286 27970 25338
rect 29430 25286 29482 25338
rect 30606 25286 30658 25338
rect 31838 25286 31890 25338
rect 33630 25286 33682 25338
rect 37084 25342 37136 25394
rect 37998 25342 38050 25394
rect 26518 25230 26570 25282
rect 10538 25062 10590 25114
rect 10642 25062 10694 25114
rect 10746 25062 10798 25114
rect 19862 25062 19914 25114
rect 19966 25062 20018 25114
rect 20070 25062 20122 25114
rect 29186 25062 29238 25114
rect 29290 25062 29342 25114
rect 29394 25062 29446 25114
rect 38510 25062 38562 25114
rect 38614 25062 38666 25114
rect 38718 25062 38770 25114
rect 13078 24894 13130 24946
rect 14366 24894 14418 24946
rect 14702 24894 14754 24946
rect 15206 24894 15258 24946
rect 24614 24894 24666 24946
rect 30830 24894 30882 24946
rect 32174 24894 32226 24946
rect 33742 24894 33794 24946
rect 4734 24782 4786 24834
rect 5574 24782 5626 24834
rect 23998 24782 24050 24834
rect 2046 24670 2098 24722
rect 2830 24670 2882 24722
rect 5070 24670 5122 24722
rect 5294 24670 5346 24722
rect 7758 24670 7810 24722
rect 8318 24670 8370 24722
rect 6638 24558 6690 24610
rect 8822 24614 8874 24666
rect 8990 24670 9042 24722
rect 12686 24670 12738 24722
rect 15038 24670 15090 24722
rect 17614 24714 17666 24766
rect 18286 24726 18338 24778
rect 17838 24670 17890 24722
rect 18398 24698 18450 24750
rect 18678 24705 18730 24757
rect 18846 24726 18898 24778
rect 19518 24726 19570 24778
rect 19630 24698 19682 24750
rect 19910 24705 19962 24757
rect 20078 24726 20130 24778
rect 30158 24782 30210 24834
rect 34694 24782 34746 24834
rect 20358 24670 20410 24722
rect 20638 24670 20690 24722
rect 21310 24670 21362 24722
rect 29038 24670 29090 24722
rect 29262 24714 29314 24766
rect 29822 24670 29874 24722
rect 30494 24670 30546 24722
rect 31390 24670 31442 24722
rect 31614 24714 31666 24766
rect 32510 24670 32562 24722
rect 33406 24670 33458 24722
rect 34974 24670 35026 24722
rect 35198 24670 35250 24722
rect 37214 24670 37266 24722
rect 37886 24670 37938 24722
rect 17502 24558 17554 24610
rect 20974 24558 21026 24610
rect 22094 24558 22146 24610
rect 29374 24558 29426 24610
rect 31726 24558 31778 24610
rect 37550 24558 37602 24610
rect 38278 24558 38330 24610
rect 8076 24446 8128 24498
rect 12350 24446 12402 24498
rect 19126 24446 19178 24498
rect 25342 24446 25394 24498
rect 26238 24446 26290 24498
rect 26574 24446 26626 24498
rect 27134 24446 27186 24498
rect 27694 24446 27746 24498
rect 36094 24446 36146 24498
rect 5876 24278 5928 24330
rect 5980 24278 6032 24330
rect 6084 24278 6136 24330
rect 15200 24278 15252 24330
rect 15304 24278 15356 24330
rect 15408 24278 15460 24330
rect 24524 24278 24576 24330
rect 24628 24278 24680 24330
rect 24732 24278 24784 24330
rect 33848 24278 33900 24330
rect 33952 24278 34004 24330
rect 34056 24278 34108 24330
rect 3838 24110 3890 24162
rect 5742 24110 5794 24162
rect 18416 24110 18468 24162
rect 19574 24110 19626 24162
rect 20022 24110 20074 24162
rect 25342 24110 25394 24162
rect 32286 24110 32338 24162
rect 7198 23998 7250 24050
rect 10278 23998 10330 24050
rect 11510 23998 11562 24050
rect 4958 23886 5010 23938
rect 6078 23886 6130 23938
rect 9102 23886 9154 23938
rect 9886 23886 9938 23938
rect 12238 23886 12290 23938
rect 12742 23942 12794 23994
rect 12910 23886 12962 23938
rect 13638 23942 13690 23994
rect 14142 23886 14194 23938
rect 14702 23886 14754 23938
rect 16718 23886 16770 23938
rect 17502 23886 17554 23938
rect 17670 23942 17722 23994
rect 23886 23998 23938 24050
rect 24502 23998 24554 24050
rect 18174 23886 18226 23938
rect 18846 23886 18898 23938
rect 19014 23942 19066 23994
rect 26910 23998 26962 24050
rect 28142 24054 28194 24106
rect 29654 23998 29706 24050
rect 30830 24054 30882 24106
rect 30326 23998 30378 24050
rect 34582 23998 34634 24050
rect 34862 23998 34914 24050
rect 19182 23886 19234 23938
rect 19294 23886 19346 23938
rect 20302 23886 20354 23938
rect 20414 23886 20466 23938
rect 21198 23886 21250 23938
rect 21982 23886 22034 23938
rect 25678 23886 25730 23938
rect 26574 23886 26626 23938
rect 27246 23886 27298 23938
rect 11996 23774 12048 23826
rect 27022 23830 27074 23882
rect 27582 23886 27634 23938
rect 28254 23886 28306 23938
rect 28590 23886 28642 23938
rect 30718 23886 30770 23938
rect 30942 23886 30994 23938
rect 31838 23886 31890 23938
rect 31950 23886 32002 23938
rect 34974 23842 35026 23894
rect 35310 23886 35362 23938
rect 35646 23886 35698 23938
rect 35814 23942 35866 23994
rect 35982 23886 36034 23938
rect 36094 23886 36146 23938
rect 36374 23886 36426 23938
rect 37326 23886 37378 23938
rect 37830 23942 37882 23994
rect 37998 23886 38050 23938
rect 14384 23774 14436 23826
rect 6470 23662 6522 23714
rect 13582 23718 13634 23770
rect 37084 23774 37136 23826
rect 10838 23662 10890 23714
rect 15038 23662 15090 23714
rect 17054 23662 17106 23714
rect 31502 23662 31554 23714
rect 10538 23494 10590 23546
rect 10642 23494 10694 23546
rect 10746 23494 10798 23546
rect 19862 23494 19914 23546
rect 19966 23494 20018 23546
rect 20070 23494 20122 23546
rect 29186 23494 29238 23546
rect 29290 23494 29342 23546
rect 29394 23494 29446 23546
rect 38510 23494 38562 23546
rect 38614 23494 38666 23546
rect 38718 23494 38770 23546
rect 4286 23326 4338 23378
rect 8654 23326 8706 23378
rect 11118 23326 11170 23378
rect 15654 23326 15706 23378
rect 16606 23326 16658 23378
rect 20750 23326 20802 23378
rect 28646 23326 28698 23378
rect 37998 23326 38050 23378
rect 6246 23214 6298 23266
rect 10558 23214 10610 23266
rect 14254 23214 14306 23266
rect 18342 23214 18394 23266
rect 18790 23214 18842 23266
rect 20078 23214 20130 23266
rect 36412 23214 36464 23266
rect 4622 23102 4674 23154
rect 6582 23102 6634 23154
rect 6862 23102 6914 23154
rect 7086 23102 7138 23154
rect 7198 23102 7250 23154
rect 9886 23102 9938 23154
rect 5014 22990 5066 23042
rect 10390 23046 10442 23098
rect 10782 23102 10834 23154
rect 11566 23102 11618 23154
rect 12350 23102 12402 23154
rect 14590 23102 14642 23154
rect 14814 23102 14866 23154
rect 16942 23102 16994 23154
rect 17950 23102 18002 23154
rect 18062 23102 18114 23154
rect 19070 23102 19122 23154
rect 19294 23102 19346 23154
rect 19742 23102 19794 23154
rect 20414 23102 20466 23154
rect 22430 23102 22482 23154
rect 22766 23102 22818 23154
rect 25566 23102 25618 23154
rect 26350 23102 26402 23154
rect 27134 23102 27186 23154
rect 27806 23158 27858 23210
rect 37326 23214 37378 23266
rect 27470 23102 27522 23154
rect 28030 23102 28082 23154
rect 29038 23102 29090 23154
rect 29262 23102 29314 23154
rect 29822 23146 29874 23198
rect 30158 23102 30210 23154
rect 30494 23102 30546 23154
rect 31054 23102 31106 23154
rect 31614 23102 31666 23154
rect 32286 23102 32338 23154
rect 34526 23102 34578 23154
rect 35422 23102 35474 23154
rect 35758 23102 35810 23154
rect 37158 23158 37210 23210
rect 36654 23102 36706 23154
rect 38334 23102 38386 23154
rect 16102 22990 16154 23042
rect 22318 22934 22370 22986
rect 25342 22990 25394 23042
rect 27918 22990 27970 23042
rect 29710 22990 29762 23042
rect 29038 22934 29090 22986
rect 31278 22934 31330 22986
rect 32398 22934 32450 22986
rect 9644 22878 9696 22930
rect 15094 22878 15146 22930
rect 34862 22878 34914 22930
rect 5876 22710 5928 22762
rect 5980 22710 6032 22762
rect 6084 22710 6136 22762
rect 15200 22710 15252 22762
rect 15304 22710 15356 22762
rect 15408 22710 15460 22762
rect 24524 22710 24576 22762
rect 24628 22710 24680 22762
rect 24732 22710 24784 22762
rect 33848 22710 33900 22762
rect 33952 22710 34004 22762
rect 34056 22710 34108 22762
rect 12406 22542 12458 22594
rect 19966 22542 20018 22594
rect 11006 22430 11058 22482
rect 18734 22430 18786 22482
rect 19462 22430 19514 22482
rect 29150 22486 29202 22538
rect 26014 22430 26066 22482
rect 27918 22430 27970 22482
rect 31502 22486 31554 22538
rect 32174 22430 32226 22482
rect 38278 22430 38330 22482
rect 2942 22318 2994 22370
rect 3166 22318 3218 22370
rect 5182 22318 5234 22370
rect 7982 22318 8034 22370
rect 8206 22318 8258 22370
rect 8318 22318 8370 22370
rect 9102 22318 9154 22370
rect 11902 22318 11954 22370
rect 12126 22318 12178 22370
rect 14030 22318 14082 22370
rect 15486 22318 15538 22370
rect 16046 22318 16098 22370
rect 16830 22318 16882 22370
rect 19630 22318 19682 22370
rect 23214 22318 23266 22370
rect 23438 22318 23490 22370
rect 23718 22318 23770 22370
rect 25678 22318 25730 22370
rect 26350 22318 26402 22370
rect 27582 22318 27634 22370
rect 28142 22318 28194 22370
rect 29262 22318 29314 22370
rect 29486 22318 29538 22370
rect 30494 22318 30546 22370
rect 26126 22262 26178 22314
rect 30714 22280 30766 22332
rect 31390 22318 31442 22370
rect 31838 22318 31890 22370
rect 32510 22318 32562 22370
rect 32174 22262 32226 22314
rect 32846 22318 32898 22370
rect 33406 22318 33458 22370
rect 34078 22318 34130 22370
rect 33574 22262 33626 22314
rect 34638 22318 34690 22370
rect 34862 22318 34914 22370
rect 2662 22206 2714 22258
rect 4062 22206 4114 22258
rect 7702 22206 7754 22258
rect 34320 22206 34372 22258
rect 35142 22206 35194 22258
rect 5798 22094 5850 22146
rect 7366 22094 7418 22146
rect 30158 22094 30210 22146
rect 10538 21926 10590 21978
rect 10642 21926 10694 21978
rect 10746 21926 10798 21978
rect 19862 21926 19914 21978
rect 19966 21926 20018 21978
rect 20070 21926 20122 21978
rect 29186 21926 29238 21978
rect 29290 21926 29342 21978
rect 29394 21926 29446 21978
rect 38510 21926 38562 21978
rect 38614 21926 38666 21978
rect 38718 21926 38770 21978
rect 6694 21758 6746 21810
rect 15878 21758 15930 21810
rect 18342 21758 18394 21810
rect 19070 21758 19122 21810
rect 5276 21646 5328 21698
rect 6190 21646 6242 21698
rect 2046 21534 2098 21586
rect 6022 21590 6074 21642
rect 12686 21646 12738 21698
rect 33350 21646 33402 21698
rect 5518 21534 5570 21586
rect 11566 21534 11618 21586
rect 11790 21534 11842 21586
rect 13806 21534 13858 21586
rect 14478 21534 14530 21586
rect 18174 21534 18226 21586
rect 19406 21534 19458 21586
rect 19798 21534 19850 21586
rect 21646 21534 21698 21586
rect 25230 21534 25282 21586
rect 25510 21563 25562 21615
rect 26126 21534 26178 21586
rect 26574 21573 26626 21625
rect 26798 21534 26850 21586
rect 27134 21534 27186 21586
rect 27582 21534 27634 21586
rect 30382 21590 30434 21642
rect 31950 21590 32002 21642
rect 27806 21534 27858 21586
rect 28590 21534 28642 21586
rect 28926 21534 28978 21586
rect 30158 21534 30210 21586
rect 30718 21534 30770 21586
rect 31614 21534 31666 21586
rect 32286 21534 32338 21586
rect 33630 21534 33682 21586
rect 33742 21534 33794 21586
rect 33966 21534 34018 21586
rect 35982 21534 36034 21586
rect 2830 21422 2882 21474
rect 4734 21422 4786 21474
rect 8374 21422 8426 21474
rect 24054 21422 24106 21474
rect 25678 21422 25730 21474
rect 26238 21422 26290 21474
rect 28086 21422 28138 21474
rect 30606 21422 30658 21474
rect 31334 21422 31386 21474
rect 11286 21310 11338 21362
rect 14142 21310 14194 21362
rect 21982 21310 22034 21362
rect 28478 21366 28530 21418
rect 31950 21422 32002 21474
rect 35422 21310 35474 21362
rect 37438 21310 37490 21362
rect 5876 21142 5928 21194
rect 5980 21142 6032 21194
rect 6084 21142 6136 21194
rect 15200 21142 15252 21194
rect 15304 21142 15356 21194
rect 15408 21142 15460 21194
rect 24524 21142 24576 21194
rect 24628 21142 24680 21194
rect 24732 21142 24784 21194
rect 33848 21142 33900 21194
rect 33952 21142 34004 21194
rect 34056 21142 34108 21194
rect 3166 20974 3218 21026
rect 9326 20974 9378 21026
rect 13564 20974 13616 21026
rect 19406 20974 19458 21026
rect 22094 20974 22146 21026
rect 24838 20974 24890 21026
rect 37904 20974 37956 21026
rect 25678 20918 25730 20970
rect 2046 20750 2098 20802
rect 4958 20750 5010 20802
rect 5182 20750 5234 20802
rect 5724 20750 5776 20802
rect 5966 20750 6018 20802
rect 6470 20806 6522 20858
rect 20190 20862 20242 20914
rect 35758 20862 35810 20914
rect 6638 20750 6690 20802
rect 7310 20750 7362 20802
rect 7814 20750 7866 20802
rect 8206 20750 8258 20802
rect 11118 20750 11170 20802
rect 13806 20750 13858 20802
rect 14478 20750 14530 20802
rect 4678 20638 4730 20690
rect 7068 20638 7120 20690
rect 14310 20694 14362 20746
rect 19070 20750 19122 20802
rect 19854 20750 19906 20802
rect 20526 20750 20578 20802
rect 20302 20694 20354 20746
rect 23774 20722 23826 20774
rect 24110 20750 24162 20802
rect 24558 20750 24610 20802
rect 25566 20750 25618 20802
rect 25790 20750 25842 20802
rect 26126 20750 26178 20802
rect 24278 20694 24330 20746
rect 30326 20750 30378 20802
rect 31390 20750 31442 20802
rect 32062 20750 32114 20802
rect 32286 20750 32338 20802
rect 33854 20750 33906 20802
rect 36542 20750 36594 20802
rect 36990 20750 37042 20802
rect 37158 20750 37210 20802
rect 37662 20750 37714 20802
rect 7982 20638 8034 20690
rect 24446 20638 24498 20690
rect 31726 20638 31778 20690
rect 32566 20638 32618 20690
rect 12574 20526 12626 20578
rect 14982 20526 15034 20578
rect 15318 20526 15370 20578
rect 15934 20526 15986 20578
rect 26462 20526 26514 20578
rect 27078 20526 27130 20578
rect 10538 20358 10590 20410
rect 10642 20358 10694 20410
rect 10746 20358 10798 20410
rect 19862 20358 19914 20410
rect 19966 20358 20018 20410
rect 20070 20358 20122 20410
rect 29186 20358 29238 20410
rect 29290 20358 29342 20410
rect 29394 20358 29446 20410
rect 38510 20358 38562 20410
rect 38614 20358 38666 20410
rect 38718 20358 38770 20410
rect 6862 20078 6914 20130
rect 7310 20078 7362 20130
rect 9606 20134 9658 20186
rect 15318 20190 15370 20242
rect 14702 20078 14754 20130
rect 19910 20134 19962 20186
rect 25846 20190 25898 20242
rect 3838 19966 3890 20018
rect 4062 19966 4114 20018
rect 7478 20022 7530 20074
rect 33294 20078 33346 20130
rect 4174 19966 4226 20018
rect 7982 19966 8034 20018
rect 9438 19966 9490 20018
rect 12014 19966 12066 20018
rect 12798 19966 12850 20018
rect 20078 19966 20130 20018
rect 20302 20001 20354 20053
rect 20414 19994 20466 20046
rect 20638 19994 20690 20046
rect 20912 19994 20964 20046
rect 21422 19966 21474 20018
rect 22878 19966 22930 20018
rect 23438 19966 23490 20018
rect 24110 19966 24162 20018
rect 25454 19966 25506 20018
rect 29038 19966 29090 20018
rect 30270 20022 30322 20074
rect 34208 20078 34260 20130
rect 29262 19966 29314 20018
rect 29542 19966 29594 20018
rect 29934 19966 29986 20018
rect 30606 19966 30658 20018
rect 30942 19966 30994 20018
rect 31390 19966 31442 20018
rect 33462 20022 33514 20074
rect 35646 20078 35698 20130
rect 31614 19966 31666 20018
rect 33966 19966 34018 20018
rect 37550 19966 37602 20018
rect 38334 19966 38386 20018
rect 4958 19854 5010 19906
rect 15766 19854 15818 19906
rect 30270 19854 30322 19906
rect 31894 19854 31946 19906
rect 35254 19854 35306 19906
rect 3558 19742 3610 19794
rect 8224 19742 8276 19794
rect 21142 19742 21194 19794
rect 23774 19742 23826 19794
rect 24446 19742 24498 19794
rect 25286 19742 25338 19794
rect 5876 19574 5928 19626
rect 5980 19574 6032 19626
rect 6084 19574 6136 19626
rect 15200 19574 15252 19626
rect 15304 19574 15356 19626
rect 15408 19574 15460 19626
rect 24524 19574 24576 19626
rect 24628 19574 24680 19626
rect 24732 19574 24784 19626
rect 33848 19574 33900 19626
rect 33952 19574 34004 19626
rect 34056 19574 34108 19626
rect 4734 19406 4786 19458
rect 21366 19406 21418 19458
rect 21814 19406 21866 19458
rect 29486 19406 29538 19458
rect 29990 19406 30042 19458
rect 37998 19406 38050 19458
rect 10670 19294 10722 19346
rect 17166 19294 17218 19346
rect 23102 19294 23154 19346
rect 3278 19182 3330 19234
rect 5518 19182 5570 19234
rect 7982 19182 8034 19234
rect 8766 19182 8818 19234
rect 11902 19182 11954 19234
rect 12574 19182 12626 19234
rect 13414 19238 13466 19290
rect 25006 19294 25058 19346
rect 13806 19182 13858 19234
rect 12070 19126 12122 19178
rect 14142 19144 14194 19196
rect 14478 19182 14530 19234
rect 15262 19182 15314 19234
rect 17782 19182 17834 19234
rect 18846 19182 18898 19234
rect 19518 19182 19570 19234
rect 19966 19182 20018 19234
rect 20526 19182 20578 19234
rect 21534 19182 21586 19234
rect 21982 19182 22034 19234
rect 22430 19182 22482 19234
rect 12816 19070 12868 19122
rect 19070 19126 19122 19178
rect 20190 19126 20242 19178
rect 22766 19182 22818 19234
rect 22990 19143 23042 19195
rect 23438 19182 23490 19234
rect 23774 19182 23826 19234
rect 23998 19182 24050 19234
rect 24782 19182 24834 19234
rect 25342 19182 25394 19234
rect 25902 19182 25954 19234
rect 26574 19182 26626 19234
rect 25006 19126 25058 19178
rect 26350 19126 26402 19178
rect 27022 19182 27074 19234
rect 27246 19182 27298 19234
rect 29150 19182 29202 19234
rect 30270 19182 30322 19234
rect 30382 19182 30434 19234
rect 30550 19182 30602 19234
rect 31054 19238 31106 19290
rect 31894 19238 31946 19290
rect 32342 19294 32394 19346
rect 37158 19294 37210 19346
rect 30718 19182 30770 19234
rect 31166 19144 31218 19196
rect 37606 19182 37658 19234
rect 38334 19182 38386 19234
rect 13582 19070 13634 19122
rect 24278 19070 24330 19122
rect 27526 19070 27578 19122
rect 31726 19070 31778 19122
rect 6638 18958 6690 19010
rect 7814 18958 7866 19010
rect 19406 19014 19458 19066
rect 20638 19014 20690 19066
rect 26686 19014 26738 19066
rect 11286 18958 11338 19010
rect 10538 18790 10590 18842
rect 10642 18790 10694 18842
rect 10746 18790 10798 18842
rect 19862 18790 19914 18842
rect 19966 18790 20018 18842
rect 20070 18790 20122 18842
rect 29186 18790 29238 18842
rect 29290 18790 29342 18842
rect 29394 18790 29446 18842
rect 38510 18790 38562 18842
rect 38614 18790 38666 18842
rect 38718 18790 38770 18842
rect 15262 18622 15314 18674
rect 8430 18510 8482 18562
rect 12462 18510 12514 18562
rect 5742 18398 5794 18450
rect 6526 18398 6578 18450
rect 9046 18398 9098 18450
rect 9438 18398 9490 18450
rect 9662 18398 9714 18450
rect 11006 18398 11058 18450
rect 11118 18398 11170 18450
rect 12294 18454 12346 18506
rect 19966 18510 20018 18562
rect 23382 18510 23434 18562
rect 29486 18510 29538 18562
rect 11790 18398 11842 18450
rect 12910 18398 12962 18450
rect 13134 18398 13186 18450
rect 13414 18398 13466 18450
rect 13806 18398 13858 18450
rect 21982 18454 22034 18506
rect 17278 18398 17330 18450
rect 20414 18398 20466 18450
rect 20750 18398 20802 18450
rect 21198 18398 21250 18450
rect 21534 18398 21586 18450
rect 22094 18426 22146 18478
rect 22318 18426 22370 18478
rect 22542 18426 22594 18478
rect 23662 18398 23714 18450
rect 23774 18398 23826 18450
rect 24110 18398 24162 18450
rect 25902 18454 25954 18506
rect 24334 18398 24386 18450
rect 24614 18398 24666 18450
rect 25566 18398 25618 18450
rect 26238 18398 26290 18450
rect 26686 18398 26738 18450
rect 26910 18398 26962 18450
rect 28030 18398 28082 18450
rect 29374 18398 29426 18450
rect 18062 18286 18114 18338
rect 20302 18286 20354 18338
rect 22822 18286 22874 18338
rect 25902 18286 25954 18338
rect 27694 18286 27746 18338
rect 29654 18342 29706 18394
rect 29822 18398 29874 18450
rect 30270 18398 30322 18450
rect 31010 18436 31062 18488
rect 31166 18398 31218 18450
rect 33966 18398 34018 18450
rect 34190 18398 34242 18450
rect 34470 18398 34522 18450
rect 34750 18398 34802 18450
rect 35758 18398 35810 18450
rect 9942 18174 9994 18226
rect 10726 18174 10778 18226
rect 11548 18174 11600 18226
rect 27190 18174 27242 18226
rect 29094 18174 29146 18226
rect 30158 18230 30210 18282
rect 31334 18230 31386 18282
rect 33798 18286 33850 18338
rect 35086 18174 35138 18226
rect 35926 18230 35978 18282
rect 5876 18006 5928 18058
rect 5980 18006 6032 18058
rect 6084 18006 6136 18058
rect 15200 18006 15252 18058
rect 15304 18006 15356 18058
rect 15408 18006 15460 18058
rect 24524 18006 24576 18058
rect 24628 18006 24680 18058
rect 24732 18006 24784 18058
rect 33848 18006 33900 18058
rect 33952 18006 34004 18058
rect 34056 18006 34108 18058
rect 8542 17838 8594 17890
rect 17838 17838 17890 17890
rect 24334 17782 24386 17834
rect 12686 17726 12738 17778
rect 9662 17614 9714 17666
rect 9998 17614 10050 17666
rect 10782 17614 10834 17666
rect 13358 17614 13410 17666
rect 13582 17614 13634 17666
rect 14142 17614 14194 17666
rect 15094 17614 15146 17666
rect 18174 17614 18226 17666
rect 20750 17614 20802 17666
rect 23886 17614 23938 17666
rect 24222 17614 24274 17666
rect 25174 17614 25226 17666
rect 27078 17670 27130 17722
rect 28646 17726 28698 17778
rect 30494 17726 30546 17778
rect 31110 17726 31162 17778
rect 34414 17726 34466 17778
rect 37158 17726 37210 17778
rect 25454 17614 25506 17666
rect 25566 17614 25618 17666
rect 25902 17614 25954 17666
rect 25734 17558 25786 17610
rect 26462 17586 26514 17638
rect 26686 17614 26738 17666
rect 29374 17614 29426 17666
rect 29822 17614 29874 17666
rect 29934 17614 29986 17666
rect 13862 17502 13914 17554
rect 20022 17502 20074 17554
rect 30100 17558 30152 17610
rect 33686 17588 33738 17640
rect 38334 17614 38386 17666
rect 26910 17502 26962 17554
rect 36318 17502 36370 17554
rect 14478 17390 14530 17442
rect 20414 17390 20466 17442
rect 27470 17390 27522 17442
rect 27806 17390 27858 17442
rect 29206 17390 29258 17442
rect 37606 17390 37658 17442
rect 37998 17390 38050 17442
rect 10538 17222 10590 17274
rect 10642 17222 10694 17274
rect 10746 17222 10798 17274
rect 19862 17222 19914 17274
rect 19966 17222 20018 17274
rect 20070 17222 20122 17274
rect 29186 17222 29238 17274
rect 29290 17222 29342 17274
rect 29394 17222 29446 17274
rect 38510 17222 38562 17274
rect 38614 17222 38666 17274
rect 38718 17222 38770 17274
rect 9718 17054 9770 17106
rect 11006 17054 11058 17106
rect 17558 17054 17610 17106
rect 12350 16942 12402 16994
rect 13264 16942 13316 16994
rect 8654 16830 8706 16882
rect 8990 16830 9042 16882
rect 12518 16886 12570 16938
rect 20078 16998 20130 17050
rect 22486 16998 22538 17050
rect 23046 17054 23098 17106
rect 28142 17054 28194 17106
rect 31110 17054 31162 17106
rect 33686 17054 33738 17106
rect 16382 16942 16434 16994
rect 25902 16942 25954 16994
rect 9886 16830 9938 16882
rect 13022 16830 13074 16882
rect 13694 16830 13746 16882
rect 18790 16830 18842 16882
rect 20414 16886 20466 16938
rect 19294 16830 19346 16882
rect 19966 16830 20018 16882
rect 20526 16858 20578 16910
rect 20750 16886 20802 16938
rect 20974 16886 21026 16938
rect 21254 16830 21306 16882
rect 21758 16874 21810 16926
rect 21982 16830 22034 16882
rect 22318 16830 22370 16882
rect 23550 16830 23602 16882
rect 23662 16830 23714 16882
rect 25734 16886 25786 16938
rect 25566 16830 25618 16882
rect 26014 16830 26066 16882
rect 26294 16830 26346 16882
rect 27806 16830 27858 16882
rect 28590 16830 28642 16882
rect 28926 16830 28978 16882
rect 29554 16870 29606 16922
rect 29710 16866 29762 16918
rect 30158 16866 30210 16918
rect 30494 16886 30546 16938
rect 34414 16830 34466 16882
rect 34526 16830 34578 16882
rect 14478 16718 14530 16770
rect 21646 16718 21698 16770
rect 29486 16718 29538 16770
rect 34078 16718 34130 16770
rect 35310 16718 35362 16770
rect 37214 16718 37266 16770
rect 29038 16662 29090 16714
rect 23942 16606 23994 16658
rect 5876 16438 5928 16490
rect 5980 16438 6032 16490
rect 6084 16438 6136 16490
rect 15200 16438 15252 16490
rect 15304 16438 15356 16490
rect 15408 16438 15460 16490
rect 24524 16438 24576 16490
rect 24628 16438 24680 16490
rect 24732 16438 24784 16490
rect 33848 16438 33900 16490
rect 33952 16438 34004 16490
rect 34056 16438 34108 16490
rect 14478 16270 14530 16322
rect 18398 16270 18450 16322
rect 22224 16270 22276 16322
rect 19630 16214 19682 16266
rect 22766 16270 22818 16322
rect 35068 16270 35120 16322
rect 37382 16270 37434 16322
rect 20638 16158 20690 16210
rect 27414 16158 27466 16210
rect 28366 16158 28418 16210
rect 31390 16158 31442 16210
rect 32006 16158 32058 16210
rect 33798 16158 33850 16210
rect 36486 16158 36538 16210
rect 11342 16046 11394 16098
rect 11734 16046 11786 16098
rect 13358 16046 13410 16098
rect 15374 16046 15426 16098
rect 18062 16046 18114 16098
rect 18846 16046 18898 16098
rect 19518 16046 19570 16098
rect 20414 16046 20466 16098
rect 20246 15990 20298 16042
rect 20806 15990 20858 16042
rect 21310 16046 21362 16098
rect 21982 16046 22034 16098
rect 21478 15990 21530 16042
rect 23102 16046 23154 16098
rect 24577 16046 24629 16098
rect 25454 16046 25506 16098
rect 27918 16046 27970 16098
rect 28590 16046 28642 16098
rect 11006 15934 11058 15986
rect 28254 15990 28306 16042
rect 29330 16013 29382 16065
rect 29486 16009 29538 16061
rect 29934 16009 29986 16061
rect 30382 16013 30434 16065
rect 30718 16046 30770 16098
rect 30830 16046 30882 16098
rect 30996 16046 31048 16098
rect 32846 16046 32898 16098
rect 34526 16046 34578 16098
rect 35310 16046 35362 16098
rect 36878 16046 36930 16098
rect 24334 15934 24386 15986
rect 35814 15990 35866 16042
rect 37102 16046 37154 16098
rect 29150 15934 29202 15986
rect 35982 15934 36034 15986
rect 15710 15822 15762 15874
rect 23494 15822 23546 15874
rect 33182 15822 33234 15874
rect 34190 15822 34242 15874
rect 10538 15654 10590 15706
rect 10642 15654 10694 15706
rect 10746 15654 10798 15706
rect 19862 15654 19914 15706
rect 19966 15654 20018 15706
rect 20070 15654 20122 15706
rect 29186 15654 29238 15706
rect 29290 15654 29342 15706
rect 29394 15654 29446 15706
rect 38510 15654 38562 15706
rect 38614 15654 38666 15706
rect 38718 15654 38770 15706
rect 12126 15486 12178 15538
rect 15206 15486 15258 15538
rect 23326 15486 23378 15538
rect 23942 15486 23994 15538
rect 25510 15486 25562 15538
rect 26014 15486 26066 15538
rect 26350 15486 26402 15538
rect 19966 15374 20018 15426
rect 21758 15374 21810 15426
rect 22672 15374 22724 15426
rect 27470 15374 27522 15426
rect 31502 15374 31554 15426
rect 33854 15374 33906 15426
rect 35292 15374 35344 15426
rect 36206 15374 36258 15426
rect 12462 15262 12514 15314
rect 17278 15262 17330 15314
rect 18062 15262 18114 15314
rect 21124 15300 21176 15352
rect 21310 15262 21362 15314
rect 21422 15262 21474 15314
rect 20750 15150 20802 15202
rect 21926 15206 21978 15258
rect 22430 15262 22482 15314
rect 22990 15262 23042 15314
rect 25342 15262 25394 15314
rect 24390 15150 24442 15202
rect 27638 15206 27690 15258
rect 28142 15262 28194 15314
rect 28814 15262 28866 15314
rect 29598 15262 29650 15314
rect 32958 15262 33010 15314
rect 32342 15150 32394 15202
rect 34022 15206 34074 15258
rect 34526 15262 34578 15314
rect 35534 15262 35586 15314
rect 36038 15206 36090 15258
rect 28384 15038 28436 15090
rect 34768 15038 34820 15090
rect 5876 14870 5928 14922
rect 5980 14870 6032 14922
rect 6084 14870 6136 14922
rect 15200 14870 15252 14922
rect 15304 14870 15356 14922
rect 15408 14870 15460 14922
rect 24524 14870 24576 14922
rect 24628 14870 24680 14922
rect 24732 14870 24784 14922
rect 33848 14870 33900 14922
rect 33952 14870 34004 14922
rect 34056 14870 34108 14922
rect 11510 14702 11562 14754
rect 13582 14702 13634 14754
rect 20582 14702 20634 14754
rect 36336 14702 36388 14754
rect 12070 14590 12122 14642
rect 17726 14590 17778 14642
rect 19630 14590 19682 14642
rect 24502 14590 24554 14642
rect 27078 14590 27130 14642
rect 29318 14590 29370 14642
rect 33630 14590 33682 14642
rect 37158 14590 37210 14642
rect 7086 14478 7138 14530
rect 7870 14478 7922 14530
rect 10894 14478 10946 14530
rect 11006 14478 11058 14530
rect 11230 14478 11282 14530
rect 13918 14478 13970 14530
rect 16942 14478 16994 14530
rect 20078 14478 20130 14530
rect 20302 14478 20354 14530
rect 21310 14478 21362 14530
rect 21982 14478 22034 14530
rect 21478 14422 21530 14474
rect 22224 14478 22276 14530
rect 22654 14478 22706 14530
rect 23326 14478 23378 14530
rect 23102 14422 23154 14474
rect 25118 14478 25170 14530
rect 25342 14478 25394 14530
rect 25902 14478 25954 14530
rect 26574 14478 26626 14530
rect 26406 14422 26458 14474
rect 28590 14478 28642 14530
rect 31502 14478 31554 14530
rect 32622 14450 32674 14502
rect 36094 14478 36146 14530
rect 9774 14366 9826 14418
rect 24838 14366 24890 14418
rect 25660 14366 25712 14418
rect 10558 14254 10610 14306
rect 22766 14310 22818 14362
rect 35590 14422 35642 14474
rect 38334 14478 38386 14530
rect 35422 14366 35474 14418
rect 37998 14366 38050 14418
rect 14310 14254 14362 14306
rect 24054 14254 24106 14306
rect 28254 14254 28306 14306
rect 31838 14254 31890 14306
rect 37606 14254 37658 14306
rect 10538 14086 10590 14138
rect 10642 14086 10694 14138
rect 10746 14086 10798 14138
rect 19862 14086 19914 14138
rect 19966 14086 20018 14138
rect 20070 14086 20122 14138
rect 29186 14086 29238 14138
rect 29290 14086 29342 14138
rect 29394 14086 29446 14138
rect 38510 14086 38562 14138
rect 38614 14086 38666 14138
rect 38718 14086 38770 14138
rect 7982 13918 8034 13970
rect 15094 13918 15146 13970
rect 18006 13918 18058 13970
rect 23942 13918 23994 13970
rect 19630 13806 19682 13858
rect 21310 13806 21362 13858
rect 22318 13806 22370 13858
rect 29934 13806 29986 13858
rect 36300 13806 36352 13858
rect 9102 13694 9154 13746
rect 9998 13694 10050 13746
rect 10502 13638 10554 13690
rect 10670 13694 10722 13746
rect 14142 13694 14194 13746
rect 16494 13694 16546 13746
rect 18174 13694 18226 13746
rect 20190 13694 20242 13746
rect 11454 13582 11506 13634
rect 13358 13582 13410 13634
rect 14534 13582 14586 13634
rect 22486 13638 22538 13690
rect 22990 13694 23042 13746
rect 23232 13694 23284 13746
rect 23774 13694 23826 13746
rect 25678 13694 25730 13746
rect 25790 13694 25842 13746
rect 27246 13694 27298 13746
rect 28030 13694 28082 13746
rect 31278 13694 31330 13746
rect 31390 13694 31442 13746
rect 32174 13694 32226 13746
rect 33070 13694 33122 13746
rect 33854 13694 33906 13746
rect 35758 13694 35810 13746
rect 37046 13750 37098 13802
rect 36542 13694 36594 13746
rect 37214 13694 37266 13746
rect 37438 13694 37490 13746
rect 24502 13582 24554 13634
rect 30662 13582 30714 13634
rect 9756 13470 9808 13522
rect 16158 13470 16210 13522
rect 25342 13470 25394 13522
rect 26126 13470 26178 13522
rect 30998 13470 31050 13522
rect 31838 13470 31890 13522
rect 37774 13470 37826 13522
rect 5876 13302 5928 13354
rect 5980 13302 6032 13354
rect 6084 13302 6136 13354
rect 15200 13302 15252 13354
rect 15304 13302 15356 13354
rect 15408 13302 15460 13354
rect 24524 13302 24576 13354
rect 24628 13302 24680 13354
rect 24732 13302 24784 13354
rect 33848 13302 33900 13354
rect 33952 13302 34004 13354
rect 34056 13302 34108 13354
rect 8598 13134 8650 13186
rect 10502 13134 10554 13186
rect 12574 13134 12626 13186
rect 19406 13134 19458 13186
rect 22430 13134 22482 13186
rect 36374 13134 36426 13186
rect 13638 13022 13690 13074
rect 14198 13022 14250 13074
rect 15822 13022 15874 13074
rect 22878 13022 22930 13074
rect 24334 13022 24386 13074
rect 26238 13022 26290 13074
rect 8878 12910 8930 12962
rect 9102 12910 9154 12962
rect 10222 12910 10274 12962
rect 10782 12910 10834 12962
rect 11006 12910 11058 12962
rect 11118 12910 11170 12962
rect 14366 12910 14418 12962
rect 15038 12910 15090 12962
rect 17726 12910 17778 12962
rect 20862 12910 20914 12962
rect 21310 12910 21362 12962
rect 22186 12854 22238 12906
rect 22990 12895 23042 12947
rect 23214 12910 23266 12962
rect 23550 12910 23602 12962
rect 28702 12910 28754 12962
rect 29598 12910 29650 12962
rect 29934 12910 29986 12962
rect 30046 12910 30098 12962
rect 30830 12910 30882 12962
rect 33182 12910 33234 12962
rect 33854 12910 33906 12962
rect 18342 12798 18394 12850
rect 33350 12854 33402 12906
rect 34638 12910 34690 12962
rect 35310 12910 35362 12962
rect 32734 12798 32786 12850
rect 34806 12854 34858 12906
rect 35552 12910 35604 12962
rect 35870 12910 35922 12962
rect 36094 12910 36146 12962
rect 36990 12910 37042 12962
rect 37158 12910 37210 12962
rect 37662 12910 37714 12962
rect 34096 12798 34148 12850
rect 37904 12798 37956 12850
rect 7814 12686 7866 12738
rect 9550 12686 9602 12738
rect 14702 12686 14754 12738
rect 10538 12518 10590 12570
rect 10642 12518 10694 12570
rect 10746 12518 10798 12570
rect 19862 12518 19914 12570
rect 19966 12518 20018 12570
rect 20070 12518 20122 12570
rect 29186 12518 29238 12570
rect 29290 12518 29342 12570
rect 29394 12518 29446 12570
rect 38510 12518 38562 12570
rect 38614 12518 38666 12570
rect 38718 12518 38770 12570
rect 7310 12350 7362 12402
rect 15094 12350 15146 12402
rect 11902 12294 11954 12346
rect 22934 12350 22986 12402
rect 23382 12350 23434 12402
rect 33910 12350 33962 12402
rect 35254 12350 35306 12402
rect 10670 12238 10722 12290
rect 16214 12238 16266 12290
rect 18062 12238 18114 12290
rect 22318 12238 22370 12290
rect 27806 12238 27858 12290
rect 31166 12238 31218 12290
rect 32080 12238 32132 12290
rect 34246 12238 34298 12290
rect 35646 12238 35698 12290
rect 7646 12126 7698 12178
rect 7870 12126 7922 12178
rect 8038 12126 8090 12178
rect 8542 12126 8594 12178
rect 9606 12126 9658 12178
rect 9886 12126 9938 12178
rect 9998 12126 10050 12178
rect 11006 12126 11058 12178
rect 11566 12126 11618 12178
rect 12070 12126 12122 12178
rect 13806 12126 13858 12178
rect 14086 12126 14138 12178
rect 14366 12126 14418 12178
rect 14590 12126 14642 12178
rect 15262 12126 15314 12178
rect 16494 12126 16546 12178
rect 16718 12126 16770 12178
rect 19182 12126 19234 12178
rect 19630 12126 19682 12178
rect 20414 12126 20466 12178
rect 25118 12126 25170 12178
rect 25902 12126 25954 12178
rect 28590 12153 28642 12205
rect 11324 12014 11376 12066
rect 12742 12014 12794 12066
rect 13134 12014 13186 12066
rect 31334 12070 31386 12122
rect 31838 12126 31890 12178
rect 34526 12126 34578 12178
rect 34638 12126 34690 12178
rect 37550 12126 37602 12178
rect 38334 12126 38386 12178
rect 8784 11902 8836 11954
rect 29374 11902 29426 11954
rect 5876 11734 5928 11786
rect 5980 11734 6032 11786
rect 6084 11734 6136 11786
rect 15200 11734 15252 11786
rect 15304 11734 15356 11786
rect 15408 11734 15460 11786
rect 24524 11734 24576 11786
rect 24628 11734 24680 11786
rect 24732 11734 24784 11786
rect 33848 11734 33900 11786
rect 33952 11734 34004 11786
rect 34056 11734 34108 11786
rect 22430 11566 22482 11618
rect 37998 11566 38050 11618
rect 14590 11454 14642 11506
rect 17670 11454 17722 11506
rect 23046 11454 23098 11506
rect 28086 11454 28138 11506
rect 5854 11342 5906 11394
rect 6638 11342 6690 11394
rect 9326 11342 9378 11394
rect 9438 11342 9490 11394
rect 9998 11342 10050 11394
rect 10110 11342 10162 11394
rect 10390 11342 10442 11394
rect 10670 11342 10722 11394
rect 11902 11342 11954 11394
rect 12070 11342 12122 11394
rect 12574 11342 12626 11394
rect 12816 11342 12868 11394
rect 14030 11342 14082 11394
rect 14142 11342 14194 11394
rect 16494 11342 16546 11394
rect 17278 11342 17330 11394
rect 17950 11342 18002 11394
rect 18734 11342 18786 11394
rect 20638 11342 20690 11394
rect 21310 11342 21362 11394
rect 22186 11342 22238 11394
rect 26350 11342 26402 11394
rect 26574 11342 26626 11394
rect 27246 11342 27298 11394
rect 30046 11342 30098 11394
rect 30158 11342 30210 11394
rect 38334 11342 38386 11394
rect 8542 11230 8594 11282
rect 9046 11230 9098 11282
rect 13750 11230 13802 11282
rect 26070 11230 26122 11282
rect 37606 11230 37658 11282
rect 26910 11118 26962 11170
rect 29710 11118 29762 11170
rect 30494 11118 30546 11170
rect 35254 11118 35306 11170
rect 10538 10950 10590 11002
rect 10642 10950 10694 11002
rect 10746 10950 10798 11002
rect 19862 10950 19914 11002
rect 19966 10950 20018 11002
rect 20070 10950 20122 11002
rect 29186 10950 29238 11002
rect 29290 10950 29342 11002
rect 29394 10950 29446 11002
rect 38510 10950 38562 11002
rect 38614 10950 38666 11002
rect 38718 10950 38770 11002
rect 6526 10782 6578 10834
rect 12238 10782 12290 10834
rect 15822 10782 15874 10834
rect 17558 10782 17610 10834
rect 18902 10782 18954 10834
rect 21030 10782 21082 10834
rect 37270 10782 37322 10834
rect 9550 10670 9602 10722
rect 29542 10670 29594 10722
rect 30848 10670 30900 10722
rect 36654 10670 36706 10722
rect 7982 10558 8034 10610
rect 8430 10558 8482 10610
rect 8654 10558 8706 10610
rect 9718 10502 9770 10554
rect 10222 10558 10274 10610
rect 11230 10585 11282 10637
rect 14254 10558 14306 10610
rect 14366 10558 14418 10610
rect 19294 10558 19346 10610
rect 19630 10558 19682 10610
rect 19742 10558 19794 10610
rect 23886 10558 23938 10610
rect 25118 10558 25170 10610
rect 25902 10558 25954 10610
rect 28702 10558 28754 10610
rect 29150 10558 29202 10610
rect 29262 10558 29314 10610
rect 29934 10558 29986 10610
rect 30102 10502 30154 10554
rect 30606 10558 30658 10610
rect 33966 10558 34018 10610
rect 27806 10446 27858 10498
rect 34750 10446 34802 10498
rect 8934 10334 8986 10386
rect 10464 10334 10516 10386
rect 13918 10334 13970 10386
rect 20078 10334 20130 10386
rect 23550 10334 23602 10386
rect 28366 10334 28418 10386
rect 5876 10166 5928 10218
rect 5980 10166 6032 10218
rect 6084 10166 6136 10218
rect 15200 10166 15252 10218
rect 15304 10166 15356 10218
rect 15408 10166 15460 10218
rect 24524 10166 24576 10218
rect 24628 10166 24680 10218
rect 24732 10166 24784 10218
rect 33848 10166 33900 10218
rect 33952 10166 34004 10218
rect 34056 10166 34108 10218
rect 34862 9998 34914 10050
rect 10166 9886 10218 9938
rect 12966 9886 13018 9938
rect 14422 9886 14474 9938
rect 14870 9886 14922 9938
rect 20470 9886 20522 9938
rect 23214 9886 23266 9938
rect 5518 9774 5570 9826
rect 6302 9774 6354 9826
rect 8990 9774 9042 9826
rect 9662 9774 9714 9826
rect 8206 9662 8258 9714
rect 9494 9718 9546 9770
rect 10446 9774 10498 9826
rect 13806 9774 13858 9826
rect 13918 9774 13970 9826
rect 15486 9746 15538 9798
rect 17502 9774 17554 9826
rect 20078 9774 20130 9826
rect 22430 9774 22482 9826
rect 25118 9774 25170 9826
rect 26126 9774 26178 9826
rect 26630 9830 26682 9882
rect 29262 9886 29314 9938
rect 31166 9886 31218 9938
rect 27302 9830 27354 9882
rect 27806 9774 27858 9826
rect 31950 9774 32002 9826
rect 32622 9774 32674 9826
rect 32846 9774 32898 9826
rect 33126 9774 33178 9826
rect 33406 9774 33458 9826
rect 37662 9774 37714 9826
rect 8748 9662 8800 9714
rect 13526 9662 13578 9714
rect 25884 9662 25936 9714
rect 26798 9662 26850 9714
rect 27134 9662 27186 9714
rect 37158 9718 37210 9770
rect 37904 9774 37956 9826
rect 28048 9662 28100 9714
rect 11566 9550 11618 9602
rect 18958 9550 19010 9602
rect 37326 9606 37378 9658
rect 32342 9550 32394 9602
rect 10538 9382 10590 9434
rect 10642 9382 10694 9434
rect 10746 9382 10798 9434
rect 19862 9382 19914 9434
rect 19966 9382 20018 9434
rect 20070 9382 20122 9434
rect 29186 9382 29238 9434
rect 29290 9382 29342 9434
rect 29394 9382 29446 9434
rect 38510 9382 38562 9434
rect 38614 9382 38666 9434
rect 38718 9382 38770 9434
rect 5966 9214 6018 9266
rect 17558 9214 17610 9266
rect 18230 9214 18282 9266
rect 35254 9214 35306 9266
rect 26574 9158 26626 9210
rect 8934 9102 8986 9154
rect 9774 9102 9826 9154
rect 27302 9102 27354 9154
rect 29038 9102 29090 9154
rect 29468 9102 29520 9154
rect 30382 9102 30434 9154
rect 7086 8990 7138 9042
rect 7814 8990 7866 9042
rect 8094 8990 8146 9042
rect 8318 8990 8370 9042
rect 8430 8990 8482 9042
rect 8654 8990 8706 9042
rect 11678 8990 11730 9042
rect 12462 8990 12514 9042
rect 12798 8990 12850 9042
rect 16942 8990 16994 9042
rect 20638 8990 20690 9042
rect 26238 8990 26290 9042
rect 26742 8934 26794 8986
rect 27582 8990 27634 9042
rect 27806 8990 27858 9042
rect 28124 8990 28176 9042
rect 28366 8990 28418 9042
rect 28870 8934 28922 8986
rect 29710 8990 29762 9042
rect 30214 8990 30266 9042
rect 30718 8990 30770 9042
rect 38334 8990 38386 9042
rect 35646 8878 35698 8930
rect 37550 8878 37602 8930
rect 14254 8766 14306 8818
rect 15822 8766 15874 8818
rect 19182 8766 19234 8818
rect 25996 8766 26048 8818
rect 32174 8766 32226 8818
rect 5876 8598 5928 8650
rect 5980 8598 6032 8650
rect 6084 8598 6136 8650
rect 15200 8598 15252 8650
rect 15304 8598 15356 8650
rect 15408 8598 15460 8650
rect 24524 8598 24576 8650
rect 24628 8598 24680 8650
rect 24732 8598 24784 8650
rect 33848 8598 33900 8650
rect 33952 8598 34004 8650
rect 34056 8598 34108 8650
rect 11510 8430 11562 8482
rect 13564 8430 13616 8482
rect 8560 8318 8612 8370
rect 7646 8206 7698 8258
rect 8318 8206 8370 8258
rect 7814 8150 7866 8202
rect 9326 8206 9378 8258
rect 9438 8206 9490 8258
rect 11790 8206 11842 8258
rect 12014 8206 12066 8258
rect 13806 8206 13858 8258
rect 14310 8262 14362 8314
rect 14982 8318 15034 8370
rect 18734 8318 18786 8370
rect 26070 8318 26122 8370
rect 36000 8318 36052 8370
rect 37904 8318 37956 8370
rect 17950 8206 18002 8258
rect 22206 8206 22258 8258
rect 23326 8206 23378 8258
rect 23550 8206 23602 8258
rect 26350 8206 26402 8258
rect 26462 8206 26514 8258
rect 27134 8206 27186 8258
rect 27246 8206 27298 8258
rect 29038 8206 29090 8258
rect 32062 8206 32114 8258
rect 32174 8206 32226 8258
rect 34190 8206 34242 8258
rect 34414 8206 34466 8258
rect 35758 8206 35810 8258
rect 9046 8094 9098 8146
rect 14478 8094 14530 8146
rect 35254 8150 35306 8202
rect 37662 8206 37714 8258
rect 20638 8094 20690 8146
rect 23046 8094 23098 8146
rect 26854 8094 26906 8146
rect 34694 8094 34746 8146
rect 35086 8094 35138 8146
rect 37158 8150 37210 8202
rect 36990 8094 37042 8146
rect 9942 7982 9994 8034
rect 17110 7982 17162 8034
rect 17782 7982 17834 8034
rect 22542 7982 22594 8034
rect 29374 7982 29426 8034
rect 30606 7982 30658 8034
rect 32510 7982 32562 8034
rect 10538 7814 10590 7866
rect 10642 7814 10694 7866
rect 10746 7814 10798 7866
rect 19862 7814 19914 7866
rect 19966 7814 20018 7866
rect 20070 7814 20122 7866
rect 29186 7814 29238 7866
rect 29290 7814 29342 7866
rect 29394 7814 29446 7866
rect 38510 7814 38562 7866
rect 38614 7814 38666 7866
rect 38718 7814 38770 7866
rect 11062 7646 11114 7698
rect 36654 7646 36706 7698
rect 7590 7534 7642 7586
rect 7982 7534 8034 7586
rect 12462 7534 12514 7586
rect 25436 7534 25488 7586
rect 27022 7590 27074 7642
rect 37998 7646 38050 7698
rect 26350 7534 26402 7586
rect 7086 7422 7138 7474
rect 7310 7422 7362 7474
rect 8150 7422 8202 7474
rect 8654 7422 8706 7474
rect 9438 7422 9490 7474
rect 9662 7422 9714 7474
rect 9942 7422 9994 7474
rect 11902 7422 11954 7474
rect 12126 7422 12178 7474
rect 14366 7422 14418 7474
rect 15150 7422 15202 7474
rect 16718 7422 16770 7474
rect 16942 7422 16994 7474
rect 17278 7422 17330 7474
rect 20750 7422 20802 7474
rect 21254 7366 21306 7418
rect 21422 7422 21474 7474
rect 21870 7422 21922 7474
rect 24558 7422 24610 7474
rect 26182 7478 26234 7530
rect 29038 7534 29090 7586
rect 35216 7534 35268 7586
rect 25678 7422 25730 7474
rect 15542 7310 15594 7362
rect 18062 7310 18114 7362
rect 19966 7310 20018 7362
rect 26854 7366 26906 7418
rect 27358 7422 27410 7474
rect 28366 7422 28418 7474
rect 22654 7310 22706 7362
rect 28870 7366 28922 7418
rect 30942 7422 30994 7474
rect 34302 7422 34354 7474
rect 34470 7366 34522 7418
rect 34974 7422 35026 7474
rect 35534 7422 35586 7474
rect 38334 7422 38386 7474
rect 8896 7198 8948 7250
rect 11622 7198 11674 7250
rect 16438 7198 16490 7250
rect 20508 7198 20560 7250
rect 27600 7198 27652 7250
rect 28124 7198 28176 7250
rect 30606 7198 30658 7250
rect 5876 7030 5928 7082
rect 5980 7030 6032 7082
rect 6084 7030 6136 7082
rect 15200 7030 15252 7082
rect 15304 7030 15356 7082
rect 15408 7030 15460 7082
rect 24524 7030 24576 7082
rect 24628 7030 24680 7082
rect 24732 7030 24784 7082
rect 33848 7030 33900 7082
rect 33952 7030 34004 7082
rect 34056 7030 34108 7082
rect 15356 6862 15408 6914
rect 17950 6862 18002 6914
rect 22542 6862 22594 6914
rect 8094 6638 8146 6690
rect 10110 6638 10162 6690
rect 10390 6638 10442 6690
rect 10670 6638 10722 6690
rect 10782 6638 10834 6690
rect 11118 6638 11170 6690
rect 13806 6638 13858 6690
rect 15598 6638 15650 6690
rect 14310 6582 14362 6634
rect 16270 6638 16322 6690
rect 13564 6526 13616 6578
rect 16102 6582 16154 6634
rect 16494 6638 16546 6690
rect 18846 6638 18898 6690
rect 19014 6694 19066 6746
rect 19518 6638 19570 6690
rect 19760 6638 19812 6690
rect 20078 6638 20130 6690
rect 20302 6638 20354 6690
rect 20582 6638 20634 6690
rect 21758 6638 21810 6690
rect 23998 6638 24050 6690
rect 24670 6638 24722 6690
rect 26686 6638 26738 6690
rect 29486 6638 29538 6690
rect 29654 6638 29706 6690
rect 30158 6638 30210 6690
rect 30718 6638 30770 6690
rect 30942 6638 30994 6690
rect 33294 6638 33346 6690
rect 33966 6638 34018 6690
rect 14478 6526 14530 6578
rect 33462 6582 33514 6634
rect 34638 6638 34690 6690
rect 36990 6638 37042 6690
rect 37662 6638 37714 6690
rect 37158 6582 37210 6634
rect 30400 6526 30452 6578
rect 31222 6526 31274 6578
rect 34208 6526 34260 6578
rect 37904 6526 37956 6578
rect 6638 6414 6690 6466
rect 8990 6414 9042 6466
rect 12238 6414 12290 6466
rect 21422 6414 21474 6466
rect 25790 6414 25842 6466
rect 27806 6414 27858 6466
rect 36094 6414 36146 6466
rect 10538 6246 10590 6298
rect 10642 6246 10694 6298
rect 10746 6246 10798 6298
rect 19862 6246 19914 6298
rect 19966 6246 20018 6298
rect 20070 6246 20122 6298
rect 29186 6246 29238 6298
rect 29290 6246 29342 6298
rect 29394 6246 29446 6298
rect 38510 6246 38562 6298
rect 38614 6246 38666 6298
rect 38718 6246 38770 6298
rect 9998 6022 10050 6074
rect 8542 5966 8594 6018
rect 10688 5966 10740 6018
rect 13694 5966 13746 6018
rect 30046 6022 30098 6074
rect 21422 5966 21474 6018
rect 24614 5966 24666 6018
rect 29468 5966 29520 6018
rect 5854 5854 5906 5906
rect 6638 5854 6690 5906
rect 9942 5854 9994 5906
rect 10446 5854 10498 5906
rect 11006 5854 11058 5906
rect 11790 5854 11842 5906
rect 14142 5881 14194 5933
rect 17502 5881 17554 5933
rect 20302 5854 20354 5906
rect 20414 5854 20466 5906
rect 21590 5854 21642 5906
rect 22094 5854 22146 5906
rect 22766 5854 22818 5906
rect 22878 5854 22930 5906
rect 24110 5854 24162 5906
rect 24334 5854 24386 5906
rect 25230 5881 25282 5933
rect 28124 5854 28176 5906
rect 28870 5910 28922 5962
rect 30718 5966 30770 6018
rect 28366 5854 28418 5906
rect 29038 5854 29090 5906
rect 30214 5910 30266 5962
rect 31632 5966 31684 6018
rect 30886 5910 30938 5962
rect 33164 5966 33216 6018
rect 35142 5966 35194 6018
rect 38110 5966 38162 6018
rect 29710 5854 29762 5906
rect 31390 5854 31442 5906
rect 31950 5854 32002 5906
rect 32174 5854 32226 5906
rect 33910 5910 33962 5962
rect 33406 5854 33458 5906
rect 34078 5854 34130 5906
rect 34638 5854 34690 5906
rect 34862 5854 34914 5906
rect 35422 5854 35474 5906
rect 36206 5854 36258 5906
rect 20974 5742 21026 5794
rect 21198 5742 21250 5794
rect 15150 5630 15202 5682
rect 18510 5630 18562 5682
rect 20694 5630 20746 5682
rect 22336 5630 22388 5682
rect 23158 5630 23210 5682
rect 26238 5630 26290 5682
rect 32454 5630 32506 5682
rect 5876 5462 5928 5514
rect 5980 5462 6032 5514
rect 6084 5462 6136 5514
rect 15200 5462 15252 5514
rect 15304 5462 15356 5514
rect 15408 5462 15460 5514
rect 24524 5462 24576 5514
rect 24628 5462 24680 5514
rect 24732 5462 24784 5514
rect 33848 5462 33900 5514
rect 33952 5462 34004 5514
rect 34056 5462 34108 5514
rect 37998 5294 38050 5346
rect 8318 5182 8370 5234
rect 10222 5182 10274 5234
rect 14254 5182 14306 5234
rect 16270 5182 16322 5234
rect 18174 5182 18226 5234
rect 25566 5182 25618 5234
rect 27470 5182 27522 5234
rect 32622 5182 32674 5234
rect 35646 5182 35698 5234
rect 36262 5182 36314 5234
rect 37158 5182 37210 5234
rect 1934 5070 1986 5122
rect 4174 5042 4226 5094
rect 6638 5070 6690 5122
rect 7310 5070 7362 5122
rect 7982 5070 8034 5122
rect 11006 5070 11058 5122
rect 13022 5070 13074 5122
rect 15374 5070 15426 5122
rect 15486 5070 15538 5122
rect 20862 5070 20914 5122
rect 23662 5070 23714 5122
rect 24782 5070 24834 5122
rect 29934 5070 29986 5122
rect 30718 5070 30770 5122
rect 32958 5070 33010 5122
rect 33742 5070 33794 5122
rect 38334 5070 38386 5122
rect 6302 4846 6354 4898
rect 6974 4846 7026 4898
rect 7646 4846 7698 4898
rect 11902 4846 11954 4898
rect 18790 4846 18842 4898
rect 19406 4846 19458 4898
rect 22542 4846 22594 4898
rect 37606 4846 37658 4898
rect 10538 4678 10590 4730
rect 10642 4678 10694 4730
rect 10746 4678 10798 4730
rect 19862 4678 19914 4730
rect 19966 4678 20018 4730
rect 20070 4678 20122 4730
rect 29186 4678 29238 4730
rect 29290 4678 29342 4730
rect 29394 4678 29446 4730
rect 38510 4678 38562 4730
rect 38614 4678 38666 4730
rect 38718 4678 38770 4730
rect 2774 4510 2826 4562
rect 30718 4510 30770 4562
rect 34078 4510 34130 4562
rect 38278 4510 38330 4562
rect 15822 4398 15874 4450
rect 17446 4398 17498 4450
rect 21758 4398 21810 4450
rect 26518 4398 26570 4450
rect 29598 4398 29650 4450
rect 35086 4398 35138 4450
rect 36000 4398 36052 4450
rect 3502 4286 3554 4338
rect 5854 4313 5906 4365
rect 6526 4313 6578 4365
rect 10110 4313 10162 4365
rect 12574 4286 12626 4338
rect 13358 4286 13410 4338
rect 15262 4286 15314 4338
rect 15990 4286 16042 4338
rect 16494 4286 16546 4338
rect 16736 4286 16788 4338
rect 17726 4286 17778 4338
rect 17950 4286 18002 4338
rect 18342 4286 18394 4338
rect 18510 4286 18562 4338
rect 19294 4286 19346 4338
rect 23662 4286 23714 4338
rect 24446 4286 24498 4338
rect 26014 4286 26066 4338
rect 26238 4286 26290 4338
rect 26910 4286 26962 4338
rect 27694 4286 27746 4338
rect 31838 4286 31890 4338
rect 35254 4342 35306 4394
rect 32958 4286 33010 4338
rect 35758 4286 35810 4338
rect 21198 4174 21250 4226
rect 37830 4174 37882 4226
rect 3166 4062 3218 4114
rect 4846 4062 4898 4114
rect 7534 4062 7586 4114
rect 10894 4062 10946 4114
rect 5876 3894 5928 3946
rect 5980 3894 6032 3946
rect 6084 3894 6136 3946
rect 15200 3894 15252 3946
rect 15304 3894 15356 3946
rect 15408 3894 15460 3946
rect 24524 3894 24576 3946
rect 24628 3894 24680 3946
rect 24732 3894 24784 3946
rect 33848 3894 33900 3946
rect 33952 3894 34004 3946
rect 34056 3894 34108 3946
rect 5742 3726 5794 3778
rect 9550 3726 9602 3778
rect 13190 3726 13242 3778
rect 27470 3726 27522 3778
rect 28478 3726 28530 3778
rect 30158 3726 30210 3778
rect 32398 3726 32450 3778
rect 33854 3726 33906 3778
rect 36206 3726 36258 3778
rect 37438 3726 37490 3778
rect 3502 3614 3554 3666
rect 22094 3614 22146 3666
rect 25566 3614 25618 3666
rect 2830 3474 2882 3526
rect 6078 3502 6130 3554
rect 6638 3474 6690 3526
rect 8318 3502 8370 3554
rect 9886 3502 9938 3554
rect 10222 3474 10274 3526
rect 13470 3502 13522 3554
rect 13582 3502 13634 3554
rect 13918 3474 13970 3526
rect 18062 3474 18114 3526
rect 21086 3474 21138 3526
rect 24558 3474 24610 3526
rect 27806 3502 27858 3554
rect 28814 3502 28866 3554
rect 29654 3502 29706 3554
rect 30494 3502 30546 3554
rect 30886 3502 30938 3554
rect 31670 3502 31722 3554
rect 32062 3502 32114 3554
rect 33518 3502 33570 3554
rect 35870 3502 35922 3554
rect 37102 3502 37154 3554
rect 37998 3502 38050 3554
rect 38334 3502 38386 3554
rect 29206 3390 29258 3442
rect 33350 3390 33402 3442
rect 35478 3390 35530 3442
rect 36934 3390 36986 3442
rect 11790 3278 11842 3330
rect 15598 3278 15650 3330
rect 19070 3278 19122 3330
rect 10538 3110 10590 3162
rect 10642 3110 10694 3162
rect 10746 3110 10798 3162
rect 19862 3110 19914 3162
rect 19966 3110 20018 3162
rect 20070 3110 20122 3162
rect 29186 3110 29238 3162
rect 29290 3110 29342 3162
rect 29394 3110 29446 3162
rect 38510 3110 38562 3162
rect 38614 3110 38666 3162
rect 38718 3110 38770 3162
<< metal2 >>
rect 3136 39200 3248 40000
rect 4256 39200 4368 40000
rect 5376 39200 5488 40000
rect 6496 39200 6608 40000
rect 7616 39200 7728 40000
rect 8736 39200 8848 40000
rect 9856 39200 9968 40000
rect 10976 39200 11088 40000
rect 12096 39200 12208 40000
rect 13216 39200 13328 40000
rect 14336 39200 14448 40000
rect 15456 39200 15568 40000
rect 16576 39200 16688 40000
rect 17696 39200 17808 40000
rect 17948 39228 18340 39284
rect 3164 36820 3220 39200
rect 4284 37380 4340 39200
rect 5404 37716 5460 39200
rect 5404 37660 5684 37716
rect 4284 37324 4564 37380
rect 4508 36932 4564 37324
rect 5628 36932 5684 37660
rect 6524 36932 6580 39200
rect 7644 37828 7700 39200
rect 7644 37772 7924 37828
rect 7868 36932 7924 37772
rect 8764 36932 8820 39200
rect 4508 36876 4620 36932
rect 5628 36876 5740 36932
rect 3164 36764 3500 36820
rect 3444 36314 3500 36764
rect 3444 36262 3446 36314
rect 3498 36262 3500 36314
rect 3444 36250 3500 36262
rect 4564 36314 4620 36876
rect 4564 36262 4566 36314
rect 4618 36262 4620 36314
rect 4564 36250 4620 36262
rect 5684 36314 5740 36876
rect 5874 36876 6138 36886
rect 6524 36876 6860 36932
rect 7868 36876 7980 36932
rect 5930 36820 5978 36876
rect 6034 36820 6082 36876
rect 5874 36810 6138 36820
rect 5684 36262 5686 36314
rect 5738 36262 5740 36314
rect 5684 36250 5740 36262
rect 6804 36314 6860 36876
rect 6804 36262 6806 36314
rect 6858 36262 6860 36314
rect 6804 36250 6860 36262
rect 7924 36314 7980 36876
rect 7924 36262 7926 36314
rect 7978 36262 7980 36314
rect 7924 36250 7980 36262
rect 8708 36876 8820 36932
rect 8708 36314 8764 36876
rect 9884 36484 9940 39200
rect 11004 37604 11060 39200
rect 11004 37548 11284 37604
rect 8708 36262 8710 36314
rect 8762 36262 8764 36314
rect 9716 36428 9940 36484
rect 10220 36454 10276 36466
rect 9716 36314 9772 36428
rect 8708 36250 8764 36262
rect 8876 36260 8932 36270
rect 9716 36262 9718 36314
rect 9770 36262 9772 36314
rect 9716 36250 9772 36262
rect 10220 36402 10222 36454
rect 10274 36402 10276 36454
rect 8876 35810 8932 36204
rect 8876 35758 8878 35810
rect 8930 35758 8932 35810
rect 2492 35698 2548 35710
rect 2492 35646 2494 35698
rect 2546 35646 2548 35698
rect 2380 32564 2436 32574
rect 2492 32564 2548 35646
rect 5516 35700 5572 35710
rect 3276 35588 3332 35598
rect 2940 35586 3332 35588
rect 2940 35534 3278 35586
rect 3330 35534 3332 35586
rect 2940 35532 3332 35534
rect 2940 35138 2996 35532
rect 3276 35522 3332 35532
rect 5180 35586 5236 35598
rect 5180 35534 5182 35586
rect 5234 35534 5236 35586
rect 5180 35476 5236 35534
rect 5180 35410 5236 35420
rect 2940 35086 2942 35138
rect 2994 35086 2996 35138
rect 2940 35074 2996 35086
rect 4060 34916 4116 34926
rect 4060 34914 4340 34916
rect 4060 34862 4062 34914
rect 4114 34862 4340 34914
rect 4060 34860 4340 34862
rect 4060 34850 4116 34860
rect 2380 32562 2660 32564
rect 2380 32510 2382 32562
rect 2434 32510 2660 32562
rect 2380 32508 2660 32510
rect 2380 32498 2436 32508
rect 2492 31892 2548 31902
rect 1988 31108 2044 31118
rect 1988 31050 2044 31052
rect 1820 30996 1876 31006
rect 1708 30994 1876 30996
rect 1708 30942 1822 30994
rect 1874 30942 1876 30994
rect 1708 30940 1876 30942
rect 1708 30098 1764 30940
rect 1820 30930 1876 30940
rect 1988 30998 1990 31050
rect 2042 30998 2044 31050
rect 1988 30436 2044 30998
rect 2492 30994 2548 31836
rect 2492 30942 2494 30994
rect 2546 30942 2548 30994
rect 2492 30930 2548 30942
rect 2604 30548 2660 32508
rect 3164 32450 3220 32462
rect 3164 32398 3166 32450
rect 3218 32398 3220 32450
rect 3164 32002 3220 32398
rect 3164 31950 3166 32002
rect 3218 31950 3220 32002
rect 3164 31938 3220 31950
rect 4284 32004 4340 34860
rect 5516 34914 5572 35644
rect 5796 35700 5852 35710
rect 5796 35606 5852 35644
rect 6188 35700 6244 35710
rect 6188 35606 6244 35644
rect 6972 35588 7028 35598
rect 6972 35494 7028 35532
rect 8764 35588 8820 35598
rect 7532 35364 7588 35374
rect 5874 35308 6138 35318
rect 5930 35252 5978 35308
rect 6034 35252 6082 35308
rect 5874 35242 6138 35252
rect 6300 34916 6356 34926
rect 5516 34862 5518 34914
rect 5570 34862 5572 34914
rect 5516 32788 5572 34862
rect 5964 34914 6356 34916
rect 5964 34862 6302 34914
rect 6354 34862 6356 34914
rect 5964 34860 6356 34862
rect 5964 34354 6020 34860
rect 6300 34850 6356 34860
rect 5964 34302 5966 34354
rect 6018 34302 6020 34354
rect 5964 34290 6020 34302
rect 7084 34132 7140 34142
rect 7084 34130 7476 34132
rect 7084 34078 7086 34130
rect 7138 34078 7476 34130
rect 7084 34076 7476 34078
rect 7084 34066 7140 34076
rect 7420 33906 7476 34076
rect 7420 33854 7422 33906
rect 7474 33854 7476 33906
rect 7420 33842 7476 33854
rect 5874 33740 6138 33750
rect 5930 33684 5978 33740
rect 6034 33684 6082 33740
rect 5874 33674 6138 33684
rect 7532 33236 7588 35308
rect 8764 35138 8820 35532
rect 8764 35086 8766 35138
rect 8818 35086 8820 35138
rect 8764 35074 8820 35086
rect 8204 34804 8260 34814
rect 8876 34804 8932 35758
rect 9548 35700 9604 35710
rect 9548 35588 9604 35644
rect 9716 35588 9772 35598
rect 9492 35586 9772 35588
rect 9492 35534 9718 35586
rect 9770 35534 9772 35586
rect 9492 35532 9772 35534
rect 9492 35026 9548 35532
rect 9716 35522 9772 35532
rect 10108 35252 10164 35262
rect 9492 34974 9494 35026
rect 9546 34974 9548 35026
rect 9492 34962 9548 34974
rect 9940 35028 9996 35038
rect 10108 35028 10164 35196
rect 9940 35026 10164 35028
rect 9940 34974 9942 35026
rect 9994 34974 10164 35026
rect 9940 34972 10164 34974
rect 9940 34962 9996 34972
rect 8204 34710 8260 34748
rect 8764 34748 8932 34804
rect 9100 34914 9156 34926
rect 9100 34862 9102 34914
rect 9154 34862 9156 34914
rect 8596 34132 8652 34142
rect 8596 34038 8652 34076
rect 7756 33908 7812 33918
rect 7756 33906 7924 33908
rect 7756 33854 7758 33906
rect 7810 33854 7924 33906
rect 7756 33852 7924 33854
rect 7756 33842 7812 33852
rect 5684 32788 5740 32798
rect 5516 32786 5740 32788
rect 5516 32734 5686 32786
rect 5738 32734 5740 32786
rect 5516 32732 5740 32734
rect 5628 32722 5740 32732
rect 5068 32452 5124 32462
rect 5068 32450 5236 32452
rect 5068 32398 5070 32450
rect 5122 32398 5236 32450
rect 5068 32396 5236 32398
rect 5068 32386 5124 32396
rect 4284 31938 4340 31948
rect 5180 31892 5236 32396
rect 5180 31826 5236 31836
rect 5404 31892 5460 31902
rect 4284 31778 4340 31790
rect 4284 31726 4286 31778
rect 4338 31726 4340 31778
rect 4284 31444 4340 31726
rect 4284 31378 4340 31388
rect 4396 31778 4452 31790
rect 4396 31726 4398 31778
rect 4450 31726 4452 31778
rect 4396 31220 4452 31726
rect 4620 31780 4676 31790
rect 4620 31686 4676 31724
rect 5068 31780 5124 31790
rect 4900 31668 4956 31678
rect 4900 31666 5012 31668
rect 4900 31614 4902 31666
rect 4954 31614 5012 31666
rect 4900 31602 5012 31614
rect 4060 31164 4452 31220
rect 3052 30996 3108 31006
rect 2734 30884 2790 30894
rect 2734 30790 2790 30828
rect 3052 30660 3108 30940
rect 2828 30604 3108 30660
rect 3836 30882 3892 30894
rect 3836 30830 3838 30882
rect 3890 30830 3892 30882
rect 2828 30548 2884 30604
rect 2268 30492 2884 30548
rect 1988 30380 2100 30436
rect 2044 30324 2100 30380
rect 2044 30258 2100 30268
rect 1876 30212 1932 30222
rect 1876 30118 1932 30156
rect 1708 30046 1710 30098
rect 1762 30046 1764 30098
rect 1708 26292 1764 30046
rect 1708 26226 1764 26236
rect 2268 28642 2324 30492
rect 3724 30436 3780 30446
rect 3836 30436 3892 30830
rect 3724 30434 3892 30436
rect 3724 30382 3726 30434
rect 3778 30382 3892 30434
rect 3724 30380 3892 30382
rect 3724 30370 3780 30380
rect 2380 30324 2436 30334
rect 2380 30210 2436 30268
rect 2380 30158 2382 30210
rect 2434 30158 2436 30210
rect 2380 30146 2436 30158
rect 2622 30324 2678 30334
rect 2622 30210 2678 30268
rect 4060 30324 4116 31164
rect 4060 30258 4116 30268
rect 2622 30158 2624 30210
rect 2676 30158 2678 30210
rect 2622 30146 2678 30158
rect 4844 30212 4900 30222
rect 4956 30212 5012 31602
rect 4844 30210 5012 30212
rect 4844 30158 4846 30210
rect 4898 30158 5012 30210
rect 4844 30156 5012 30158
rect 5068 31220 5124 31724
rect 4844 30146 4900 30156
rect 5068 30100 5124 31164
rect 4956 30044 5124 30100
rect 4956 29764 5012 30044
rect 4844 29708 5012 29764
rect 2492 29428 2548 29438
rect 2492 29426 2996 29428
rect 2492 29374 2494 29426
rect 2546 29374 2996 29426
rect 2492 29372 2996 29374
rect 2492 29362 2548 29372
rect 2268 28590 2270 28642
rect 2322 28590 2324 28642
rect 2044 25284 2100 25294
rect 2044 24722 2100 25228
rect 2268 25284 2324 28590
rect 2940 27982 2996 29372
rect 3052 29204 3108 29214
rect 3052 28754 3108 29148
rect 3612 29204 3668 29214
rect 4714 29204 4770 29214
rect 3612 29110 3668 29148
rect 4172 29202 4770 29204
rect 4172 29150 4716 29202
rect 4768 29150 4770 29202
rect 4172 29148 4770 29150
rect 3052 28702 3054 28754
rect 3106 28702 3108 28754
rect 3052 28690 3108 28702
rect 4172 28420 4228 29148
rect 4714 29138 4770 29148
rect 3500 28364 4228 28420
rect 2940 27970 3052 27982
rect 2940 27918 2998 27970
rect 3050 27918 3052 27970
rect 2940 27916 3052 27918
rect 2996 27906 3052 27916
rect 3276 27860 3332 27870
rect 3276 27766 3332 27804
rect 3500 27858 3556 28364
rect 3500 27806 3502 27858
rect 3554 27806 3556 27858
rect 3500 27794 3556 27806
rect 4396 27858 4452 27870
rect 4396 27806 4398 27858
rect 4450 27806 4452 27858
rect 3612 27636 3668 27646
rect 3108 26404 3164 26414
rect 3108 26346 3164 26348
rect 2940 26292 2996 26302
rect 3108 26294 3110 26346
rect 3162 26294 3164 26346
rect 3108 26282 3164 26294
rect 3612 26290 3668 27580
rect 4228 27636 4284 27646
rect 4228 27186 4284 27580
rect 4228 27134 4230 27186
rect 4282 27134 4284 27186
rect 4228 27122 4284 27134
rect 4396 26908 4452 27806
rect 4844 27860 4900 29708
rect 5404 29494 5460 31836
rect 5628 30996 5684 32722
rect 7196 32562 7252 32574
rect 7196 32510 7198 32562
rect 7250 32510 7252 32562
rect 7196 32452 7252 32510
rect 7196 32386 7252 32396
rect 7364 32564 7420 32574
rect 7364 32394 7420 32508
rect 7364 32342 7366 32394
rect 7418 32342 7420 32394
rect 7364 32330 7420 32342
rect 5874 32172 6138 32182
rect 5930 32116 5978 32172
rect 6034 32116 6082 32172
rect 5874 32106 6138 32116
rect 7252 31722 7308 31734
rect 7084 31668 7140 31678
rect 6860 31612 7084 31668
rect 6580 31444 6636 31454
rect 6300 31220 6356 31230
rect 5740 31108 5796 31118
rect 5740 31014 5796 31052
rect 5628 30436 5684 30940
rect 6076 30994 6132 31006
rect 6076 30942 6078 30994
rect 6130 30942 6132 30994
rect 6076 30884 6132 30942
rect 6300 30994 6356 31164
rect 6580 31106 6636 31388
rect 6580 31054 6582 31106
rect 6634 31054 6636 31106
rect 6580 31042 6636 31054
rect 6300 30942 6302 30994
rect 6354 30942 6356 30994
rect 6300 30930 6356 30942
rect 6076 30818 6132 30828
rect 5874 30604 6138 30614
rect 5930 30548 5978 30604
rect 6034 30548 6082 30604
rect 5874 30538 6138 30548
rect 5628 30380 6188 30436
rect 5404 29482 5516 29494
rect 4396 26852 4676 26908
rect 2940 26198 2996 26236
rect 3612 26238 3614 26290
rect 3666 26238 3668 26290
rect 2268 25218 2324 25228
rect 2828 25282 2884 25294
rect 2828 25230 2830 25282
rect 2882 25230 2884 25282
rect 2044 24670 2046 24722
rect 2098 24670 2100 24722
rect 2044 22148 2100 24670
rect 2828 24722 2884 25230
rect 3612 25060 3668 26238
rect 4060 26292 4116 26302
rect 3854 26068 3910 26078
rect 3612 24994 3668 25004
rect 3836 26066 3910 26068
rect 3836 26014 3856 26066
rect 3908 26014 3910 26066
rect 3836 26002 3910 26014
rect 3836 24948 3892 26002
rect 3836 24882 3892 24892
rect 3948 25506 4004 25518
rect 3948 25454 3950 25506
rect 4002 25454 4004 25506
rect 3948 24836 4004 25454
rect 3948 24770 4004 24780
rect 2828 24670 2830 24722
rect 2882 24670 2884 24722
rect 2828 24658 2884 24670
rect 3836 24164 3892 24174
rect 4060 24164 4116 26236
rect 4508 26290 4564 26302
rect 4508 26238 4510 26290
rect 4562 26238 4564 26290
rect 4340 25284 4396 25294
rect 4508 25284 4564 26238
rect 4620 25742 4676 26852
rect 4620 25730 4732 25742
rect 4620 25678 4678 25730
rect 4730 25678 4732 25730
rect 4620 25676 4732 25678
rect 4676 25666 4732 25676
rect 4844 25508 4900 27804
rect 4956 29428 5012 29438
rect 5404 29430 5462 29482
rect 5514 29430 5516 29482
rect 5404 29428 5516 29430
rect 5460 29418 5516 29428
rect 5628 29426 5684 29438
rect 4956 28754 5012 29372
rect 4956 28702 4958 28754
rect 5010 28702 5012 28754
rect 4956 26404 5012 28702
rect 5628 29374 5630 29426
rect 5682 29374 5684 29426
rect 5516 27636 5572 27646
rect 4956 26338 5012 26348
rect 5292 27634 5572 27636
rect 5292 27582 5518 27634
rect 5570 27582 5572 27634
rect 5292 27580 5572 27582
rect 5292 26290 5348 27580
rect 5516 27570 5572 27580
rect 5628 26908 5684 29374
rect 5740 28766 5796 30380
rect 6132 30210 6188 30380
rect 6132 30158 6134 30210
rect 6186 30158 6188 30210
rect 6132 30146 6188 30158
rect 6748 30212 6804 30222
rect 6580 29092 6636 29102
rect 5874 29036 6138 29046
rect 5930 28980 5978 29036
rect 6034 28980 6082 29036
rect 5874 28970 6138 28980
rect 5740 28754 5852 28766
rect 5740 28702 5798 28754
rect 5850 28702 5852 28754
rect 5740 28700 5852 28702
rect 5796 28690 5852 28700
rect 6580 28756 6636 29036
rect 6748 28868 6804 30156
rect 6860 30210 6916 31612
rect 7084 31574 7140 31612
rect 7252 31670 7254 31722
rect 7306 31670 7308 31722
rect 7252 31332 7308 31670
rect 7252 31276 7476 31332
rect 7420 31162 7476 31276
rect 7420 31110 7422 31162
rect 7474 31110 7476 31162
rect 7420 31098 7476 31110
rect 7308 31009 7364 31021
rect 7308 30996 7310 31009
rect 7362 30996 7364 31009
rect 7308 30917 7364 30940
rect 7532 30772 7588 33180
rect 7756 32788 7812 32798
rect 7756 32562 7812 32732
rect 7756 32510 7758 32562
rect 7810 32510 7812 32562
rect 7756 32498 7812 32510
rect 7644 32452 7700 32462
rect 7644 30994 7700 32396
rect 7756 31778 7812 31790
rect 7756 31726 7758 31778
rect 7810 31726 7812 31778
rect 7756 31108 7812 31726
rect 7756 31042 7812 31052
rect 7644 30942 7646 30994
rect 7698 30942 7700 30994
rect 7644 30930 7700 30942
rect 7532 30716 7700 30772
rect 6860 30158 6862 30210
rect 6914 30158 6916 30210
rect 7532 30212 7588 30222
rect 6860 29652 6916 30158
rect 7028 30154 7084 30166
rect 7028 30102 7030 30154
rect 7082 30102 7084 30154
rect 7532 30118 7588 30156
rect 7028 29764 7084 30102
rect 7644 30100 7700 30716
rect 7868 30324 7924 33852
rect 8764 33346 8820 34748
rect 8764 33294 8766 33346
rect 8818 33294 8820 33346
rect 8764 33282 8820 33294
rect 8876 34130 8932 34142
rect 8876 34078 8878 34130
rect 8930 34078 8932 34130
rect 8428 33122 8484 33134
rect 8428 33070 8430 33122
rect 8482 33070 8484 33122
rect 8428 32788 8484 33070
rect 8428 32722 8484 32732
rect 8764 33124 8820 33134
rect 8092 32577 8148 32589
rect 8092 32525 8094 32577
rect 8146 32525 8148 32577
rect 8092 32340 8148 32525
rect 8428 32564 8484 32574
rect 8428 32470 8484 32508
rect 8652 32564 8708 32574
rect 8764 32564 8820 33068
rect 8652 32562 8820 32564
rect 8652 32510 8654 32562
rect 8706 32510 8820 32562
rect 8652 32508 8820 32510
rect 8876 32564 8932 34078
rect 8988 34130 9044 34142
rect 8988 34078 8990 34130
rect 9042 34078 9044 34130
rect 8988 33796 9044 34078
rect 8988 33730 9044 33740
rect 9100 33582 9156 34862
rect 10108 34914 10164 34972
rect 10108 34862 10110 34914
rect 10162 34862 10164 34914
rect 10108 34850 10164 34862
rect 10220 34804 10276 36402
rect 10536 36092 10800 36102
rect 10592 36036 10640 36092
rect 10696 36036 10744 36092
rect 10536 36026 10800 36036
rect 11228 35934 11284 37548
rect 12124 37380 12180 39200
rect 12124 37324 12628 37380
rect 12348 36484 12404 36494
rect 12348 36390 12404 36428
rect 11228 35922 11340 35934
rect 11228 35870 11286 35922
rect 11338 35870 11340 35922
rect 11228 35868 11340 35870
rect 11284 35858 11340 35868
rect 12236 35698 12292 35710
rect 12236 35646 12238 35698
rect 12290 35646 12292 35698
rect 10948 35586 11004 35598
rect 10948 35534 10950 35586
rect 11002 35534 11004 35586
rect 10948 35252 11004 35534
rect 11900 35476 11956 35486
rect 12236 35476 12292 35646
rect 11900 35474 12068 35476
rect 11900 35422 11902 35474
rect 11954 35422 12068 35474
rect 11900 35420 12068 35422
rect 11900 35410 11956 35420
rect 10948 35186 11004 35196
rect 9436 34132 9492 34142
rect 9436 34038 9492 34076
rect 9044 33570 9156 33582
rect 9044 33518 9046 33570
rect 9098 33518 9156 33570
rect 9044 33516 9156 33518
rect 9436 33796 9492 33806
rect 9044 33506 9100 33516
rect 9436 33460 9492 33740
rect 9324 33346 9380 33358
rect 9324 33294 9326 33346
rect 9378 33294 9380 33346
rect 9324 32788 9380 33294
rect 9436 33346 9492 33404
rect 9436 33294 9438 33346
rect 9490 33294 9492 33346
rect 9436 33282 9492 33294
rect 10052 33348 10108 33358
rect 10052 33254 10108 33292
rect 9324 32732 9660 32788
rect 9604 32674 9660 32732
rect 9604 32622 9606 32674
rect 9658 32622 9660 32674
rect 9604 32610 9660 32622
rect 9884 32676 9940 32686
rect 9884 32618 9940 32620
rect 9884 32566 9886 32618
rect 9938 32566 9940 32618
rect 10108 32590 10164 32602
rect 8876 32508 9492 32564
rect 9884 32554 9940 32566
rect 9996 32564 10052 32574
rect 8652 32498 8708 32508
rect 8204 32452 8260 32462
rect 8204 32450 8372 32452
rect 8204 32398 8206 32450
rect 8258 32398 8372 32450
rect 8204 32396 8372 32398
rect 8204 32386 8260 32396
rect 8092 32274 8148 32284
rect 8204 32004 8260 32014
rect 7998 31780 8054 31790
rect 7998 31686 8054 31724
rect 8204 31556 8260 31948
rect 8316 31892 8372 32396
rect 8316 31836 8652 31892
rect 8596 31834 8652 31836
rect 8596 31782 8598 31834
rect 8650 31782 8652 31834
rect 8596 31770 8652 31782
rect 8428 31668 8484 31678
rect 8428 31574 8484 31612
rect 8036 31500 8260 31556
rect 8036 31106 8092 31500
rect 8036 31054 8038 31106
rect 8090 31054 8092 31106
rect 8036 31042 8092 31054
rect 8316 30996 8372 31006
rect 8260 30994 8372 30996
rect 8260 30942 8318 30994
rect 8370 30942 8372 30994
rect 8260 30930 8372 30942
rect 8540 30996 8596 31006
rect 8764 30996 8820 32508
rect 9436 32452 9492 32508
rect 9436 32396 9884 32452
rect 8932 32340 8988 32350
rect 8932 32246 8988 32284
rect 9342 32228 9398 32238
rect 9100 31892 9156 31902
rect 9100 31778 9156 31836
rect 9342 31890 9398 32172
rect 9342 31838 9344 31890
rect 9396 31838 9398 31890
rect 9342 31826 9398 31838
rect 9828 31890 9884 32396
rect 9828 31838 9830 31890
rect 9882 31838 9884 31890
rect 9828 31826 9884 31838
rect 9996 31892 10052 32508
rect 10108 32538 10110 32590
rect 10162 32538 10164 32590
rect 10108 32116 10164 32538
rect 10108 32050 10164 32060
rect 9996 31836 10164 31892
rect 9100 31726 9102 31778
rect 9154 31726 9156 31778
rect 9100 31714 9156 31726
rect 10108 31750 10164 31836
rect 10108 31698 10110 31750
rect 10162 31698 10164 31750
rect 10108 31686 10164 31698
rect 10052 31556 10108 31566
rect 8540 30994 8708 30996
rect 8540 30942 8542 30994
rect 8594 30942 8708 30994
rect 8540 30940 8708 30942
rect 8540 30930 8596 30940
rect 8260 30434 8316 30930
rect 8260 30382 8262 30434
rect 8314 30382 8316 30434
rect 8260 30370 8316 30382
rect 7868 30268 8148 30324
rect 7774 30212 7830 30222
rect 7774 30118 7830 30156
rect 7028 29708 7252 29764
rect 6860 29596 7140 29652
rect 7084 28868 7140 29596
rect 7196 29314 7252 29708
rect 7196 29262 7198 29314
rect 7250 29262 7252 29314
rect 7196 29250 7252 29262
rect 7308 29441 7364 29453
rect 7308 29389 7310 29441
rect 7362 29389 7364 29441
rect 7308 29316 7364 29389
rect 7644 29426 7700 30044
rect 7644 29374 7646 29426
rect 7698 29374 7700 29426
rect 7644 29362 7700 29374
rect 7980 29652 8036 29662
rect 7308 29250 7364 29260
rect 7980 28868 8036 29596
rect 8092 29550 8148 30268
rect 8540 30154 8596 30166
rect 8540 30102 8542 30154
rect 8594 30102 8596 30154
rect 8540 30100 8596 30102
rect 8540 30034 8596 30044
rect 8092 29538 8204 29550
rect 8092 29486 8150 29538
rect 8202 29486 8204 29538
rect 8092 29484 8204 29486
rect 8148 29474 8204 29484
rect 8428 29426 8484 29438
rect 8428 29374 8430 29426
rect 8482 29374 8484 29426
rect 8428 28878 8484 29374
rect 8652 29428 8708 30940
rect 8764 30930 8820 30940
rect 9660 31332 9716 31342
rect 9660 30882 9716 31276
rect 9660 30830 9662 30882
rect 9714 30830 9716 30882
rect 9660 30818 9716 30830
rect 10052 30994 10108 31500
rect 10220 31164 10276 34748
rect 10892 34914 10948 34926
rect 10892 34862 10894 34914
rect 10946 34862 10948 34914
rect 10536 34524 10800 34534
rect 10592 34468 10640 34524
rect 10696 34468 10744 34524
rect 10536 34458 10800 34468
rect 10892 34354 10948 34862
rect 10892 34302 10894 34354
rect 10946 34302 10948 34354
rect 10892 34290 10948 34302
rect 11788 34157 11844 34169
rect 11788 34105 11790 34157
rect 11842 34105 11844 34157
rect 11228 33572 11284 33582
rect 10444 33460 10500 33470
rect 10444 33366 10500 33404
rect 10780 33348 10836 33358
rect 10780 33254 10836 33292
rect 11116 33124 11172 33134
rect 11116 33030 11172 33068
rect 10536 32956 10800 32966
rect 10592 32900 10640 32956
rect 10696 32900 10744 32956
rect 10536 32890 10800 32900
rect 10892 32900 10948 32910
rect 10892 32676 10948 32844
rect 11228 32676 11284 33516
rect 10332 32590 10388 32602
rect 10332 32538 10334 32590
rect 10386 32538 10388 32590
rect 10332 32228 10388 32538
rect 10500 32578 10556 32590
rect 10500 32526 10502 32578
rect 10554 32564 10556 32578
rect 10554 32526 10724 32564
rect 10500 32508 10724 32526
rect 10332 32162 10388 32172
rect 10668 32228 10724 32508
rect 10892 32562 10948 32620
rect 10892 32510 10894 32562
rect 10946 32510 10948 32562
rect 10892 32498 10948 32510
rect 11116 32620 11284 32676
rect 11340 33348 11396 33358
rect 11116 32564 11172 32620
rect 11116 32470 11172 32508
rect 11228 32452 11284 32462
rect 11228 32394 11284 32396
rect 11228 32342 11230 32394
rect 11282 32342 11284 32394
rect 11228 32330 11284 32342
rect 10668 32162 10724 32172
rect 10444 32116 10500 32126
rect 10444 32004 10500 32060
rect 11116 32004 11172 32014
rect 10444 32002 11172 32004
rect 10444 31950 11118 32002
rect 11170 31950 11172 32002
rect 10444 31948 11172 31950
rect 11116 31938 11172 31948
rect 10556 31780 10612 31790
rect 10332 31722 10388 31734
rect 10332 31670 10334 31722
rect 10386 31670 10388 31722
rect 10556 31698 10558 31724
rect 10610 31698 10612 31724
rect 10724 31762 11172 31780
rect 10724 31710 10726 31762
rect 10778 31724 11172 31762
rect 10778 31710 10780 31724
rect 10724 31698 10780 31710
rect 10556 31686 10612 31698
rect 10332 31332 10388 31670
rect 10536 31388 10800 31398
rect 10592 31332 10640 31388
rect 10696 31332 10744 31388
rect 10536 31322 10800 31332
rect 10332 31266 10388 31276
rect 10220 31108 10500 31164
rect 10052 30942 10054 30994
rect 10106 30942 10108 30994
rect 10052 30436 10108 30942
rect 10220 30994 10276 31006
rect 10220 30942 10222 30994
rect 10274 30942 10276 30994
rect 10220 30884 10276 30942
rect 10220 30818 10276 30828
rect 10332 30938 10388 30950
rect 10332 30886 10334 30938
rect 10386 30886 10388 30938
rect 9996 30380 10108 30436
rect 9548 30322 9604 30334
rect 9548 30270 9550 30322
rect 9602 30270 9604 30322
rect 8988 30212 9044 30222
rect 8764 30154 8820 30166
rect 8764 30102 8766 30154
rect 8818 30102 8820 30154
rect 8988 30130 8990 30156
rect 9042 30130 9044 30156
rect 8988 30118 9044 30130
rect 9100 30154 9156 30166
rect 8764 30100 8820 30102
rect 8764 30034 8820 30044
rect 9100 30102 9102 30154
rect 9154 30102 9156 30154
rect 8652 29426 8820 29428
rect 8652 29374 8654 29426
rect 8706 29374 8820 29426
rect 8652 29372 8820 29374
rect 8652 29362 8708 29372
rect 6748 28812 6916 28868
rect 6580 28754 6804 28756
rect 6580 28702 6582 28754
rect 6634 28702 6804 28754
rect 6580 28700 6804 28702
rect 6580 28690 6636 28700
rect 6748 28642 6804 28700
rect 6748 28590 6750 28642
rect 6802 28590 6804 28642
rect 6748 28578 6804 28590
rect 5874 27468 6138 27478
rect 5930 27412 5978 27468
rect 6034 27412 6082 27468
rect 5874 27402 6138 27412
rect 5292 26238 5294 26290
rect 5346 26238 5348 26290
rect 5292 26226 5348 26238
rect 5516 26852 5684 26908
rect 6860 26908 6916 28812
rect 7084 28866 7588 28868
rect 7084 28814 7086 28866
rect 7138 28814 7588 28866
rect 7084 28812 7588 28814
rect 7084 28802 7140 28812
rect 7532 27972 7588 28812
rect 7644 28756 7700 28766
rect 7644 28627 7700 28700
rect 7644 28575 7646 28627
rect 7698 28575 7700 28627
rect 7980 28642 8036 28812
rect 8372 28866 8484 28878
rect 8372 28814 8374 28866
rect 8426 28814 8484 28866
rect 8372 28812 8484 28814
rect 8540 29204 8596 29214
rect 8372 28802 8428 28812
rect 7980 28590 7982 28642
rect 8034 28590 8036 28642
rect 7980 28578 8036 28590
rect 8204 28644 8260 28654
rect 8540 28644 8596 29148
rect 8764 28980 8820 29372
rect 8764 28914 8820 28924
rect 7644 28563 7700 28575
rect 7644 28474 7700 28486
rect 7644 28422 7646 28474
rect 7698 28422 7700 28474
rect 7644 28308 7700 28422
rect 7644 28252 7868 28308
rect 7644 27972 7700 27982
rect 7532 27970 7700 27972
rect 7532 27918 7646 27970
rect 7698 27918 7700 27970
rect 7532 27916 7700 27918
rect 7644 27906 7700 27916
rect 7812 27914 7868 28252
rect 7812 27862 7814 27914
rect 7866 27862 7868 27914
rect 7812 27850 7868 27862
rect 8204 27298 8260 28588
rect 8428 28588 8596 28644
rect 8652 28868 8708 28878
rect 9100 28868 9156 30102
rect 9548 30100 9604 30270
rect 9548 30034 9604 30044
rect 9772 30324 9828 30334
rect 9548 29652 9604 29662
rect 9548 29426 9604 29596
rect 9548 29374 9550 29426
rect 9602 29374 9604 29426
rect 9548 29362 9604 29374
rect 9772 29428 9828 30268
rect 9996 30212 10052 30380
rect 9942 30156 10052 30212
rect 10108 30210 10164 30222
rect 10108 30158 10110 30210
rect 10162 30158 10164 30210
rect 9942 30154 9998 30156
rect 9942 30102 9944 30154
rect 9996 30102 9998 30154
rect 9942 29876 9998 30102
rect 9942 29820 10052 29876
rect 9772 29362 9828 29372
rect 9884 29540 9940 29550
rect 9884 29426 9940 29484
rect 9884 29374 9886 29426
rect 9938 29374 9940 29426
rect 9884 29362 9940 29374
rect 9660 29316 9716 29326
rect 9660 29258 9716 29260
rect 9660 29206 9662 29258
rect 9714 29206 9716 29258
rect 9660 29194 9716 29206
rect 9996 29204 10052 29820
rect 10108 29316 10164 30158
rect 10220 30212 10276 30222
rect 10332 30212 10388 30886
rect 10220 30210 10388 30212
rect 10220 30158 10222 30210
rect 10274 30158 10388 30210
rect 10220 30156 10388 30158
rect 10444 30210 10500 31108
rect 10444 30158 10446 30210
rect 10498 30158 10500 30210
rect 10220 30100 10276 30156
rect 10444 30146 10500 30158
rect 10220 30034 10276 30044
rect 10780 29988 10836 29998
rect 10780 29986 11060 29988
rect 10780 29934 10782 29986
rect 10834 29934 11060 29986
rect 10780 29932 11060 29934
rect 10780 29922 10836 29932
rect 11004 29876 11060 29932
rect 10536 29820 10800 29830
rect 10592 29764 10640 29820
rect 10696 29764 10744 29820
rect 11004 29810 11060 29820
rect 10536 29754 10800 29764
rect 10780 29428 10836 29438
rect 10780 29334 10836 29372
rect 10892 29426 10948 29438
rect 10892 29374 10894 29426
rect 10946 29374 10948 29426
rect 10108 29250 10164 29260
rect 9996 29138 10052 29148
rect 10444 29204 10500 29214
rect 10444 29110 10500 29148
rect 10892 29092 10948 29374
rect 10892 29026 10948 29036
rect 9436 28980 9492 28990
rect 9212 28868 9268 28878
rect 9100 28812 9212 28868
rect 8652 28614 8708 28812
rect 8204 27246 8206 27298
rect 8258 27246 8260 27298
rect 8204 27234 8260 27246
rect 8316 27858 8372 27870
rect 8316 27806 8318 27858
rect 8370 27806 8372 27858
rect 6860 26852 7028 26908
rect 5516 26292 5572 26852
rect 5516 26226 5572 26236
rect 6972 26404 7028 26852
rect 7196 26404 7252 26414
rect 6972 26402 7252 26404
rect 6972 26350 7198 26402
rect 7250 26350 7252 26402
rect 6972 26348 7252 26350
rect 5874 25900 6138 25910
rect 5930 25844 5978 25900
rect 6034 25844 6082 25900
rect 5874 25834 6138 25844
rect 6188 25620 6244 25630
rect 4956 25508 5012 25518
rect 4844 25506 5012 25508
rect 4844 25454 4958 25506
rect 5010 25454 5012 25506
rect 4844 25452 5012 25454
rect 4396 25228 4564 25284
rect 4956 25284 5012 25452
rect 5180 25508 5236 25518
rect 5946 25508 6002 25518
rect 5180 25506 6002 25508
rect 5180 25454 5182 25506
rect 5234 25454 5948 25506
rect 6000 25454 6002 25506
rect 5180 25452 6002 25454
rect 5180 25442 5236 25452
rect 5946 25442 6002 25452
rect 6188 25506 6244 25564
rect 6972 25620 7028 26348
rect 7196 26338 7252 26348
rect 7812 26180 7868 26190
rect 6972 25554 7028 25564
rect 7756 26178 7868 26180
rect 7756 26126 7814 26178
rect 7866 26126 7868 26178
rect 7756 26114 7868 26126
rect 6188 25454 6190 25506
rect 6242 25454 6244 25506
rect 6188 25442 6244 25454
rect 6692 25508 6748 25546
rect 6692 25442 6748 25452
rect 7196 25508 7252 25518
rect 6636 25338 6692 25350
rect 4340 25190 4396 25228
rect 4956 25218 5012 25228
rect 5740 25284 5796 25294
rect 3836 24162 4116 24164
rect 3836 24110 3838 24162
rect 3890 24110 4116 24162
rect 3836 24108 4116 24110
rect 4732 25060 4788 25070
rect 4732 24834 4788 25004
rect 4732 24782 4734 24834
rect 4786 24782 4788 24834
rect 3836 24098 3892 24108
rect 4732 23716 4788 24782
rect 5068 24948 5124 24958
rect 4956 24724 5012 24734
rect 4956 23940 5012 24668
rect 5068 24722 5124 24892
rect 5572 24836 5628 24846
rect 5572 24742 5628 24780
rect 5068 24670 5070 24722
rect 5122 24670 5124 24722
rect 5068 24658 5124 24670
rect 5292 24722 5348 24734
rect 5292 24670 5294 24722
rect 5346 24670 5348 24722
rect 4956 23938 5236 23940
rect 4956 23886 4958 23938
rect 5010 23886 5236 23938
rect 4956 23884 5236 23886
rect 4956 23874 5012 23884
rect 4732 23650 4788 23660
rect 2940 23380 2996 23390
rect 2940 22370 2996 23324
rect 4284 23380 4340 23390
rect 4284 23286 4340 23324
rect 4844 23380 4900 23390
rect 4620 23154 4676 23166
rect 4620 23102 4622 23154
rect 4674 23102 4676 23154
rect 4620 23044 4676 23102
rect 4620 22978 4676 22988
rect 2940 22318 2942 22370
rect 2994 22318 2996 22370
rect 2940 22306 2996 22318
rect 3164 22370 3220 22382
rect 3164 22318 3166 22370
rect 3218 22318 3220 22370
rect 2660 22260 2716 22270
rect 2044 21588 2100 22092
rect 2492 22258 2716 22260
rect 2492 22206 2662 22258
rect 2714 22206 2716 22258
rect 2492 22204 2716 22206
rect 2044 21586 2212 21588
rect 2044 21534 2046 21586
rect 2098 21534 2212 21586
rect 2044 21532 2212 21534
rect 2044 21522 2100 21532
rect 2044 20804 2100 20814
rect 2044 20710 2100 20748
rect 2156 20020 2212 21532
rect 2492 20804 2548 22204
rect 2660 22194 2716 22204
rect 3164 21812 3220 22318
rect 3164 21746 3220 21756
rect 4060 22258 4116 22270
rect 4060 22206 4062 22258
rect 4114 22206 4116 22258
rect 4060 21700 4116 22206
rect 4060 21634 4116 21644
rect 2828 21474 2884 21486
rect 2828 21422 2830 21474
rect 2882 21422 2884 21474
rect 2828 21028 2884 21422
rect 4732 21476 4788 21486
rect 4732 21382 4788 21420
rect 3164 21028 3220 21038
rect 2828 21026 3220 21028
rect 2828 20974 3166 21026
rect 3218 20974 3220 21026
rect 2828 20972 3220 20974
rect 3164 20962 3220 20972
rect 4844 20916 4900 23324
rect 5012 23044 5068 23054
rect 5012 22950 5068 22988
rect 5180 22370 5236 23884
rect 5292 23380 5348 24670
rect 5740 24162 5796 25228
rect 6636 25286 6638 25338
rect 6690 25286 6692 25338
rect 6636 24612 6692 25286
rect 6636 24518 6692 24556
rect 7084 24500 7140 24510
rect 5874 24332 6138 24342
rect 5930 24276 5978 24332
rect 6034 24276 6082 24332
rect 5874 24266 6138 24276
rect 5740 24110 5742 24162
rect 5794 24110 5796 24162
rect 5740 24098 5796 24110
rect 6076 23938 6132 23950
rect 6076 23886 6078 23938
rect 6130 23886 6132 23938
rect 5292 23314 5348 23324
rect 5740 23716 5796 23726
rect 5180 22318 5182 22370
rect 5234 22318 5236 22370
rect 5180 22306 5236 22318
rect 5740 22372 5796 23660
rect 6076 23716 6132 23886
rect 6468 23716 6524 23726
rect 6076 23714 6524 23716
rect 6076 23662 6470 23714
rect 6522 23662 6524 23714
rect 6076 23660 6524 23662
rect 6076 23044 6132 23660
rect 6468 23650 6524 23660
rect 6244 23268 6300 23278
rect 6244 23174 6300 23212
rect 6860 23268 6916 23278
rect 6580 23156 6636 23166
rect 6580 23062 6636 23100
rect 6860 23154 6916 23212
rect 6860 23102 6862 23154
rect 6914 23102 6916 23154
rect 6860 23090 6916 23102
rect 7084 23154 7140 24444
rect 7196 24050 7252 25452
rect 7196 23998 7198 24050
rect 7250 23998 7252 24050
rect 7196 23986 7252 23998
rect 7420 25508 7476 25518
rect 7756 25508 7812 26114
rect 7420 25506 7812 25508
rect 7420 25454 7422 25506
rect 7474 25454 7812 25506
rect 7420 25452 7812 25454
rect 8316 25508 8372 27806
rect 8428 27076 8484 28588
rect 8652 28562 8654 28614
rect 8706 28562 8708 28614
rect 8652 28550 8708 28562
rect 8876 28644 8932 28654
rect 9212 28607 9268 28812
rect 8876 28562 8878 28588
rect 8930 28562 8932 28588
rect 8876 28550 8932 28562
rect 9044 28586 9100 28598
rect 9044 28534 9046 28586
rect 9098 28534 9100 28586
rect 9212 28555 9214 28607
rect 9266 28555 9268 28607
rect 9212 28543 9268 28555
rect 9044 28532 9100 28534
rect 8988 28476 9100 28532
rect 8558 27972 8614 27982
rect 8988 27972 9044 28476
rect 8558 27970 9044 27972
rect 8558 27918 8560 27970
rect 8612 27918 9044 27970
rect 8558 27916 9044 27918
rect 8558 27906 8614 27916
rect 9100 27188 9156 27198
rect 8596 27076 8652 27086
rect 8428 27074 8652 27076
rect 8428 27022 8598 27074
rect 8650 27022 8652 27074
rect 8428 27020 8652 27022
rect 8596 27010 8652 27020
rect 8764 27074 8820 27086
rect 8764 27022 8766 27074
rect 8818 27022 8820 27074
rect 8764 26964 8820 27022
rect 8876 27076 8932 27086
rect 8876 26982 8932 27020
rect 9100 27074 9156 27132
rect 9100 27022 9102 27074
rect 9154 27022 9156 27074
rect 9100 27010 9156 27022
rect 8764 26898 8820 26908
rect 7084 23102 7086 23154
rect 7138 23102 7140 23154
rect 7084 23090 7140 23102
rect 7196 23156 7252 23166
rect 7196 23062 7252 23100
rect 6076 22978 6132 22988
rect 5874 22764 6138 22774
rect 5930 22708 5978 22764
rect 6034 22708 6082 22764
rect 5874 22698 6138 22708
rect 5740 22316 6020 22372
rect 5796 22148 5852 22158
rect 5796 22054 5852 22092
rect 5964 21924 6020 22316
rect 7420 22158 7476 25452
rect 7756 24724 7812 24734
rect 7756 24630 7812 24668
rect 8316 24722 8372 25452
rect 8316 24670 8318 24722
rect 8370 24670 8372 24722
rect 8988 24722 9044 24734
rect 8316 24658 8372 24670
rect 8820 24666 8876 24678
rect 8820 24614 8822 24666
rect 8874 24614 8876 24666
rect 8074 24500 8130 24510
rect 8074 24406 8130 24444
rect 8820 24388 8876 24614
rect 8988 24670 8990 24722
rect 9042 24670 9044 24722
rect 8988 24612 9044 24670
rect 8988 24500 9044 24556
rect 8988 24444 9380 24500
rect 8820 24332 9268 24388
rect 9100 23940 9156 23950
rect 8876 23938 9156 23940
rect 8876 23886 9102 23938
rect 9154 23886 9156 23938
rect 8876 23884 9156 23886
rect 8652 23380 8708 23390
rect 8876 23380 8932 23884
rect 9100 23874 9156 23884
rect 8652 23378 8932 23380
rect 8652 23326 8654 23378
rect 8706 23326 8932 23378
rect 8652 23324 8932 23326
rect 8652 23314 8708 23324
rect 7980 23268 8036 23278
rect 7980 22708 8036 23212
rect 9212 23156 9268 24332
rect 9324 23828 9380 24444
rect 9324 23762 9380 23772
rect 9436 23380 9492 28924
rect 10892 28868 10948 28878
rect 11116 28868 11172 31724
rect 11340 30996 11396 33292
rect 11452 33346 11508 33358
rect 11452 33294 11454 33346
rect 11506 33294 11508 33346
rect 11452 32676 11508 33294
rect 11676 32676 11732 32686
rect 11452 32620 11676 32676
rect 11676 32562 11732 32620
rect 11676 32510 11678 32562
rect 11730 32510 11732 32562
rect 11676 32498 11732 32510
rect 11676 32340 11732 32350
rect 11676 31778 11732 32284
rect 11788 32004 11844 34105
rect 12012 33572 12068 35420
rect 12236 35410 12292 35420
rect 12348 35698 12404 35710
rect 12348 35646 12350 35698
rect 12402 35646 12404 35698
rect 12348 35252 12404 35646
rect 12348 34916 12404 35196
rect 12348 34850 12404 34860
rect 12572 34018 12628 37324
rect 13244 36484 13300 39200
rect 13244 36418 13300 36428
rect 13692 36482 13748 36494
rect 13692 36430 13694 36482
rect 13746 36430 13748 36482
rect 13356 36258 13412 36270
rect 13356 36206 13358 36258
rect 13410 36206 13412 36258
rect 13356 35700 13412 36206
rect 13692 35924 13748 36430
rect 13916 36454 13972 36466
rect 13916 36402 13918 36454
rect 13970 36402 13972 36454
rect 13916 36260 13972 36402
rect 13916 36194 13972 36204
rect 13692 35868 14308 35924
rect 13132 35586 13188 35598
rect 13132 35534 13134 35586
rect 13186 35534 13188 35586
rect 12796 35476 12852 35486
rect 12796 35026 12852 35420
rect 12796 34974 12798 35026
rect 12850 34974 12852 35026
rect 12796 34962 12852 34974
rect 12572 33966 12574 34018
rect 12626 33966 12628 34018
rect 12572 33954 12628 33966
rect 12012 33506 12068 33516
rect 12460 33572 12516 33582
rect 12348 33458 12404 33470
rect 12348 33406 12350 33458
rect 12402 33406 12404 33458
rect 11900 33348 11956 33358
rect 11900 33346 12180 33348
rect 11900 33294 11902 33346
rect 11954 33294 12180 33346
rect 11900 33292 12180 33294
rect 11900 33282 11956 33292
rect 11900 32577 11956 32589
rect 11900 32525 11902 32577
rect 11954 32525 11956 32577
rect 11900 32452 11956 32525
rect 12124 32564 12180 33292
rect 12236 33290 12292 33302
rect 12236 33238 12238 33290
rect 12290 33238 12292 33290
rect 12236 33012 12292 33238
rect 12236 32946 12292 32956
rect 12348 32676 12404 33406
rect 12460 33346 12516 33516
rect 12460 33294 12462 33346
rect 12514 33294 12516 33346
rect 12460 33236 12516 33294
rect 12460 33170 12516 33180
rect 12348 32610 12404 32620
rect 12908 33012 12964 33022
rect 12124 32508 12292 32564
rect 11900 32386 11956 32396
rect 12012 32452 12068 32462
rect 12012 32450 12180 32452
rect 12012 32398 12014 32450
rect 12066 32398 12180 32450
rect 12012 32396 12180 32398
rect 12012 32386 12068 32396
rect 11788 31948 12068 32004
rect 11508 31722 11564 31734
rect 11508 31670 11510 31722
rect 11562 31670 11564 31722
rect 11676 31726 11678 31778
rect 11730 31726 11732 31778
rect 11676 31714 11732 31726
rect 11788 31778 11844 31790
rect 11788 31726 11790 31778
rect 11842 31726 11844 31778
rect 11508 31556 11564 31670
rect 11508 31490 11564 31500
rect 11658 31220 11714 31230
rect 11658 31106 11714 31164
rect 11658 31054 11660 31106
rect 11712 31054 11714 31106
rect 11658 31042 11714 31054
rect 11340 30940 11620 30996
rect 11228 29988 11284 29998
rect 11228 29650 11284 29932
rect 11396 29988 11452 29998
rect 11396 29986 11508 29988
rect 11396 29934 11398 29986
rect 11450 29934 11508 29986
rect 11396 29922 11508 29934
rect 11228 29598 11230 29650
rect 11282 29598 11284 29650
rect 11228 29586 11284 29598
rect 11452 29092 11508 29922
rect 11452 29026 11508 29036
rect 11340 28868 11396 28878
rect 10948 28866 11396 28868
rect 10948 28814 11342 28866
rect 11394 28814 11396 28866
rect 10948 28812 11396 28814
rect 10220 28756 10276 28766
rect 9884 28754 10276 28756
rect 9884 28702 10222 28754
rect 10274 28702 10276 28754
rect 9884 28700 10276 28702
rect 9716 28644 9772 28654
rect 9716 28082 9772 28588
rect 9716 28030 9718 28082
rect 9770 28030 9772 28082
rect 9716 27076 9772 28030
rect 9884 28084 9940 28700
rect 10220 28690 10276 28700
rect 10444 28644 10500 28654
rect 10052 28586 10108 28598
rect 10052 28534 10054 28586
rect 10106 28534 10108 28586
rect 10444 28550 10500 28588
rect 10780 28586 10836 28598
rect 10052 28084 10108 28534
rect 10780 28534 10782 28586
rect 10834 28534 10836 28586
rect 10780 28420 10836 28534
rect 10780 28354 10836 28364
rect 10536 28252 10800 28262
rect 10592 28196 10640 28252
rect 10696 28196 10744 28252
rect 10536 28186 10800 28196
rect 10892 28084 10948 28812
rect 11340 28802 11396 28812
rect 11564 28420 11620 30940
rect 11788 30212 11844 31726
rect 11900 30994 11956 31006
rect 11900 30942 11902 30994
rect 11954 30942 11956 30994
rect 11900 30324 11956 30942
rect 11900 30258 11956 30268
rect 11676 30156 11844 30212
rect 11676 29988 11732 30156
rect 11676 29922 11732 29932
rect 11844 29986 11900 29998
rect 11844 29934 11846 29986
rect 11898 29934 11900 29986
rect 11844 29764 11900 29934
rect 11844 29698 11900 29708
rect 11676 28868 11732 28878
rect 11676 28642 11732 28812
rect 11676 28590 11678 28642
rect 11730 28590 11732 28642
rect 11676 28578 11732 28590
rect 11788 28644 11844 28654
rect 12012 28644 12068 31948
rect 12124 31780 12180 32396
rect 12124 31686 12180 31724
rect 12236 30548 12292 32508
rect 12684 31892 12740 31902
rect 12684 31778 12740 31836
rect 12684 31726 12686 31778
rect 12738 31726 12740 31778
rect 12684 31714 12740 31726
rect 12796 31668 12852 31678
rect 12572 31610 12628 31622
rect 12572 31558 12574 31610
rect 12626 31558 12628 31610
rect 12572 31332 12628 31558
rect 12404 31276 12628 31332
rect 12684 31556 12740 31566
rect 12404 31050 12460 31276
rect 12404 30998 12406 31050
rect 12458 30998 12460 31050
rect 12404 30986 12460 30998
rect 12572 30994 12628 31006
rect 12236 30482 12292 30492
rect 12572 30942 12574 30994
rect 12626 30942 12628 30994
rect 12236 30212 12292 30222
rect 12124 30154 12180 30166
rect 12124 30102 12126 30154
rect 12178 30102 12180 30154
rect 12236 30118 12292 30156
rect 12404 30154 12460 30166
rect 12124 29988 12180 30102
rect 12124 29922 12180 29932
rect 12404 30102 12406 30154
rect 12458 30102 12460 30154
rect 12404 29764 12460 30102
rect 12404 29698 12460 29708
rect 12572 30100 12628 30942
rect 12124 29652 12180 29662
rect 12124 29558 12180 29596
rect 12236 29540 12292 29550
rect 11788 28642 12068 28644
rect 11788 28590 11790 28642
rect 11842 28590 12068 28642
rect 11788 28588 12068 28590
rect 12124 28868 12180 28878
rect 12236 28868 12292 29484
rect 12124 28866 12292 28868
rect 12124 28814 12126 28866
rect 12178 28814 12292 28866
rect 12124 28812 12292 28814
rect 12460 29426 12516 29438
rect 12460 29374 12462 29426
rect 12514 29374 12516 29426
rect 12460 28868 12516 29374
rect 12572 29428 12628 30044
rect 12684 29652 12740 31500
rect 12796 30434 12852 31612
rect 12796 30382 12798 30434
rect 12850 30382 12852 30434
rect 12796 30370 12852 30382
rect 12908 29876 12964 32956
rect 13020 32788 13076 32798
rect 13132 32788 13188 35534
rect 13020 32786 13188 32788
rect 13020 32734 13022 32786
rect 13074 32734 13188 32786
rect 13020 32732 13188 32734
rect 13020 32722 13076 32732
rect 13356 32564 13412 35644
rect 14252 35252 14308 35868
rect 14252 35186 14308 35196
rect 14364 35140 14420 39200
rect 15484 37044 15540 39200
rect 16604 37828 16660 39200
rect 17724 39060 17780 39200
rect 17948 39060 18004 39228
rect 17724 39004 18004 39060
rect 16156 37772 16660 37828
rect 15484 36988 16100 37044
rect 15198 36876 15462 36886
rect 15254 36820 15302 36876
rect 15358 36820 15406 36876
rect 15198 36810 15462 36820
rect 16044 36148 16100 36988
rect 16156 36482 16212 37772
rect 16156 36430 16158 36482
rect 16210 36430 16212 36482
rect 16156 36418 16212 36430
rect 17388 36482 17444 36494
rect 17388 36430 17390 36482
rect 17442 36430 17444 36482
rect 17052 36260 17108 36270
rect 16716 36258 17108 36260
rect 16716 36206 17054 36258
rect 17106 36206 17108 36258
rect 16716 36204 17108 36206
rect 16044 36092 16212 36148
rect 15708 35700 15764 35710
rect 15708 35698 15876 35700
rect 15708 35646 15710 35698
rect 15762 35646 15876 35698
rect 15708 35644 15876 35646
rect 15708 35634 15764 35644
rect 14364 35074 14420 35084
rect 15036 35586 15092 35598
rect 15036 35534 15038 35586
rect 15090 35534 15092 35586
rect 15036 35252 15092 35534
rect 15596 35588 15652 35598
rect 15198 35308 15462 35318
rect 15254 35252 15302 35308
rect 15358 35252 15406 35308
rect 15198 35242 15462 35252
rect 13748 34916 13804 34926
rect 13748 34822 13804 34860
rect 13916 34914 13972 34926
rect 13916 34862 13918 34914
rect 13970 34862 13972 34914
rect 13916 33572 13972 34862
rect 14364 34157 14420 34169
rect 14364 34105 14366 34157
rect 14418 34105 14420 34157
rect 14364 33796 14420 34105
rect 15036 33908 15092 35196
rect 15372 35140 15428 35150
rect 15596 35140 15652 35532
rect 15820 35476 15876 35644
rect 15372 35138 15652 35140
rect 15372 35086 15374 35138
rect 15426 35086 15652 35138
rect 15372 35084 15652 35086
rect 15708 35140 15764 35150
rect 15372 35074 15428 35084
rect 15708 34354 15764 35084
rect 15708 34302 15710 34354
rect 15762 34302 15764 34354
rect 15708 34290 15764 34302
rect 15036 33842 15092 33852
rect 14364 33730 14420 33740
rect 15198 33740 15462 33750
rect 15254 33684 15302 33740
rect 15358 33684 15406 33740
rect 15198 33674 15462 33684
rect 14756 33572 14812 33582
rect 15820 33572 15876 35420
rect 16044 35698 16100 35710
rect 16044 35646 16046 35698
rect 16098 35646 16100 35698
rect 15932 34916 15988 34926
rect 15932 34692 15988 34860
rect 15932 34626 15988 34636
rect 13916 33570 14812 33572
rect 13916 33518 14758 33570
rect 14810 33518 14812 33570
rect 13916 33516 14812 33518
rect 14756 33506 14812 33516
rect 15484 33516 15876 33572
rect 15932 34356 15988 34366
rect 13804 33346 13860 33358
rect 13804 33294 13806 33346
rect 13858 33294 13860 33346
rect 13524 33236 13580 33246
rect 13524 33234 13748 33236
rect 13524 33182 13526 33234
rect 13578 33182 13748 33234
rect 13524 33180 13748 33182
rect 13524 33170 13580 33180
rect 13692 32564 13748 33180
rect 13804 32788 13860 33294
rect 13916 33348 13972 33358
rect 13916 33254 13972 33292
rect 14252 33348 14308 33358
rect 14252 33254 14308 33292
rect 14476 33346 14532 33358
rect 14476 33294 14478 33346
rect 14530 33294 14532 33346
rect 13804 32732 14308 32788
rect 14140 32564 14196 32574
rect 13692 32562 14196 32564
rect 13692 32510 14142 32562
rect 14194 32510 14196 32562
rect 13692 32508 14196 32510
rect 13356 32498 13412 32508
rect 14140 32498 14196 32508
rect 14028 32340 14084 32350
rect 14028 31892 14084 32284
rect 14252 32014 14308 32732
rect 14364 32564 14420 32574
rect 14364 32470 14420 32508
rect 14252 32002 14364 32014
rect 14252 31950 14310 32002
rect 14362 31950 14364 32002
rect 14252 31948 14364 31950
rect 14308 31938 14364 31948
rect 13692 31780 13748 31790
rect 13468 31722 13524 31734
rect 13468 31670 13470 31722
rect 13522 31670 13524 31722
rect 13468 31556 13524 31670
rect 13468 31490 13524 31500
rect 13580 31722 13636 31734
rect 13580 31670 13582 31722
rect 13634 31670 13636 31722
rect 13580 31220 13636 31670
rect 13580 31154 13636 31164
rect 14028 31750 14084 31836
rect 13020 31108 13076 31118
rect 13076 31052 13188 31108
rect 13020 31042 13076 31052
rect 12908 29810 12964 29820
rect 12684 29586 12740 29596
rect 13132 29494 13188 31052
rect 13244 30994 13300 31006
rect 13244 30942 13246 30994
rect 13298 30942 13300 30994
rect 13244 29876 13300 30942
rect 13356 30994 13412 31006
rect 13356 30942 13358 30994
rect 13410 30942 13412 30994
rect 13356 30548 13412 30942
rect 13524 30994 13580 31006
rect 13524 30942 13526 30994
rect 13578 30942 13580 30994
rect 13524 30660 13580 30942
rect 13524 30594 13580 30604
rect 13356 30482 13412 30492
rect 13524 30378 13580 30390
rect 13524 30326 13526 30378
rect 13578 30326 13580 30378
rect 13524 30212 13580 30326
rect 13524 30146 13580 30156
rect 13692 30210 13748 31724
rect 13804 31722 13860 31734
rect 13804 31670 13806 31722
rect 13858 31670 13860 31722
rect 14028 31698 14030 31750
rect 14082 31698 14084 31750
rect 14028 31686 14084 31698
rect 13804 31668 13860 31670
rect 13804 31602 13860 31612
rect 14364 31556 14420 31566
rect 13692 30158 13694 30210
rect 13746 30158 13748 30210
rect 13692 30146 13748 30158
rect 13804 31220 13860 31230
rect 13244 29810 13300 29820
rect 13804 29540 13860 31164
rect 14364 31050 14420 31500
rect 14476 31444 14532 33294
rect 15484 33318 15540 33516
rect 15932 33460 15988 34300
rect 15484 33266 15486 33318
rect 15538 33266 15540 33318
rect 15484 33254 15540 33266
rect 15708 33404 15988 33460
rect 14700 32564 14756 32574
rect 14700 32562 14980 32564
rect 14700 32510 14702 32562
rect 14754 32510 14980 32562
rect 14700 32508 14980 32510
rect 14700 32498 14756 32508
rect 14700 32394 14756 32406
rect 14700 32342 14702 32394
rect 14754 32342 14756 32394
rect 14476 31378 14532 31388
rect 14588 31778 14644 31790
rect 14588 31726 14590 31778
rect 14642 31726 14644 31778
rect 14588 31332 14644 31726
rect 14700 31556 14756 32342
rect 14812 32340 14868 32350
rect 14812 31778 14868 32284
rect 14812 31726 14814 31778
rect 14866 31726 14868 31778
rect 14812 31714 14868 31726
rect 14924 31780 14980 32508
rect 15708 32562 15764 33404
rect 16044 32900 16100 35646
rect 16156 33570 16212 36092
rect 16268 35737 16324 35749
rect 16268 35700 16270 35737
rect 16322 35700 16324 35737
rect 16268 35634 16324 35644
rect 16604 35698 16660 35710
rect 16604 35646 16606 35698
rect 16658 35646 16660 35698
rect 16156 33518 16158 33570
rect 16210 33518 16212 33570
rect 16156 33506 16212 33518
rect 16492 35586 16548 35598
rect 16492 35534 16494 35586
rect 16546 35534 16548 35586
rect 16044 32834 16100 32844
rect 15708 32510 15710 32562
rect 15762 32510 15764 32562
rect 15708 32498 15764 32510
rect 15932 32577 15988 32589
rect 15932 32525 15934 32577
rect 15986 32525 15988 32577
rect 15316 32452 15372 32462
rect 15260 32450 15372 32452
rect 15260 32398 15318 32450
rect 15370 32398 15372 32450
rect 15260 32386 15372 32398
rect 15260 32340 15316 32386
rect 15036 32284 15316 32340
rect 15036 31892 15092 32284
rect 15198 32172 15462 32182
rect 15254 32116 15302 32172
rect 15358 32116 15406 32172
rect 15198 32106 15462 32116
rect 15932 31948 15988 32525
rect 16492 32577 16548 35534
rect 16604 34804 16660 35646
rect 16716 35026 16772 36204
rect 17052 36194 17108 36204
rect 17276 35698 17332 35710
rect 17276 35646 17278 35698
rect 17330 35646 17332 35698
rect 17276 35252 17332 35646
rect 17388 35364 17444 36430
rect 18060 35588 18116 35598
rect 18060 35494 18116 35532
rect 17388 35308 18004 35364
rect 16716 34974 16718 35026
rect 16770 34974 16772 35026
rect 16716 34962 16772 34974
rect 16940 35196 17332 35252
rect 16604 34356 16660 34748
rect 16940 34692 16996 35196
rect 16940 34626 16996 34636
rect 17276 34692 17332 34702
rect 16604 34290 16660 34300
rect 16828 33572 16884 33582
rect 16492 32525 16494 32577
rect 16546 32525 16548 32577
rect 16044 32452 16100 32462
rect 16044 32358 16100 32396
rect 16380 32450 16436 32462
rect 16380 32398 16382 32450
rect 16434 32398 16436 32450
rect 15036 31826 15092 31836
rect 15820 31892 15876 31902
rect 15932 31892 16212 31948
rect 14924 31714 14980 31724
rect 15820 31778 15876 31836
rect 15820 31726 15822 31778
rect 15874 31726 15876 31778
rect 15820 31714 15876 31726
rect 15932 31778 15988 31790
rect 15932 31726 15934 31778
rect 15986 31726 15988 31778
rect 15092 31668 15148 31678
rect 14700 31490 14756 31500
rect 15036 31666 15148 31668
rect 15036 31614 15094 31666
rect 15146 31614 15148 31666
rect 15036 31602 15148 31614
rect 15540 31666 15596 31678
rect 15540 31614 15542 31666
rect 15594 31614 15596 31666
rect 14588 31266 14644 31276
rect 14364 30998 14366 31050
rect 14418 30998 14420 31050
rect 14364 30986 14420 30998
rect 14476 31220 14532 31230
rect 14476 31050 14532 31164
rect 14476 30998 14478 31050
rect 14530 30998 14532 31050
rect 14476 30986 14532 30998
rect 14700 31022 14756 31034
rect 14700 30970 14702 31022
rect 14754 30970 14756 31022
rect 13916 30884 13972 30894
rect 14700 30884 14756 30970
rect 14924 31022 14980 31034
rect 14924 30996 14926 31022
rect 14978 30996 14980 31022
rect 14924 30930 14980 30940
rect 13916 30882 14756 30884
rect 13916 30830 13918 30882
rect 13970 30830 14756 30882
rect 13916 30828 14756 30830
rect 13916 30818 13972 30828
rect 14364 30660 14420 30670
rect 14196 30548 14252 30558
rect 14196 30266 14252 30492
rect 14196 30214 14198 30266
rect 14250 30214 14252 30266
rect 14196 30202 14252 30214
rect 14028 30100 14084 30110
rect 14028 30006 14084 30044
rect 14364 29764 14420 30604
rect 15036 30548 15092 31602
rect 15204 31444 15260 31454
rect 15204 31106 15260 31388
rect 15204 31054 15206 31106
rect 15258 31054 15260 31106
rect 15204 31042 15260 31054
rect 15540 31108 15596 31614
rect 15540 31042 15596 31052
rect 15708 31556 15764 31566
rect 15708 31050 15764 31500
rect 15708 30998 15710 31050
rect 15762 30998 15764 31050
rect 15708 30986 15764 30998
rect 15198 30604 15462 30614
rect 15254 30548 15302 30604
rect 15358 30548 15406 30604
rect 15198 30538 15462 30548
rect 15036 30436 15092 30492
rect 15260 30436 15316 30446
rect 15036 30380 15204 30436
rect 14942 30324 14998 30334
rect 14942 30230 14998 30268
rect 14700 30212 14756 30222
rect 13934 29540 13990 29550
rect 13804 29538 13990 29540
rect 13132 29482 13244 29494
rect 13804 29486 13936 29538
rect 13988 29486 13990 29538
rect 13804 29484 13990 29486
rect 13020 29428 13076 29438
rect 13132 29430 13190 29482
rect 13242 29430 13244 29482
rect 13934 29474 13990 29484
rect 13132 29428 13244 29430
rect 12572 29426 13076 29428
rect 12572 29374 13022 29426
rect 13074 29374 13076 29426
rect 13188 29418 13244 29428
rect 13356 29428 13412 29438
rect 13692 29428 13748 29438
rect 12572 29372 13076 29374
rect 11564 28364 11732 28420
rect 9884 28028 9996 28084
rect 10052 28028 10220 28084
rect 9940 27972 9996 28028
rect 9940 27916 10052 27972
rect 9828 27860 9884 27870
rect 9828 27766 9884 27804
rect 9996 27636 10052 27916
rect 10164 27970 10220 28028
rect 10164 27918 10166 27970
rect 10218 27918 10220 27970
rect 10164 27906 10220 27918
rect 10556 28028 10948 28084
rect 10556 27970 10612 28028
rect 10556 27918 10558 27970
rect 10610 27918 10612 27970
rect 10556 27906 10612 27918
rect 9884 27580 10052 27636
rect 10444 27858 10500 27870
rect 10444 27806 10446 27858
rect 10498 27806 10500 27858
rect 9884 27186 9940 27580
rect 10444 27412 10500 27806
rect 10724 27860 10780 27870
rect 10724 27766 10780 27804
rect 10892 27858 10948 27870
rect 10892 27806 10894 27858
rect 10946 27806 10948 27858
rect 10108 27356 10500 27412
rect 10892 27412 10948 27806
rect 9884 27134 9886 27186
rect 9938 27134 9940 27186
rect 9884 27122 9940 27134
rect 9996 27188 10052 27198
rect 9716 27010 9772 27020
rect 9660 26068 9716 26078
rect 9660 25478 9716 26012
rect 9660 25426 9662 25478
rect 9714 25426 9716 25478
rect 9660 25414 9716 25426
rect 9996 24052 10052 27132
rect 10108 26852 10164 27356
rect 10892 27346 10948 27356
rect 11228 27858 11284 27870
rect 11228 27806 11230 27858
rect 11282 27806 11284 27858
rect 10108 26796 10388 26852
rect 10332 26122 10388 26796
rect 11228 26740 11284 27806
rect 10536 26684 10800 26694
rect 10592 26628 10640 26684
rect 10696 26628 10744 26684
rect 10536 26618 10800 26628
rect 10892 26684 11284 26740
rect 11340 27858 11396 27870
rect 11340 27806 11342 27858
rect 11394 27806 11396 27858
rect 11340 26740 11396 27806
rect 11508 27860 11564 27870
rect 11508 27766 11564 27804
rect 11564 27412 11620 27422
rect 11340 26684 11508 26740
rect 10444 26404 10500 26414
rect 10444 26290 10500 26348
rect 10668 26292 10724 26302
rect 10444 26238 10446 26290
rect 10498 26238 10500 26290
rect 10444 26226 10500 26238
rect 10556 26290 10724 26292
rect 10556 26238 10670 26290
rect 10722 26238 10724 26290
rect 10556 26236 10724 26238
rect 10164 26068 10220 26078
rect 10332 26070 10334 26122
rect 10386 26070 10388 26122
rect 10332 26058 10388 26070
rect 10164 25618 10220 26012
rect 10164 25566 10166 25618
rect 10218 25566 10220 25618
rect 10164 25554 10220 25566
rect 10556 25508 10612 26236
rect 10668 26226 10724 26236
rect 10892 26068 10948 26684
rect 11284 26516 11340 26526
rect 11284 26422 11340 26460
rect 11452 26404 11508 26684
rect 11564 26516 11620 27356
rect 11564 26450 11620 26460
rect 11452 26338 11508 26348
rect 10724 26012 10948 26068
rect 10724 25730 10780 26012
rect 10724 25678 10726 25730
rect 10778 25678 10780 25730
rect 10724 25666 10780 25678
rect 11004 25508 11060 25518
rect 10556 25506 10948 25508
rect 10556 25454 10558 25506
rect 10610 25454 10948 25506
rect 10556 25452 10948 25454
rect 10556 25442 10612 25452
rect 10892 25172 10948 25452
rect 11004 25414 11060 25452
rect 10536 25116 10800 25126
rect 10892 25116 11060 25172
rect 10592 25060 10640 25116
rect 10696 25060 10744 25116
rect 10536 25050 10800 25060
rect 10276 24052 10332 24062
rect 9884 24050 10332 24052
rect 9884 23998 10278 24050
rect 10330 23998 10332 24050
rect 9884 23996 10332 23998
rect 9884 23938 9940 23996
rect 9884 23886 9886 23938
rect 9938 23886 9940 23938
rect 9884 23874 9940 23886
rect 10220 23986 10332 23996
rect 9436 23314 9492 23324
rect 9212 23090 9268 23100
rect 9884 23156 9940 23166
rect 9884 23062 9940 23100
rect 8652 23044 8708 23054
rect 7980 22372 8036 22652
rect 8204 22932 8260 22942
rect 7980 22370 8148 22372
rect 7980 22318 7982 22370
rect 8034 22318 8148 22370
rect 7980 22316 8148 22318
rect 7980 22306 8036 22316
rect 7700 22260 7756 22270
rect 7700 22258 7924 22260
rect 7700 22206 7702 22258
rect 7754 22206 7924 22258
rect 7700 22204 7924 22206
rect 7700 22194 7756 22204
rect 7364 22148 7476 22158
rect 7420 22092 7476 22148
rect 7364 22054 7420 22092
rect 5964 21868 6748 21924
rect 5274 21812 5330 21822
rect 5274 21698 5330 21756
rect 5274 21646 5276 21698
rect 5328 21646 5330 21698
rect 5274 21634 5330 21646
rect 5964 21700 6020 21868
rect 6692 21810 6748 21868
rect 6692 21758 6694 21810
rect 6746 21758 6748 21810
rect 6692 21746 6748 21758
rect 6188 21700 6244 21710
rect 5964 21644 6076 21700
rect 6020 21642 6076 21644
rect 5516 21586 5572 21598
rect 5516 21534 5518 21586
rect 5570 21534 5572 21586
rect 6020 21590 6022 21642
rect 6074 21590 6076 21642
rect 6188 21606 6244 21644
rect 6524 21700 6580 21710
rect 6020 21578 6076 21590
rect 5516 21476 5572 21534
rect 5516 21028 5572 21420
rect 6524 21252 6580 21644
rect 7868 21364 7924 22204
rect 8092 21924 8148 22316
rect 8204 22370 8260 22876
rect 8204 22318 8206 22370
rect 8258 22318 8260 22370
rect 8204 22306 8260 22318
rect 8316 22370 8372 22382
rect 8316 22318 8318 22370
rect 8370 22318 8372 22370
rect 8316 22148 8372 22318
rect 8316 22082 8372 22092
rect 8092 21868 8428 21924
rect 8372 21476 8428 21868
rect 8372 21382 8428 21420
rect 7868 21308 8260 21364
rect 5874 21196 6138 21206
rect 6524 21196 6692 21252
rect 5930 21140 5978 21196
rect 6034 21140 6082 21196
rect 5874 21130 6138 21140
rect 5516 20962 5572 20972
rect 6468 21028 6524 21038
rect 2492 20738 2548 20748
rect 3836 20860 4900 20916
rect 2156 19954 2212 19964
rect 3836 20018 3892 20860
rect 4844 20804 4900 20860
rect 6468 20858 6524 20972
rect 4956 20804 5012 20814
rect 4844 20802 5012 20804
rect 4844 20750 4958 20802
rect 5010 20750 5012 20802
rect 4844 20748 5012 20750
rect 4956 20738 5012 20748
rect 5180 20804 5236 20814
rect 5722 20804 5778 20814
rect 5180 20802 5778 20804
rect 5180 20750 5182 20802
rect 5234 20750 5724 20802
rect 5776 20750 5778 20802
rect 5180 20748 5778 20750
rect 5180 20738 5236 20748
rect 5722 20738 5778 20748
rect 5964 20804 6020 20814
rect 6468 20806 6470 20858
rect 6522 20806 6524 20858
rect 6468 20794 6524 20806
rect 6636 20802 6692 21196
rect 5964 20710 6020 20748
rect 6636 20750 6638 20802
rect 6690 20750 6692 20802
rect 3836 19966 3838 20018
rect 3890 19966 3892 20018
rect 3836 19954 3892 19966
rect 4060 20692 4116 20702
rect 4060 20018 4116 20636
rect 4676 20690 4732 20702
rect 4676 20638 4678 20690
rect 4730 20638 4732 20690
rect 4676 20188 4732 20638
rect 6636 20580 6692 20750
rect 6636 20514 6692 20524
rect 6860 21028 6916 21038
rect 4620 20132 4732 20188
rect 4060 19966 4062 20018
rect 4114 19966 4116 20018
rect 4060 19954 4116 19966
rect 4172 20020 4228 20030
rect 3556 19796 3612 19806
rect 3276 19794 3612 19796
rect 3276 19742 3558 19794
rect 3610 19742 3612 19794
rect 3276 19740 3612 19742
rect 3276 19234 3332 19740
rect 3556 19730 3612 19740
rect 3276 19182 3278 19234
rect 3330 19182 3332 19234
rect 3276 19170 3332 19182
rect 4172 18900 4228 19964
rect 4620 19236 4676 20132
rect 6860 20130 6916 20972
rect 7308 21028 7364 21038
rect 7308 20802 7364 20972
rect 7308 20750 7310 20802
rect 7362 20750 7364 20802
rect 7308 20738 7364 20750
rect 7420 20804 7476 20814
rect 7066 20692 7122 20702
rect 7066 20598 7122 20636
rect 7196 20580 7252 20590
rect 7196 20188 7252 20524
rect 7420 20356 7476 20748
rect 7812 20804 7868 20814
rect 7812 20710 7868 20748
rect 8204 20802 8260 21308
rect 8204 20750 8206 20802
rect 8258 20750 8260 20802
rect 8204 20738 8260 20750
rect 7980 20690 8036 20702
rect 7980 20638 7982 20690
rect 8034 20638 8036 20690
rect 7980 20580 8036 20638
rect 7980 20514 8036 20524
rect 7420 20188 7476 20300
rect 8428 20244 8484 20254
rect 8652 20188 8708 22988
rect 9642 22932 9698 22942
rect 9642 22838 9698 22876
rect 9100 22370 9156 22382
rect 9100 22318 9102 22370
rect 9154 22318 9156 22370
rect 7196 20132 7364 20188
rect 7420 20132 7532 20188
rect 6860 20078 6862 20130
rect 6914 20078 6916 20130
rect 6860 20066 6916 20078
rect 7308 20130 7364 20132
rect 7308 20078 7310 20130
rect 7362 20078 7364 20130
rect 7308 20066 7364 20078
rect 7476 20074 7532 20132
rect 7476 20022 7478 20074
rect 7530 20022 7532 20074
rect 7476 20010 7532 20022
rect 7980 20018 8036 20030
rect 7980 19966 7982 20018
rect 8034 19966 8036 20018
rect 4956 19908 5012 19918
rect 4732 19906 5012 19908
rect 4732 19854 4958 19906
rect 5010 19854 5012 19906
rect 4732 19852 5012 19854
rect 4732 19458 4788 19852
rect 4956 19842 5012 19852
rect 5874 19628 6138 19638
rect 5930 19572 5978 19628
rect 6034 19572 6082 19628
rect 5874 19562 6138 19572
rect 4732 19406 4734 19458
rect 4786 19406 4788 19458
rect 4732 19394 4788 19406
rect 7980 19460 8036 19966
rect 8222 19796 8278 19806
rect 7980 19394 8036 19404
rect 8204 19794 8278 19796
rect 8204 19742 8224 19794
rect 8276 19742 8278 19794
rect 8204 19730 8278 19742
rect 4620 19170 4676 19180
rect 5516 19236 5572 19246
rect 5516 19142 5572 19180
rect 7980 19236 8036 19246
rect 6636 19010 6692 19022
rect 6636 18958 6638 19010
rect 6690 18958 6692 19010
rect 4172 18834 4228 18844
rect 5740 18900 5796 18910
rect 5740 18450 5796 18844
rect 5740 18398 5742 18450
rect 5794 18398 5796 18450
rect 5740 18386 5796 18398
rect 6524 18452 6580 18462
rect 6636 18452 6692 18958
rect 7812 19012 7868 19022
rect 7980 19012 8036 19180
rect 7812 19010 8036 19012
rect 7812 18958 7814 19010
rect 7866 18958 8036 19010
rect 7812 18956 8036 18958
rect 7812 18900 7868 18956
rect 7812 18834 7868 18844
rect 6524 18450 6692 18452
rect 6524 18398 6526 18450
rect 6578 18398 6692 18450
rect 6524 18396 6692 18398
rect 8204 18452 8260 19730
rect 8428 18562 8484 20188
rect 8428 18510 8430 18562
rect 8482 18510 8484 18562
rect 8428 18498 8484 18510
rect 8540 20132 8708 20188
rect 8876 21476 8932 21486
rect 6524 18386 6580 18396
rect 8204 18386 8260 18396
rect 8540 18116 8596 20132
rect 8876 19572 8932 21420
rect 9100 21028 9156 22318
rect 10220 22148 10276 23986
rect 10332 23828 10388 23838
rect 10332 23268 10388 23772
rect 10836 23716 10892 23726
rect 10836 23714 10948 23716
rect 10836 23662 10838 23714
rect 10890 23662 10948 23714
rect 10836 23650 10948 23662
rect 10892 23604 10948 23650
rect 10536 23548 10800 23558
rect 10592 23492 10640 23548
rect 10696 23492 10744 23548
rect 10536 23482 10800 23492
rect 10556 23268 10612 23278
rect 10332 23266 10612 23268
rect 10332 23214 10558 23266
rect 10610 23214 10612 23266
rect 10332 23212 10612 23214
rect 10556 23202 10612 23212
rect 10780 23268 10836 23278
rect 10780 23154 10836 23212
rect 10388 23098 10444 23110
rect 10388 23046 10390 23098
rect 10442 23046 10444 23098
rect 10388 23044 10444 23046
rect 10388 22978 10444 22988
rect 10780 23102 10782 23154
rect 10834 23102 10836 23154
rect 10780 22148 10836 23102
rect 9996 22092 10276 22148
rect 10332 22092 10836 22148
rect 10892 23044 10948 23548
rect 9324 21028 9380 21038
rect 9100 21026 9380 21028
rect 9100 20974 9326 21026
rect 9378 20974 9380 21026
rect 9100 20972 9380 20974
rect 9324 20962 9380 20972
rect 9436 20244 9492 20254
rect 9436 20018 9492 20188
rect 9604 20186 9660 20198
rect 9604 20134 9606 20186
rect 9658 20134 9660 20186
rect 9604 20132 9660 20134
rect 9604 20066 9660 20076
rect 9436 19966 9438 20018
rect 9490 19966 9492 20018
rect 9436 19954 9492 19966
rect 5874 18060 6138 18070
rect 5930 18004 5978 18060
rect 6034 18004 6082 18060
rect 8540 18050 8596 18060
rect 8652 19516 8932 19572
rect 5874 17994 6138 18004
rect 8540 17892 8596 17902
rect 8540 17798 8596 17836
rect 8652 16882 8708 19516
rect 8764 19234 8820 19246
rect 8764 19182 8766 19234
rect 8818 19182 8820 19234
rect 8764 17892 8820 19182
rect 9044 19012 9100 19022
rect 9044 18450 9100 18956
rect 9044 18398 9046 18450
rect 9098 18398 9100 18450
rect 9044 18386 9100 18398
rect 9436 18452 9492 18462
rect 9436 18358 9492 18396
rect 9660 18452 9716 18462
rect 9996 18452 10052 22092
rect 10220 21812 10276 21822
rect 9996 18396 10164 18452
rect 9660 18358 9716 18396
rect 9940 18228 9996 18238
rect 9660 18226 9996 18228
rect 9660 18174 9942 18226
rect 9994 18174 9996 18226
rect 9660 18172 9996 18174
rect 8764 17826 8820 17836
rect 8988 18116 9044 18126
rect 8652 16830 8654 16882
rect 8706 16830 8708 16882
rect 5874 16492 6138 16502
rect 5930 16436 5978 16492
rect 6034 16436 6082 16492
rect 5874 16426 6138 16436
rect 8652 16324 8708 16830
rect 8988 17108 9044 18060
rect 9660 17666 9716 18172
rect 9940 18162 9996 18172
rect 10108 18004 10164 18396
rect 9996 17948 10164 18004
rect 9660 17614 9662 17666
rect 9714 17614 9716 17666
rect 9660 17602 9716 17614
rect 9884 17892 9940 17902
rect 8988 16882 9044 17052
rect 9716 17108 9772 17118
rect 9716 17014 9772 17052
rect 8988 16830 8990 16882
rect 9042 16830 9044 16882
rect 8988 16818 9044 16830
rect 9884 16882 9940 17836
rect 9996 17666 10052 17948
rect 9996 17614 9998 17666
rect 10050 17614 10052 17666
rect 9996 17602 10052 17614
rect 9884 16830 9886 16882
rect 9938 16830 9940 16882
rect 9884 16818 9940 16830
rect 8652 16258 8708 16268
rect 5874 14924 6138 14934
rect 5930 14868 5978 14924
rect 6034 14868 6082 14924
rect 5874 14858 6138 14868
rect 10220 14756 10276 21756
rect 10332 16100 10388 22092
rect 10536 21980 10800 21990
rect 10592 21924 10640 21980
rect 10696 21924 10744 21980
rect 10536 21914 10800 21924
rect 10892 21812 10948 22988
rect 11004 23156 11060 25116
rect 11676 24612 11732 28364
rect 11788 27186 11844 28588
rect 11900 28420 11956 28430
rect 11900 27746 11956 28364
rect 12124 27972 12180 28812
rect 12460 28802 12516 28812
rect 12740 28868 12796 28878
rect 12740 28754 12796 28812
rect 12740 28702 12742 28754
rect 12794 28702 12796 28754
rect 12740 28690 12796 28702
rect 13020 28082 13076 29372
rect 13356 28196 13412 29372
rect 13356 28130 13412 28140
rect 13468 29426 13748 29428
rect 13468 29374 13694 29426
rect 13746 29374 13748 29426
rect 13468 29372 13748 29374
rect 13020 28030 13022 28082
rect 13074 28030 13076 28082
rect 13020 28018 13076 28030
rect 12124 27906 12180 27916
rect 11900 27694 11902 27746
rect 11954 27694 11956 27746
rect 11900 27682 11956 27694
rect 11788 27134 11790 27186
rect 11842 27134 11844 27186
rect 11788 27122 11844 27134
rect 12124 27188 12180 27198
rect 12124 27074 12180 27132
rect 12852 27188 12908 27198
rect 12852 27094 12908 27132
rect 13356 27188 13412 27198
rect 12124 27022 12126 27074
rect 12178 27022 12180 27074
rect 12124 27010 12180 27022
rect 11508 24556 11732 24612
rect 11788 26852 11844 26862
rect 11788 25508 11844 26796
rect 13356 26514 13412 27132
rect 13356 26462 13358 26514
rect 13410 26462 13412 26514
rect 12348 26317 12404 26329
rect 12348 26265 12350 26317
rect 12402 26265 12404 26317
rect 12348 26068 12404 26265
rect 12348 26002 12404 26012
rect 11788 25284 11844 25452
rect 12460 25508 12516 25518
rect 12460 25414 12516 25452
rect 11508 24052 11564 24556
rect 11452 24050 11564 24052
rect 11452 23998 11510 24050
rect 11562 23998 11564 24050
rect 11452 23986 11564 23998
rect 11004 22482 11060 23100
rect 11004 22430 11006 22482
rect 11058 22430 11060 22482
rect 11004 22418 11060 22430
rect 11116 23380 11172 23390
rect 11116 22372 11172 23324
rect 11452 23268 11508 23986
rect 11788 23716 11844 25228
rect 13076 25284 13132 25294
rect 13076 24946 13132 25228
rect 13076 24894 13078 24946
rect 13130 24894 13132 24946
rect 13076 24882 13132 24894
rect 12684 24724 12740 24734
rect 12460 24722 12740 24724
rect 12460 24670 12686 24722
rect 12738 24670 12740 24722
rect 12460 24668 12740 24670
rect 12348 24498 12404 24510
rect 12348 24446 12350 24498
rect 12402 24446 12404 24498
rect 12236 23940 12292 23950
rect 12236 23846 12292 23884
rect 11994 23828 12050 23838
rect 11994 23826 12180 23828
rect 11994 23774 11996 23826
rect 12048 23774 12180 23826
rect 11994 23772 12180 23774
rect 11994 23762 12050 23772
rect 11788 23650 11844 23660
rect 11452 23202 11508 23212
rect 11564 23380 11620 23390
rect 11564 23154 11620 23324
rect 11564 23102 11566 23154
rect 11618 23102 11620 23154
rect 11564 23090 11620 23102
rect 12012 23380 12068 23390
rect 11900 22372 11956 22382
rect 11116 22306 11172 22316
rect 11788 22316 11900 22372
rect 10892 21746 10948 21756
rect 11564 21586 11620 21598
rect 11564 21534 11566 21586
rect 11618 21534 11620 21586
rect 11284 21364 11340 21374
rect 11116 21362 11340 21364
rect 11116 21310 11286 21362
rect 11338 21310 11340 21362
rect 11116 21308 11340 21310
rect 11116 20802 11172 21308
rect 11284 21298 11340 21308
rect 11564 21028 11620 21534
rect 11788 21586 11844 22316
rect 11900 22278 11956 22316
rect 11788 21534 11790 21586
rect 11842 21534 11844 21586
rect 11788 21522 11844 21534
rect 11564 20962 11620 20972
rect 11116 20750 11118 20802
rect 11170 20750 11172 20802
rect 11116 20738 11172 20750
rect 10536 20412 10800 20422
rect 10592 20356 10640 20412
rect 10696 20356 10744 20412
rect 10536 20346 10800 20356
rect 12012 20018 12068 23324
rect 12124 22370 12180 23772
rect 12124 22318 12126 22370
rect 12178 22318 12180 22370
rect 12124 22306 12180 22318
rect 12236 23716 12292 23726
rect 12236 20916 12292 23660
rect 12348 23154 12404 24446
rect 12348 23102 12350 23154
rect 12402 23102 12404 23154
rect 12348 23090 12404 23102
rect 12460 22606 12516 24668
rect 12684 24658 12740 24668
rect 12908 24724 12964 24734
rect 12740 24164 12796 24174
rect 12740 23994 12796 24108
rect 12740 23942 12742 23994
rect 12794 23942 12796 23994
rect 12740 23930 12796 23942
rect 12908 23938 12964 24668
rect 12908 23886 12910 23938
rect 12962 23886 12964 23938
rect 12908 23380 12964 23886
rect 12404 22594 12516 22606
rect 12404 22542 12406 22594
rect 12458 22542 12516 22594
rect 12404 22540 12516 22542
rect 12572 23324 12964 23380
rect 13356 23380 13412 26462
rect 12404 22530 12460 22540
rect 12572 21700 12628 23324
rect 13356 23314 13412 23324
rect 12684 21700 12740 21710
rect 12572 21698 12740 21700
rect 12572 21646 12686 21698
rect 12738 21646 12740 21698
rect 12572 21644 12740 21646
rect 12684 21634 12740 21644
rect 13468 21140 13524 29372
rect 13692 29362 13748 29372
rect 13636 28868 13692 28878
rect 13636 28754 13692 28812
rect 13636 28702 13638 28754
rect 13690 28702 13692 28754
rect 13636 28690 13692 28702
rect 14140 27858 14196 27870
rect 14140 27806 14142 27858
rect 14194 27806 14196 27858
rect 14010 27300 14066 27310
rect 14010 27206 14066 27244
rect 13636 27188 13692 27198
rect 13636 27094 13692 27132
rect 13804 26964 13860 26974
rect 13804 25730 13860 26908
rect 13804 25678 13806 25730
rect 13858 25678 13860 25730
rect 13804 25666 13860 25678
rect 14140 25508 14196 27806
rect 14140 25442 14196 25452
rect 14252 27074 14308 27086
rect 14252 27022 14254 27074
rect 14306 27022 14308 27074
rect 14252 24724 14308 27022
rect 14364 24946 14420 29708
rect 14532 30210 14756 30212
rect 14532 30158 14702 30210
rect 14754 30158 14756 30210
rect 14532 30156 14756 30158
rect 14532 29652 14588 30156
rect 14700 30146 14756 30156
rect 14476 29650 14588 29652
rect 14476 29598 14534 29650
rect 14586 29598 14588 29650
rect 14476 29586 14588 29598
rect 14812 30100 14868 30110
rect 15148 30100 15204 30380
rect 14476 27636 14532 29586
rect 14476 27570 14532 27580
rect 14588 28196 14644 28206
rect 14364 24894 14366 24946
rect 14418 24894 14420 24946
rect 14364 24882 14420 24894
rect 13804 24668 14308 24724
rect 13636 24500 13692 24510
rect 13636 23994 13692 24444
rect 13636 23942 13638 23994
rect 13690 23942 13692 23994
rect 13636 23940 13692 23942
rect 13636 23864 13692 23884
rect 13580 23770 13636 23782
rect 13580 23718 13582 23770
rect 13634 23718 13636 23770
rect 13580 23716 13636 23718
rect 13580 23650 13636 23660
rect 13804 21924 13860 24668
rect 14252 24500 14308 24510
rect 12236 20850 12292 20860
rect 13356 21084 13524 21140
rect 13692 21868 13860 21924
rect 13916 24164 13972 24174
rect 13692 21140 13748 21868
rect 13804 21700 13860 21710
rect 13804 21586 13860 21644
rect 13804 21534 13806 21586
rect 13858 21534 13860 21586
rect 13804 21522 13860 21534
rect 13356 20804 13412 21084
rect 13692 21074 13748 21084
rect 13562 21028 13618 21038
rect 13562 20934 13618 20972
rect 13356 20738 13412 20748
rect 13804 20804 13860 20814
rect 13916 20804 13972 24108
rect 14140 24052 14196 24062
rect 14140 23938 14196 23996
rect 14140 23886 14142 23938
rect 14194 23886 14196 23938
rect 14140 23874 14196 23886
rect 14252 23266 14308 24444
rect 14588 23940 14644 28140
rect 14812 28082 14868 30044
rect 15036 30044 15204 30100
rect 14812 28030 14814 28082
rect 14866 28030 14868 28082
rect 14812 28018 14868 28030
rect 14924 29594 14980 29606
rect 14924 29542 14926 29594
rect 14978 29542 14980 29594
rect 14924 27412 14980 29542
rect 15036 29426 15092 30044
rect 15036 29374 15038 29426
rect 15090 29374 15092 29426
rect 15260 29482 15316 30380
rect 15932 30436 15988 31726
rect 16156 31108 16212 31892
rect 16380 31892 16436 32398
rect 16492 32340 16548 32525
rect 16716 32676 16772 32686
rect 16716 32562 16772 32620
rect 16716 32510 16718 32562
rect 16770 32510 16772 32562
rect 16716 32498 16772 32510
rect 16828 32340 16884 33516
rect 16492 32274 16548 32284
rect 16716 32284 16884 32340
rect 16380 31826 16436 31836
rect 16716 31890 16772 32284
rect 16716 31838 16718 31890
rect 16770 31838 16772 31890
rect 16716 31826 16772 31838
rect 16268 31778 16324 31790
rect 16268 31726 16270 31778
rect 16322 31726 16324 31778
rect 17276 31778 17332 34636
rect 17948 34298 18004 35308
rect 17948 34246 17950 34298
rect 18002 34246 18004 34298
rect 17948 34234 18004 34246
rect 17836 34169 17892 34181
rect 17612 34130 17668 34142
rect 17612 34078 17614 34130
rect 17666 34078 17668 34130
rect 17500 33236 17556 33246
rect 17500 32674 17556 33180
rect 17500 32622 17502 32674
rect 17554 32622 17556 32674
rect 17500 32116 17556 32622
rect 17612 32452 17668 34078
rect 17836 34117 17838 34169
rect 17890 34117 17892 34169
rect 17836 33572 17892 34117
rect 18172 34130 18228 34142
rect 18172 34078 18174 34130
rect 18226 34078 18228 34130
rect 17836 33506 17892 33516
rect 17948 33908 18004 33918
rect 17948 33318 18004 33852
rect 17948 33266 17950 33318
rect 18002 33266 18004 33318
rect 17948 33254 18004 33266
rect 18172 33124 18228 34078
rect 18284 33684 18340 39228
rect 18816 39200 18928 40000
rect 19936 39200 20048 40000
rect 21056 39200 21168 40000
rect 22176 39200 22288 40000
rect 23296 39200 23408 40000
rect 24416 39200 24528 40000
rect 25536 39200 25648 40000
rect 26656 39200 26768 40000
rect 27776 39200 27888 40000
rect 28896 39200 29008 40000
rect 30016 39200 30128 40000
rect 31136 39200 31248 40000
rect 32256 39200 32368 40000
rect 33376 39200 33488 40000
rect 34496 39200 34608 40000
rect 35616 39200 35728 40000
rect 36736 39200 36848 40000
rect 18844 36484 18900 39200
rect 19180 36708 19236 36718
rect 19180 36614 19236 36652
rect 19964 36708 20020 39200
rect 19964 36642 20020 36652
rect 18844 36428 19236 36484
rect 18620 34804 18676 34814
rect 18620 34710 18676 34748
rect 19068 34804 19124 34814
rect 18788 34692 18844 34702
rect 18788 34354 18844 34636
rect 18788 34302 18790 34354
rect 18842 34302 18844 34354
rect 18788 34290 18844 34302
rect 19068 34157 19124 34748
rect 19180 34356 19236 36428
rect 19852 36454 19908 36466
rect 19852 36402 19854 36454
rect 19906 36402 19908 36454
rect 19852 36260 19908 36402
rect 19740 36204 19908 36260
rect 20860 36370 20916 36382
rect 20860 36318 20862 36370
rect 20914 36318 20916 36370
rect 19740 35588 19796 36204
rect 19860 36092 20124 36102
rect 19916 36036 19964 36092
rect 20020 36036 20068 36092
rect 19860 36026 20124 36036
rect 20300 35924 20356 35934
rect 19964 35588 20020 35598
rect 19740 35586 20132 35588
rect 19740 35534 19966 35586
rect 20018 35534 20132 35586
rect 19740 35532 20132 35534
rect 19964 35522 20020 35532
rect 19964 35028 20020 35038
rect 19740 35026 20020 35028
rect 19740 34974 19966 35026
rect 20018 34974 20020 35026
rect 19740 34972 20020 34974
rect 19628 34916 19684 34926
rect 19628 34822 19684 34860
rect 19180 34290 19236 34300
rect 19068 34105 19070 34157
rect 19122 34105 19124 34157
rect 19068 34093 19124 34105
rect 18284 33618 18340 33628
rect 18396 33796 18452 33806
rect 19740 33796 19796 34972
rect 19964 34962 20020 34972
rect 20076 34916 20132 35532
rect 19964 34858 20020 34870
rect 19964 34806 19966 34858
rect 20018 34806 20020 34858
rect 20076 34850 20132 34860
rect 20300 34916 20356 35868
rect 20860 35700 20916 36318
rect 20972 35924 21028 35934
rect 20972 35810 21028 35868
rect 20972 35758 20974 35810
rect 21026 35758 21028 35810
rect 20972 35746 21028 35758
rect 20580 35588 20636 35598
rect 20580 35494 20636 35532
rect 20860 35364 20916 35644
rect 20860 35308 21028 35364
rect 20804 35140 20860 35150
rect 20804 35026 20860 35084
rect 20804 34974 20806 35026
rect 20858 34974 20860 35026
rect 20804 34962 20860 34974
rect 20300 34914 20692 34916
rect 20300 34862 20302 34914
rect 20354 34862 20692 34914
rect 20300 34860 20692 34862
rect 20300 34850 20356 34860
rect 19964 34692 20020 34806
rect 19964 34636 20244 34692
rect 19860 34524 20124 34534
rect 19916 34468 19964 34524
rect 20020 34468 20068 34524
rect 19860 34458 20124 34468
rect 20188 34356 20244 34636
rect 18172 33058 18228 33068
rect 18396 32788 18452 33740
rect 18284 32732 18452 32788
rect 18732 33740 19796 33796
rect 20076 34300 20244 34356
rect 20412 34356 20468 34366
rect 18060 32676 18116 32686
rect 17612 32386 17668 32396
rect 17836 32562 17892 32574
rect 17836 32510 17838 32562
rect 17890 32510 17892 32562
rect 17500 32050 17556 32060
rect 17836 32004 17892 32510
rect 18060 32562 18116 32620
rect 18060 32510 18062 32562
rect 18114 32510 18116 32562
rect 18060 32498 18116 32510
rect 17836 31938 17892 31948
rect 16268 31332 16324 31726
rect 16604 31734 16660 31746
rect 16604 31682 16606 31734
rect 16658 31682 16660 31734
rect 16268 31276 16436 31332
rect 16268 31108 16324 31118
rect 16156 31106 16324 31108
rect 16156 31054 16270 31106
rect 16322 31054 16324 31106
rect 16156 31052 16324 31054
rect 16268 31042 16324 31052
rect 16044 30996 16100 31006
rect 16380 30996 16436 31276
rect 16044 30994 16212 30996
rect 16044 30942 16046 30994
rect 16098 30942 16212 30994
rect 16044 30940 16212 30942
rect 16380 30940 16492 30996
rect 16044 30930 16100 30940
rect 15932 30370 15988 30380
rect 15484 30212 15596 30222
rect 16044 30212 16100 30222
rect 15540 30210 15596 30212
rect 15540 30158 15542 30210
rect 15594 30158 15596 30210
rect 15540 30156 15596 30158
rect 15484 30146 15596 30156
rect 15708 30210 16100 30212
rect 15708 30158 16046 30210
rect 16098 30158 16100 30210
rect 15708 30156 16100 30158
rect 15372 30098 15428 30110
rect 15372 30046 15374 30098
rect 15426 30046 15428 30098
rect 15372 29876 15428 30046
rect 15372 29810 15428 29820
rect 15596 29876 15652 29886
rect 15260 29430 15262 29482
rect 15314 29430 15316 29482
rect 15260 29418 15316 29430
rect 15596 29426 15652 29820
rect 15036 29362 15092 29374
rect 15596 29374 15598 29426
rect 15650 29374 15652 29426
rect 15596 29362 15652 29374
rect 15198 29036 15462 29046
rect 15254 28980 15302 29036
rect 15358 28980 15406 29036
rect 15198 28970 15462 28980
rect 15708 28532 15764 30156
rect 16044 30146 16100 30156
rect 16156 29988 16212 30940
rect 16436 30938 16492 30940
rect 16436 30886 16438 30938
rect 16490 30886 16492 30938
rect 16286 30660 16342 30670
rect 16286 30210 16342 30604
rect 16436 30436 16492 30886
rect 16436 30380 16548 30436
rect 16286 30158 16288 30210
rect 16340 30158 16342 30210
rect 16286 30146 16342 30158
rect 16492 30100 16548 30380
rect 16604 30324 16660 31682
rect 17276 31726 17278 31778
rect 17330 31726 17332 31778
rect 16940 31220 16996 31230
rect 16940 30996 16996 31164
rect 16940 30902 16996 30940
rect 16772 30770 16828 30782
rect 16772 30718 16774 30770
rect 16826 30718 16828 30770
rect 16772 30436 16828 30718
rect 16772 30370 16828 30380
rect 16604 30258 16660 30268
rect 17108 30324 17164 30334
rect 17276 30324 17332 31726
rect 17500 31892 17556 31902
rect 17500 30994 17556 31836
rect 18060 31778 18116 31790
rect 18060 31726 18062 31778
rect 18114 31726 18116 31778
rect 17500 30942 17502 30994
rect 17554 30942 17556 30994
rect 17500 30930 17556 30942
rect 17836 31220 17892 31230
rect 17836 30994 17892 31164
rect 17836 30942 17838 30994
rect 17890 30942 17892 30994
rect 17836 30930 17892 30942
rect 17108 30322 17332 30324
rect 17108 30270 17110 30322
rect 17162 30270 17332 30322
rect 17108 30268 17332 30270
rect 17108 30258 17164 30268
rect 16940 30212 16996 30222
rect 16492 30044 16772 30100
rect 16156 29922 16212 29932
rect 16268 29876 16324 29886
rect 16268 29204 16324 29820
rect 16268 29148 16380 29204
rect 15596 28476 15764 28532
rect 15820 28868 15876 28878
rect 15148 27860 15204 27870
rect 14756 27356 14980 27412
rect 15036 27858 15204 27860
rect 15036 27806 15150 27858
rect 15202 27806 15204 27858
rect 15036 27804 15204 27806
rect 14756 27130 14812 27356
rect 14756 27078 14758 27130
rect 14810 27078 14812 27130
rect 14756 27066 14812 27078
rect 14924 26964 14980 27002
rect 15036 26964 15092 27804
rect 15148 27794 15204 27804
rect 15198 27468 15462 27478
rect 15254 27412 15302 27468
rect 15358 27412 15406 27468
rect 15198 27402 15462 27412
rect 15260 27076 15316 27086
rect 15260 26982 15316 27020
rect 15428 27076 15484 27086
rect 15428 26982 15484 27020
rect 14980 26908 15092 26964
rect 14924 26898 14980 26908
rect 14980 26178 15036 26190
rect 14980 26126 14982 26178
rect 15034 26126 15036 26178
rect 14980 26068 15036 26126
rect 14980 26002 15036 26012
rect 15198 25900 15462 25910
rect 15254 25844 15302 25900
rect 15358 25844 15406 25900
rect 15198 25834 15462 25844
rect 15596 25732 15652 28476
rect 15820 27076 15876 28812
rect 16324 28698 16380 29148
rect 16156 28642 16212 28654
rect 16156 28590 16158 28642
rect 16210 28590 16212 28642
rect 16324 28646 16326 28698
rect 16378 28646 16380 28698
rect 16324 28634 16380 28646
rect 16604 28644 16660 28654
rect 16156 28196 16212 28590
rect 16604 28550 16660 28588
rect 16492 28530 16548 28542
rect 16492 28478 16494 28530
rect 16546 28478 16548 28530
rect 16492 28420 16548 28478
rect 16716 28420 16772 30044
rect 16940 28878 16996 30156
rect 16884 28866 16996 28878
rect 16884 28814 16886 28866
rect 16938 28814 16996 28866
rect 16884 28812 16996 28814
rect 16884 28802 16940 28812
rect 17164 28532 17220 28542
rect 16492 28354 16548 28364
rect 16604 28364 16772 28420
rect 17052 28420 17108 28430
rect 16156 28140 16492 28196
rect 16436 27970 16492 28140
rect 16436 27918 16438 27970
rect 16490 27918 16492 27970
rect 16436 27906 16492 27918
rect 16604 27860 16660 28364
rect 16604 27794 16660 27804
rect 16716 27858 16772 27870
rect 16716 27806 16718 27858
rect 16770 27806 16772 27858
rect 16604 27412 16660 27422
rect 15820 27010 15876 27020
rect 15932 27074 15988 27086
rect 15932 27022 15934 27074
rect 15986 27022 15988 27074
rect 15932 26908 15988 27022
rect 16174 27076 16230 27086
rect 16174 26982 16230 27020
rect 15372 25676 15652 25732
rect 15708 26852 15988 26908
rect 15260 25508 15316 25518
rect 15260 25414 15316 25452
rect 15372 25284 15428 25676
rect 15204 25228 15428 25284
rect 15484 25506 15540 25518
rect 15484 25454 15486 25506
rect 15538 25454 15540 25506
rect 14700 24948 14756 24958
rect 14700 24946 14868 24948
rect 14700 24894 14702 24946
rect 14754 24894 14868 24946
rect 14700 24892 14868 24894
rect 14700 24882 14756 24892
rect 14700 23940 14756 23950
rect 14588 23938 14756 23940
rect 14588 23886 14702 23938
rect 14754 23886 14756 23938
rect 14588 23884 14756 23886
rect 14700 23874 14756 23884
rect 14382 23828 14438 23838
rect 14382 23826 14644 23828
rect 14382 23774 14384 23826
rect 14436 23774 14644 23826
rect 14382 23772 14644 23774
rect 14382 23762 14438 23772
rect 14252 23214 14254 23266
rect 14306 23214 14308 23266
rect 14252 23202 14308 23214
rect 14588 23154 14644 23772
rect 14812 23716 14868 24892
rect 15204 24946 15260 25228
rect 15204 24894 15206 24946
rect 15258 24894 15260 24946
rect 15204 24882 15260 24894
rect 15036 24722 15092 24734
rect 15036 24670 15038 24722
rect 15090 24670 15092 24722
rect 15036 24164 15092 24670
rect 15484 24500 15540 25454
rect 15484 24434 15540 24444
rect 15198 24332 15462 24342
rect 15254 24276 15302 24332
rect 15358 24276 15406 24332
rect 15198 24266 15462 24276
rect 15036 24098 15092 24108
rect 15036 23716 15092 23726
rect 14812 23714 15092 23716
rect 14812 23662 15038 23714
rect 15090 23662 15092 23714
rect 14812 23660 15092 23662
rect 14588 23102 14590 23154
rect 14642 23102 14644 23154
rect 14588 23090 14644 23102
rect 14812 23154 14868 23166
rect 14812 23102 14814 23154
rect 14866 23102 14868 23154
rect 14812 23044 14868 23102
rect 14028 22932 14084 22942
rect 14028 22370 14084 22876
rect 14812 22708 14868 22988
rect 14812 22642 14868 22652
rect 14028 22318 14030 22370
rect 14082 22318 14084 22370
rect 14028 22306 14084 22318
rect 14924 22148 14980 23660
rect 15036 23650 15092 23660
rect 15708 23604 15764 26852
rect 16604 26516 16660 27356
rect 16716 27300 16772 27806
rect 16716 27234 16772 27244
rect 16828 27858 16884 27870
rect 16828 27806 16830 27858
rect 16882 27806 16884 27858
rect 16716 26516 16772 26526
rect 16604 26514 16772 26516
rect 16604 26462 16718 26514
rect 16770 26462 16772 26514
rect 16604 26460 16772 26462
rect 16716 26450 16772 26460
rect 15820 26404 15876 26414
rect 15820 25620 15876 26348
rect 16828 26404 16884 27806
rect 16828 26338 16884 26348
rect 16380 26292 16436 26302
rect 15932 26180 15988 26190
rect 15932 25674 15988 26124
rect 15932 25622 15934 25674
rect 15986 25622 15988 25674
rect 15932 25610 15988 25622
rect 15820 25506 15876 25564
rect 15820 25454 15822 25506
rect 15874 25454 15876 25506
rect 15820 25442 15876 25454
rect 16380 25508 16436 26236
rect 16380 25442 16436 25452
rect 16716 23938 16772 23950
rect 16716 23886 16718 23938
rect 16770 23886 16772 23938
rect 15708 23548 15876 23604
rect 15652 23380 15708 23390
rect 15652 23286 15708 23324
rect 15092 22932 15148 22970
rect 15092 22866 15148 22876
rect 15198 22764 15462 22774
rect 15254 22708 15302 22764
rect 15358 22708 15406 22764
rect 15198 22698 15462 22708
rect 15484 22372 15540 22382
rect 15484 22278 15540 22316
rect 13804 20802 13916 20804
rect 13804 20750 13806 20802
rect 13858 20750 13916 20802
rect 13804 20748 13916 20750
rect 13804 20738 13860 20748
rect 13916 20710 13972 20748
rect 14028 22092 14980 22148
rect 12572 20578 12628 20590
rect 12572 20526 12574 20578
rect 12626 20526 12628 20578
rect 12572 20188 12628 20526
rect 14028 20188 14084 22092
rect 15820 22036 15876 23548
rect 15596 21980 15876 22036
rect 15932 23380 15988 23390
rect 15932 22372 15988 23324
rect 16604 23380 16660 23390
rect 16100 23044 16156 23054
rect 16100 22950 16156 22988
rect 16044 22372 16100 22382
rect 15932 22370 16100 22372
rect 15932 22318 16046 22370
rect 16098 22318 16100 22370
rect 15932 22316 16100 22318
rect 14812 21924 14868 21934
rect 14476 21700 14532 21710
rect 14476 21586 14532 21644
rect 14476 21534 14478 21586
rect 14530 21534 14532 21586
rect 14476 21522 14532 21534
rect 12572 20132 12852 20188
rect 12012 19966 12014 20018
rect 12066 19966 12068 20018
rect 12012 19954 12068 19966
rect 12796 20018 12852 20132
rect 12796 19966 12798 20018
rect 12850 19966 12852 20018
rect 12796 19954 12852 19966
rect 13916 20132 14084 20188
rect 14140 21364 14196 21374
rect 14140 21362 14532 21364
rect 14140 21310 14142 21362
rect 14194 21310 14532 21362
rect 14140 21308 14532 21310
rect 10668 19908 10724 19918
rect 10668 19460 10724 19852
rect 10668 19346 10724 19404
rect 12236 19908 12292 19918
rect 10668 19294 10670 19346
rect 10722 19294 10724 19346
rect 10668 19282 10724 19294
rect 11900 19348 11956 19358
rect 11900 19234 11956 19292
rect 11900 19182 11902 19234
rect 11954 19182 11956 19234
rect 11900 19170 11956 19182
rect 12068 19180 12124 19190
rect 12068 19178 12180 19180
rect 12068 19126 12070 19178
rect 12122 19126 12180 19178
rect 12068 19114 12180 19126
rect 11284 19012 11340 19022
rect 11284 18918 11340 18956
rect 10536 18844 10800 18854
rect 10592 18788 10640 18844
rect 10696 18788 10744 18844
rect 10536 18778 10800 18788
rect 10892 18452 10948 18462
rect 10724 18226 10780 18238
rect 10724 18174 10726 18226
rect 10778 18174 10780 18226
rect 10724 17892 10780 18174
rect 10724 17826 10780 17836
rect 10892 17780 10948 18396
rect 11004 18450 11060 18462
rect 11004 18398 11006 18450
rect 11058 18398 11060 18450
rect 11004 18228 11060 18398
rect 11116 18452 11172 18462
rect 11116 18358 11172 18396
rect 11788 18452 11844 18462
rect 11788 18450 11956 18452
rect 11788 18398 11790 18450
rect 11842 18398 11956 18450
rect 11788 18396 11956 18398
rect 11788 18386 11844 18396
rect 11546 18228 11602 18238
rect 11004 18226 11602 18228
rect 11004 18174 11548 18226
rect 11600 18174 11602 18226
rect 11004 18172 11602 18174
rect 11546 18162 11602 18172
rect 11900 17780 11956 18396
rect 10892 17724 11060 17780
rect 10780 17668 10836 17678
rect 10780 17666 10948 17668
rect 10780 17614 10782 17666
rect 10834 17614 10948 17666
rect 10780 17612 10948 17614
rect 10780 17602 10836 17612
rect 10536 17276 10800 17286
rect 10592 17220 10640 17276
rect 10696 17220 10744 17276
rect 10536 17210 10800 17220
rect 10892 17108 10948 17612
rect 11004 17332 11060 17724
rect 11900 17714 11956 17724
rect 11004 17276 11172 17332
rect 11004 17108 11060 17118
rect 10892 17106 11060 17108
rect 10892 17054 11006 17106
rect 11058 17054 11060 17106
rect 10892 17052 11060 17054
rect 11004 17042 11060 17052
rect 10332 16034 10388 16044
rect 10892 16100 10948 16110
rect 10536 15708 10800 15718
rect 10592 15652 10640 15708
rect 10696 15652 10744 15708
rect 10536 15642 10800 15652
rect 10220 14690 10276 14700
rect 7084 14530 7140 14542
rect 7084 14478 7086 14530
rect 7138 14478 7140 14530
rect 5874 13356 6138 13366
rect 5930 13300 5978 13356
rect 6034 13300 6082 13356
rect 5874 13290 6138 13300
rect 5874 11788 6138 11798
rect 5930 11732 5978 11788
rect 6034 11732 6082 11788
rect 5874 11722 6138 11732
rect 7084 11732 7140 14478
rect 7868 14530 7924 14542
rect 7868 14478 7870 14530
rect 7922 14478 7924 14530
rect 7868 13972 7924 14478
rect 10892 14530 10948 16044
rect 11004 15988 11060 15998
rect 11116 15988 11172 17276
rect 12124 16996 12180 19114
rect 12236 19124 12292 19852
rect 13916 19796 13972 20132
rect 14140 20055 14196 21308
rect 14476 20802 14532 21308
rect 14308 20746 14364 20758
rect 14308 20694 14310 20746
rect 14362 20694 14364 20746
rect 14476 20750 14478 20802
rect 14530 20750 14532 20802
rect 14476 20738 14532 20750
rect 14700 20804 14756 20814
rect 14308 20188 14364 20694
rect 12572 19684 12628 19694
rect 12460 19348 12516 19358
rect 12236 19068 12348 19124
rect 12292 18506 12348 19068
rect 12292 18454 12294 18506
rect 12346 18454 12348 18506
rect 12292 18442 12348 18454
rect 12460 18562 12516 19292
rect 12572 19234 12628 19628
rect 12572 19182 12574 19234
rect 12626 19182 12628 19234
rect 13412 19460 13468 19470
rect 13412 19290 13468 19404
rect 13916 19460 13972 19740
rect 13916 19394 13972 19404
rect 14028 19999 14196 20055
rect 14252 20132 14364 20188
rect 13412 19238 13414 19290
rect 13466 19238 13468 19290
rect 14028 19348 14084 19999
rect 14028 19282 14084 19292
rect 14252 19684 14308 20132
rect 14700 20130 14756 20748
rect 14700 20078 14702 20130
rect 14754 20078 14756 20130
rect 14700 20066 14756 20078
rect 14252 19348 14308 19628
rect 14252 19282 14308 19292
rect 14364 20020 14420 20030
rect 13412 19226 13468 19238
rect 13692 19236 13748 19246
rect 12572 19170 12628 19182
rect 12814 19124 12870 19134
rect 13580 19124 13636 19134
rect 12814 19122 13188 19124
rect 12814 19070 12816 19122
rect 12868 19070 13188 19122
rect 12814 19068 13188 19070
rect 12814 19058 12870 19068
rect 12460 18510 12462 18562
rect 12514 18510 12516 18562
rect 12460 18228 12516 18510
rect 12908 18452 12964 18462
rect 12908 18358 12964 18396
rect 13132 18450 13188 19068
rect 13580 19030 13636 19068
rect 13132 18398 13134 18450
rect 13186 18398 13188 18450
rect 13132 18386 13188 18398
rect 13244 18452 13300 18462
rect 12124 16930 12180 16940
rect 12348 18172 12516 18228
rect 12348 16994 12404 18172
rect 12684 17780 12740 17790
rect 12572 17724 12684 17780
rect 12572 17556 12628 17724
rect 12684 17686 12740 17724
rect 13244 17668 13300 18396
rect 13412 18452 13468 18462
rect 13412 18358 13468 18396
rect 13356 17668 13412 17678
rect 13580 17668 13636 17678
rect 13244 17666 13412 17668
rect 13244 17614 13358 17666
rect 13410 17614 13412 17666
rect 13244 17612 13412 17614
rect 13356 17602 13412 17612
rect 13468 17666 13636 17668
rect 13468 17614 13582 17666
rect 13634 17614 13636 17666
rect 13468 17612 13636 17614
rect 12348 16942 12350 16994
rect 12402 16942 12404 16994
rect 12348 16930 12404 16942
rect 12516 17500 12628 17556
rect 12516 16938 12572 17500
rect 13468 17108 13524 17612
rect 13580 17602 13636 17612
rect 13262 17052 13524 17108
rect 13580 17108 13636 17118
rect 12516 16886 12518 16938
rect 12570 16886 12572 16938
rect 12516 16874 12572 16886
rect 13020 16996 13076 17006
rect 13020 16882 13076 16940
rect 13262 16994 13318 17052
rect 13262 16942 13264 16994
rect 13316 16942 13318 16994
rect 13262 16930 13318 16942
rect 13580 16884 13636 17052
rect 13020 16830 13022 16882
rect 13074 16830 13076 16882
rect 13020 16818 13076 16830
rect 13356 16828 13636 16884
rect 13692 16882 13748 19180
rect 13804 19234 13860 19246
rect 13804 19182 13806 19234
rect 13858 19182 13860 19234
rect 13804 18788 13860 19182
rect 14140 19196 14196 19208
rect 14140 19144 14142 19196
rect 14194 19180 14196 19196
rect 14364 19180 14420 19964
rect 14194 19144 14420 19180
rect 13804 18722 13860 18732
rect 14028 19124 14084 19134
rect 14140 19124 14420 19144
rect 14476 19236 14532 19246
rect 14476 19142 14532 19180
rect 13804 18452 13860 18462
rect 13804 18358 13860 18396
rect 13860 17554 13916 17566
rect 13860 17502 13862 17554
rect 13914 17502 13916 17554
rect 13860 17108 13916 17502
rect 13860 17042 13916 17052
rect 13692 16830 13694 16882
rect 13746 16830 13748 16882
rect 11340 16100 11396 16110
rect 11732 16100 11788 16110
rect 11396 16098 12180 16100
rect 11396 16046 11734 16098
rect 11786 16046 12180 16098
rect 11396 16044 12180 16046
rect 11340 16006 11396 16044
rect 11732 16034 11788 16044
rect 11004 15986 11172 15988
rect 11004 15934 11006 15986
rect 11058 15934 11172 15986
rect 11004 15932 11172 15934
rect 11004 15922 11060 15932
rect 12124 15538 12180 16044
rect 13356 16098 13412 16828
rect 13356 16046 13358 16098
rect 13410 16046 13412 16098
rect 13356 16034 13412 16046
rect 12124 15486 12126 15538
rect 12178 15486 12180 15538
rect 11508 14756 11564 14766
rect 11116 14754 11564 14756
rect 11116 14702 11510 14754
rect 11562 14702 11564 14754
rect 11116 14700 11564 14702
rect 10892 14478 10894 14530
rect 10946 14478 10948 14530
rect 10892 14466 10948 14478
rect 11004 14530 11060 14542
rect 11004 14478 11006 14530
rect 11058 14478 11060 14530
rect 9772 14418 9828 14430
rect 9772 14366 9774 14418
rect 9826 14366 9828 14418
rect 7980 13972 8036 13982
rect 7868 13970 8036 13972
rect 7868 13918 7982 13970
rect 8034 13918 8036 13970
rect 7868 13916 8036 13918
rect 7980 13906 8036 13916
rect 9100 13748 9156 13758
rect 8596 13746 9156 13748
rect 8596 13694 9102 13746
rect 9154 13694 9156 13746
rect 8596 13692 9156 13694
rect 9772 13748 9828 14366
rect 10556 14308 10612 14318
rect 11004 14308 11060 14478
rect 10332 14306 11060 14308
rect 10332 14254 10558 14306
rect 10610 14254 11060 14306
rect 10332 14252 11060 14254
rect 9996 13748 10052 13758
rect 9772 13746 10052 13748
rect 9772 13694 9998 13746
rect 10050 13694 10052 13746
rect 9772 13692 10052 13694
rect 8596 13186 8652 13692
rect 9100 13682 9156 13692
rect 9754 13524 9810 13534
rect 8596 13134 8598 13186
rect 8650 13134 8652 13186
rect 8596 13122 8652 13134
rect 8876 13522 9810 13524
rect 8876 13470 9756 13522
rect 9808 13470 9810 13522
rect 8876 13468 9810 13470
rect 8876 12962 8932 13468
rect 9754 13458 9810 13468
rect 9212 13300 9268 13310
rect 8876 12910 8878 12962
rect 8930 12910 8932 12962
rect 8876 12898 8932 12910
rect 9100 12964 9156 12974
rect 9212 12964 9268 13244
rect 9100 12962 9268 12964
rect 9100 12910 9102 12962
rect 9154 12910 9268 12962
rect 9100 12908 9268 12910
rect 9100 12898 9156 12908
rect 7812 12740 7868 12750
rect 7644 12738 7868 12740
rect 7644 12686 7814 12738
rect 7866 12686 7868 12738
rect 7644 12684 7868 12686
rect 7308 12404 7364 12414
rect 7308 12310 7364 12348
rect 7644 12292 7700 12684
rect 7812 12674 7868 12684
rect 7644 12178 7700 12236
rect 8652 12404 8708 12414
rect 7644 12126 7646 12178
rect 7698 12126 7700 12178
rect 7644 12114 7700 12126
rect 7868 12178 7924 12190
rect 7868 12126 7870 12178
rect 7922 12126 7924 12178
rect 7084 11666 7140 11676
rect 7868 12068 7924 12126
rect 8036 12180 8092 12190
rect 8036 12086 8092 12124
rect 8540 12178 8596 12190
rect 8540 12126 8542 12178
rect 8594 12126 8596 12178
rect 5852 11620 5908 11630
rect 5852 11396 5908 11564
rect 6636 11396 6692 11406
rect 5516 11394 5908 11396
rect 5516 11342 5854 11394
rect 5906 11342 5908 11394
rect 5516 11340 5908 11342
rect 5516 9826 5572 11340
rect 5852 11330 5908 11340
rect 6524 11394 6692 11396
rect 6524 11342 6638 11394
rect 6690 11342 6692 11394
rect 6524 11340 6692 11342
rect 6524 10834 6580 11340
rect 6636 11330 6692 11340
rect 6524 10782 6526 10834
rect 6578 10782 6580 10834
rect 6524 10770 6580 10782
rect 5874 10220 6138 10230
rect 5930 10164 5978 10220
rect 6034 10164 6082 10220
rect 5874 10154 6138 10164
rect 7868 9940 7924 12012
rect 7980 11284 8036 11294
rect 7980 10610 8036 11228
rect 8540 11282 8596 12126
rect 8540 11230 8542 11282
rect 8594 11230 8596 11282
rect 7980 10558 7982 10610
rect 8034 10558 8036 10610
rect 7980 10546 8036 10558
rect 8316 10724 8372 10734
rect 7924 9884 8036 9940
rect 7868 9874 7924 9884
rect 6300 9828 6356 9838
rect 5516 9774 5518 9826
rect 5570 9774 5572 9826
rect 5516 5908 5572 9774
rect 5964 9826 6356 9828
rect 5964 9774 6302 9826
rect 6354 9774 6356 9826
rect 5964 9772 6356 9774
rect 5964 9266 6020 9772
rect 6300 9762 6356 9772
rect 5964 9214 5966 9266
rect 6018 9214 6020 9266
rect 5964 9202 6020 9214
rect 7084 9044 7140 9054
rect 7812 9044 7868 9054
rect 7084 9042 7868 9044
rect 7084 8990 7086 9042
rect 7138 8990 7814 9042
rect 7866 8990 7868 9042
rect 7084 8988 7868 8990
rect 7084 8978 7140 8988
rect 7812 8978 7868 8988
rect 7084 8820 7140 8830
rect 5874 8652 6138 8662
rect 5930 8596 5978 8652
rect 6034 8596 6082 8652
rect 5874 8586 6138 8596
rect 7084 7476 7140 8764
rect 7980 8428 8036 9884
rect 8204 9828 8260 9838
rect 8092 9716 8148 9726
rect 8092 9042 8148 9660
rect 8092 8990 8094 9042
rect 8146 8990 8148 9042
rect 8092 8978 8148 8990
rect 8204 9714 8260 9772
rect 8204 9662 8206 9714
rect 8258 9662 8260 9714
rect 8204 8820 8260 9662
rect 8316 9042 8372 10668
rect 8428 10610 8484 10622
rect 8428 10558 8430 10610
rect 8482 10558 8484 10610
rect 8428 10276 8484 10558
rect 8428 10210 8484 10220
rect 8316 8990 8318 9042
rect 8370 8990 8372 9042
rect 8316 8978 8372 8990
rect 8428 9044 8484 9054
rect 8540 9044 8596 11230
rect 8652 10836 8708 12348
rect 8782 11954 8838 11966
rect 8782 11902 8784 11954
rect 8836 11902 8838 11954
rect 8782 11396 8838 11902
rect 8782 11330 8838 11340
rect 9044 11284 9100 11294
rect 9044 11190 9100 11228
rect 9212 11172 9268 12908
rect 9548 12740 9604 12750
rect 9436 12684 9548 12740
rect 9436 11956 9492 12684
rect 9548 12646 9604 12684
rect 9884 12404 9940 12414
rect 9604 12180 9660 12190
rect 9604 12086 9660 12124
rect 9884 12178 9940 12348
rect 9884 12126 9886 12178
rect 9938 12126 9940 12178
rect 9884 12114 9940 12126
rect 9996 12178 10052 13692
rect 10332 13524 10388 14252
rect 10556 14242 10612 14252
rect 10536 14140 10800 14150
rect 10592 14084 10640 14140
rect 10696 14084 10744 14140
rect 10536 14074 10800 14084
rect 10668 13746 10724 13758
rect 10332 13458 10388 13468
rect 10500 13690 10556 13702
rect 10500 13638 10502 13690
rect 10554 13638 10556 13690
rect 10500 13186 10556 13638
rect 10500 13134 10502 13186
rect 10554 13134 10556 13186
rect 10500 13122 10556 13134
rect 10668 13694 10670 13746
rect 10722 13694 10724 13746
rect 10220 12962 10276 12974
rect 10220 12910 10222 12962
rect 10274 12910 10276 12962
rect 10220 12852 10276 12910
rect 10220 12786 10276 12796
rect 10668 12740 10724 13694
rect 10780 12964 10836 12974
rect 11004 12964 11060 12974
rect 10780 12962 10948 12964
rect 10780 12910 10782 12962
rect 10834 12910 10948 12962
rect 10780 12908 10948 12910
rect 10780 12898 10836 12908
rect 10668 12674 10724 12684
rect 10536 12572 10800 12582
rect 10592 12516 10640 12572
rect 10696 12516 10744 12572
rect 10536 12506 10800 12516
rect 9996 12126 9998 12178
rect 10050 12126 10052 12178
rect 9996 12114 10052 12126
rect 10108 12292 10164 12302
rect 9436 11900 9604 11956
rect 9324 11396 9380 11406
rect 9324 11302 9380 11340
rect 9436 11394 9492 11406
rect 9436 11342 9438 11394
rect 9490 11342 9492 11394
rect 9436 11172 9492 11342
rect 9212 11116 9492 11172
rect 8652 10780 8820 10836
rect 8652 10612 8708 10622
rect 8652 10518 8708 10556
rect 8764 9940 8820 10780
rect 9436 10724 9492 11116
rect 9436 10658 9492 10668
rect 9548 10722 9604 11900
rect 9548 10670 9550 10722
rect 9602 10670 9604 10722
rect 9548 10658 9604 10670
rect 9996 11394 10052 11406
rect 9996 11342 9998 11394
rect 10050 11342 10052 11394
rect 9716 10554 9772 10566
rect 9716 10502 9718 10554
rect 9770 10502 9772 10554
rect 8932 10388 8988 10398
rect 9716 10388 9772 10502
rect 8932 10386 9772 10388
rect 8932 10334 8934 10386
rect 8986 10334 9772 10386
rect 8932 10332 9772 10334
rect 9884 10500 9940 10510
rect 8932 10322 8988 10332
rect 9660 9940 9716 9950
rect 8764 9884 8932 9940
rect 8746 9716 8802 9726
rect 8746 9622 8802 9660
rect 8876 9492 8932 9884
rect 8988 9828 9044 9838
rect 9660 9826 9716 9884
rect 8988 9734 9044 9772
rect 9492 9770 9548 9782
rect 8428 9042 8596 9044
rect 8428 8990 8430 9042
rect 8482 8990 8596 9042
rect 8428 8988 8596 8990
rect 8652 9436 8932 9492
rect 9492 9718 9494 9770
rect 9546 9718 9548 9770
rect 9660 9774 9662 9826
rect 9714 9774 9716 9826
rect 9660 9762 9716 9774
rect 8652 9042 8708 9436
rect 9492 9380 9548 9718
rect 9884 9604 9940 10444
rect 8932 9324 9548 9380
rect 9772 9548 9940 9604
rect 8932 9154 8988 9324
rect 8932 9102 8934 9154
rect 8986 9102 8988 9154
rect 8932 9090 8988 9102
rect 9548 9156 9604 9166
rect 8652 8990 8654 9042
rect 8706 8990 8708 9042
rect 8204 8754 8260 8764
rect 6860 7474 7140 7476
rect 6860 7422 7086 7474
rect 7138 7422 7140 7474
rect 6860 7420 7140 7422
rect 5874 7084 6138 7094
rect 5930 7028 5978 7084
rect 6034 7028 6082 7084
rect 5874 7018 6138 7028
rect 6524 6804 6580 6814
rect 5852 5908 5908 5918
rect 5516 5852 5852 5908
rect 5852 5814 5908 5852
rect 5874 5516 6138 5526
rect 5930 5460 5978 5516
rect 6034 5460 6082 5516
rect 5874 5450 6138 5460
rect 6188 5236 6244 5246
rect 1932 5122 1988 5134
rect 1932 5070 1934 5122
rect 1986 5070 1988 5122
rect 1148 3444 1204 3454
rect 1148 800 1204 3388
rect 1932 3444 1988 5070
rect 4172 5124 4228 5134
rect 4172 5042 4174 5068
rect 4226 5042 4228 5068
rect 4172 5030 4228 5042
rect 3500 5012 3556 5022
rect 2772 4564 2828 4574
rect 2772 4470 2828 4508
rect 3500 4564 3556 4956
rect 6188 4676 6244 5180
rect 6524 5124 6580 6748
rect 6636 6466 6692 6478
rect 6636 6414 6638 6466
rect 6690 6414 6692 6466
rect 6636 5906 6692 6414
rect 6636 5854 6638 5906
rect 6690 5854 6692 5906
rect 6636 5842 6692 5854
rect 6636 5124 6692 5134
rect 6524 5122 6692 5124
rect 6524 5070 6638 5122
rect 6690 5070 6692 5122
rect 6524 5068 6692 5070
rect 6860 5124 6916 7420
rect 7084 7410 7140 7420
rect 7308 8372 7364 8382
rect 7308 7474 7364 8316
rect 7644 8372 8036 8428
rect 7644 8258 7700 8372
rect 7644 8206 7646 8258
rect 7698 8206 7700 8258
rect 7644 8194 7700 8206
rect 7812 8202 7868 8214
rect 7812 8150 7814 8202
rect 7866 8150 7868 8202
rect 7588 7588 7644 7598
rect 7812 7588 7868 8150
rect 7588 7586 7868 7588
rect 7588 7534 7590 7586
rect 7642 7534 7868 7586
rect 7588 7532 7868 7534
rect 7980 7586 8036 8372
rect 8316 8258 8372 8270
rect 8316 8206 8318 8258
rect 8370 8206 8372 8258
rect 8316 8148 8372 8206
rect 8316 8082 8372 8092
rect 7980 7534 7982 7586
rect 8034 7534 8036 7586
rect 7588 7522 7644 7532
rect 7980 7522 8036 7534
rect 8316 7588 8372 7598
rect 7308 7422 7310 7474
rect 7362 7422 7364 7474
rect 7308 7410 7364 7422
rect 8148 7476 8204 7486
rect 8148 7382 8204 7420
rect 7980 7252 8036 7262
rect 7308 5124 7364 5134
rect 6860 5122 7364 5124
rect 6860 5070 7310 5122
rect 7362 5070 7364 5122
rect 6860 5068 7364 5070
rect 6636 5058 6692 5068
rect 7308 5058 7364 5068
rect 7980 5122 8036 7196
rect 8092 6692 8148 6702
rect 8316 6692 8372 7532
rect 8428 7252 8484 8988
rect 8652 8596 8708 8990
rect 8652 8530 8708 8540
rect 8558 8372 8614 8382
rect 8558 8370 9380 8372
rect 8558 8318 8560 8370
rect 8612 8318 9380 8370
rect 8558 8316 9380 8318
rect 8558 8306 8614 8316
rect 9324 8258 9380 8316
rect 9324 8206 9326 8258
rect 9378 8206 9380 8258
rect 9324 8194 9380 8206
rect 9436 8258 9492 8270
rect 9436 8206 9438 8258
rect 9490 8206 9492 8258
rect 8428 7186 8484 7196
rect 8540 8148 8596 8158
rect 8540 7364 8596 8092
rect 9044 8146 9100 8158
rect 9044 8094 9046 8146
rect 9098 8094 9100 8146
rect 9044 7588 9100 8094
rect 9436 8036 9492 8206
rect 9436 7970 9492 7980
rect 9044 7522 9100 7532
rect 8092 6690 8372 6692
rect 8092 6638 8094 6690
rect 8146 6638 8372 6690
rect 8092 6636 8372 6638
rect 8540 6804 8596 7308
rect 8092 6626 8148 6636
rect 8540 6018 8596 6748
rect 8540 5966 8542 6018
rect 8594 5966 8596 6018
rect 8540 5954 8596 5966
rect 8652 7474 8708 7486
rect 8652 7422 8654 7474
rect 8706 7422 8708 7474
rect 8652 6580 8708 7422
rect 9436 7474 9492 7486
rect 9436 7422 9438 7474
rect 9490 7422 9492 7474
rect 9436 7364 9492 7422
rect 9436 7298 9492 7308
rect 8894 7250 8950 7262
rect 8894 7198 8896 7250
rect 8948 7198 8950 7250
rect 8894 6692 8950 7198
rect 8894 6626 8950 6636
rect 8316 5236 8372 5246
rect 8652 5236 8708 6524
rect 9548 6580 9604 9100
rect 9772 9154 9828 9548
rect 9772 9102 9774 9154
rect 9826 9102 9828 9154
rect 9660 8372 9716 8382
rect 9660 7474 9716 8316
rect 9660 7422 9662 7474
rect 9714 7422 9716 7474
rect 9660 7410 9716 7422
rect 9548 6514 9604 6524
rect 8372 5180 8708 5236
rect 8988 6466 9044 6478
rect 8988 6414 8990 6466
rect 9042 6414 9044 6466
rect 8988 5236 9044 6414
rect 9772 6132 9828 9102
rect 9996 9156 10052 11342
rect 10108 11394 10164 12236
rect 10668 12292 10724 12302
rect 10668 12198 10724 12236
rect 10892 12292 10948 12908
rect 11004 12870 11060 12908
rect 11116 12962 11172 14700
rect 11508 14690 11564 14700
rect 12124 14654 12180 15486
rect 12460 15316 12516 15326
rect 12460 15222 12516 15260
rect 13468 15316 13524 15326
rect 12068 14642 12180 14654
rect 12068 14590 12070 14642
rect 12122 14590 12180 14642
rect 12068 14588 12180 14590
rect 12068 14578 12124 14588
rect 11116 12910 11118 12962
rect 11170 12910 11172 12962
rect 11116 12898 11172 12910
rect 11228 14530 11284 14542
rect 11228 14478 11230 14530
rect 11282 14478 11284 14530
rect 10892 12226 10948 12236
rect 11004 12404 11060 12414
rect 11004 12180 11060 12348
rect 11228 12180 11284 14478
rect 11452 13634 11508 13646
rect 13356 13636 13412 13646
rect 11452 13582 11454 13634
rect 11506 13582 11508 13634
rect 11452 12964 11508 13582
rect 13132 13634 13412 13636
rect 13132 13582 13358 13634
rect 13410 13582 13412 13634
rect 13132 13580 13412 13582
rect 13132 13300 13188 13580
rect 13356 13570 13412 13580
rect 12572 13244 13188 13300
rect 12572 13186 12628 13244
rect 12572 13134 12574 13186
rect 12626 13134 12628 13186
rect 12572 13122 12628 13134
rect 11452 12180 11508 12908
rect 11900 12740 11956 12750
rect 11900 12346 11956 12684
rect 11900 12294 11902 12346
rect 11954 12294 11956 12346
rect 11564 12180 11620 12190
rect 11228 12124 11378 12180
rect 11452 12178 11620 12180
rect 11452 12126 11566 12178
rect 11618 12126 11620 12178
rect 11452 12124 11620 12126
rect 11004 12086 11060 12124
rect 11322 12066 11378 12124
rect 11564 12114 11620 12124
rect 11322 12014 11324 12066
rect 11376 12014 11378 12066
rect 11322 12002 11378 12014
rect 10668 11620 10724 11630
rect 10108 11342 10110 11394
rect 10162 11342 10164 11394
rect 10108 10836 10164 11342
rect 10388 11396 10444 11406
rect 10388 11302 10444 11340
rect 10668 11394 10724 11564
rect 10668 11342 10670 11394
rect 10722 11342 10724 11394
rect 10668 11330 10724 11342
rect 11900 11394 11956 12294
rect 12068 12180 12124 12190
rect 12068 12086 12124 12124
rect 12740 12068 12796 12078
rect 12684 12066 12796 12068
rect 12684 12014 12742 12066
rect 12794 12014 12796 12066
rect 12684 12002 12796 12014
rect 13132 12068 13188 12078
rect 12236 11620 12292 11630
rect 11900 11342 11902 11394
rect 11954 11342 11956 11394
rect 11900 11330 11956 11342
rect 12068 11396 12124 11406
rect 12068 11302 12124 11340
rect 10536 11004 10800 11014
rect 10592 10948 10640 11004
rect 10696 10948 10744 11004
rect 10536 10938 10800 10948
rect 10108 10770 10164 10780
rect 12236 10834 12292 11564
rect 12236 10782 12238 10834
rect 12290 10782 12292 10834
rect 11228 10637 11284 10649
rect 10220 10610 10276 10622
rect 10220 10558 10222 10610
rect 10274 10558 10276 10610
rect 10220 10500 10276 10558
rect 10220 10434 10276 10444
rect 11228 10585 11230 10637
rect 11282 10585 11284 10637
rect 10462 10386 10518 10398
rect 10462 10334 10464 10386
rect 10516 10334 10518 10386
rect 10164 10276 10220 10286
rect 10164 9940 10220 10220
rect 10462 10052 10518 10334
rect 11228 10164 11284 10585
rect 11228 10098 11284 10108
rect 10462 9986 10518 9996
rect 11788 10052 11844 10062
rect 10164 9938 10276 9940
rect 10164 9886 10166 9938
rect 10218 9886 10276 9938
rect 10164 9874 10276 9886
rect 9996 9090 10052 9100
rect 9940 8036 9996 8046
rect 9940 7942 9996 7980
rect 9940 7476 9996 7486
rect 9940 7382 9996 7420
rect 10220 6916 10276 9874
rect 10444 9828 10500 9838
rect 10444 9826 11508 9828
rect 10444 9774 10446 9826
rect 10498 9774 11508 9826
rect 10444 9772 11508 9774
rect 10444 9762 10500 9772
rect 10536 9436 10800 9446
rect 10592 9380 10640 9436
rect 10696 9380 10744 9436
rect 10536 9370 10800 9380
rect 11452 8494 11508 9772
rect 11564 9604 11620 9614
rect 11564 9602 11732 9604
rect 11564 9550 11566 9602
rect 11618 9550 11732 9602
rect 11564 9548 11732 9550
rect 11564 9538 11620 9548
rect 11676 9042 11732 9548
rect 11676 8990 11678 9042
rect 11730 8990 11732 9042
rect 11676 8978 11732 8990
rect 11452 8482 11564 8494
rect 11452 8430 11510 8482
rect 11562 8430 11564 8482
rect 11452 8428 11564 8430
rect 11508 8418 11564 8428
rect 11788 8258 11844 9996
rect 12236 9044 12292 10782
rect 12572 11508 12628 11518
rect 12684 11508 12740 12002
rect 13132 11974 13188 12012
rect 12628 11452 12740 11508
rect 12572 11394 12628 11452
rect 12572 11342 12574 11394
rect 12626 11342 12628 11394
rect 12572 10276 12628 11342
rect 12814 11396 12870 11406
rect 12814 11302 12870 11340
rect 13468 10612 13524 15260
rect 13580 14756 13636 14766
rect 13580 13860 13636 14700
rect 13580 13794 13636 13804
rect 13692 13412 13748 16830
rect 14028 14756 14084 19068
rect 14364 18788 14420 18798
rect 14140 18452 14196 18462
rect 14140 17668 14196 18396
rect 14140 17666 14308 17668
rect 14140 17614 14142 17666
rect 14194 17614 14308 17666
rect 14140 17612 14308 17614
rect 14140 17602 14196 17612
rect 14252 15316 14308 17612
rect 14252 15250 14308 15260
rect 13692 13346 13748 13356
rect 13804 14700 14084 14756
rect 13636 13188 13692 13198
rect 13636 13074 13692 13132
rect 13636 13022 13638 13074
rect 13690 13022 13692 13074
rect 13636 12404 13692 13022
rect 13636 12338 13692 12348
rect 13804 12852 13860 14700
rect 13916 14530 13972 14542
rect 14364 14532 14420 18732
rect 14476 17442 14532 17454
rect 14476 17390 14478 17442
rect 14530 17390 14532 17442
rect 14476 17220 14532 17390
rect 14476 17154 14532 17164
rect 14812 17108 14868 21868
rect 15198 21196 15462 21206
rect 15254 21140 15302 21196
rect 15358 21140 15406 21196
rect 15198 21130 15462 21140
rect 14980 20578 15036 20590
rect 14980 20526 14982 20578
rect 15034 20526 15036 20578
rect 14980 20188 15036 20526
rect 14924 20132 15036 20188
rect 15316 20578 15372 20590
rect 15316 20526 15318 20578
rect 15370 20526 15372 20578
rect 15316 20242 15372 20526
rect 15316 20190 15318 20242
rect 15370 20190 15372 20242
rect 14924 18788 14980 20132
rect 15316 19796 15372 20190
rect 15596 19908 15652 21980
rect 15932 21822 15988 22316
rect 16044 22306 16100 22316
rect 16604 21924 16660 23324
rect 16716 23156 16772 23886
rect 17052 23714 17108 28364
rect 17052 23662 17054 23714
rect 17106 23662 17108 23714
rect 16940 23156 16996 23166
rect 16716 23100 16940 23156
rect 16940 23062 16996 23100
rect 16828 22372 16884 22382
rect 16828 22278 16884 22316
rect 16604 21858 16660 21868
rect 15876 21810 15988 21822
rect 15876 21758 15878 21810
rect 15930 21758 15988 21810
rect 15876 21746 15988 21758
rect 15932 20578 15988 21746
rect 15932 20526 15934 20578
rect 15986 20526 15988 20578
rect 15932 20514 15988 20526
rect 15596 19842 15652 19852
rect 15764 19906 15820 19918
rect 15764 19854 15766 19906
rect 15818 19854 15820 19906
rect 15036 19740 15372 19796
rect 15764 19796 15820 19854
rect 15036 19460 15092 19740
rect 15764 19730 15820 19740
rect 15198 19628 15462 19638
rect 15254 19572 15302 19628
rect 15358 19572 15406 19628
rect 15198 19562 15462 19572
rect 15036 19404 15204 19460
rect 14924 18722 14980 18732
rect 15148 18228 15204 19404
rect 15260 19234 15316 19246
rect 15260 19182 15262 19234
rect 15314 19182 15316 19234
rect 15260 18674 15316 19182
rect 15260 18622 15262 18674
rect 15314 18622 15316 18674
rect 15260 18610 15316 18622
rect 15036 18172 15204 18228
rect 15036 17892 15092 18172
rect 15198 18060 15462 18070
rect 15254 18004 15302 18060
rect 15358 18004 15406 18060
rect 15198 17994 15462 18004
rect 15036 17836 15204 17892
rect 15148 17678 15204 17836
rect 15092 17666 15204 17678
rect 15092 17614 15094 17666
rect 15146 17614 15204 17666
rect 15092 17612 15204 17614
rect 15092 17602 15148 17612
rect 14700 17052 14868 17108
rect 15596 17220 15652 17230
rect 14476 16770 14532 16782
rect 14476 16718 14478 16770
rect 14530 16718 14532 16770
rect 14476 16322 14532 16718
rect 14476 16270 14478 16322
rect 14530 16270 14532 16322
rect 14476 16258 14532 16270
rect 13916 14478 13918 14530
rect 13970 14478 13972 14530
rect 13916 14308 13972 14478
rect 13916 13076 13972 14252
rect 14028 14476 14420 14532
rect 14028 13188 14084 14476
rect 14308 14308 14364 14318
rect 14308 14214 14364 14252
rect 14476 14196 14532 14206
rect 14476 13860 14532 14140
rect 14700 14196 14756 17052
rect 15198 16492 15462 16502
rect 15254 16436 15302 16492
rect 15358 16436 15406 16492
rect 15198 16426 15462 16436
rect 15372 16100 15428 16110
rect 15596 16100 15652 17164
rect 16380 16996 16436 17006
rect 16380 16902 16436 16940
rect 15204 16098 15652 16100
rect 15204 16046 15374 16098
rect 15426 16046 15652 16098
rect 15204 16044 15652 16046
rect 16716 16436 16772 16446
rect 15204 15538 15260 16044
rect 15372 16034 15428 16044
rect 15204 15486 15206 15538
rect 15258 15486 15260 15538
rect 15204 15474 15260 15486
rect 15708 15874 15764 15886
rect 15708 15822 15710 15874
rect 15762 15822 15764 15874
rect 15198 14924 15462 14934
rect 15254 14868 15302 14924
rect 15358 14868 15406 14924
rect 15198 14858 15462 14868
rect 14700 14084 14756 14140
rect 14700 14028 15148 14084
rect 15092 13970 15148 14028
rect 15092 13918 15094 13970
rect 15146 13918 15148 13970
rect 15092 13906 15148 13918
rect 14364 13804 14532 13860
rect 14924 13860 14980 13870
rect 14140 13746 14196 13758
rect 14140 13694 14142 13746
rect 14194 13694 14196 13746
rect 14140 13412 14196 13694
rect 14140 13346 14196 13356
rect 14028 13122 14084 13132
rect 13916 13010 13972 13020
rect 14196 13076 14252 13086
rect 14196 12982 14252 13020
rect 14364 12962 14420 13804
rect 14532 13634 14588 13646
rect 14532 13582 14534 13634
rect 14586 13582 14588 13634
rect 14532 13412 14588 13582
rect 14532 13346 14588 13356
rect 14364 12910 14366 12962
rect 14418 12910 14420 12962
rect 14364 12852 14420 12910
rect 13804 12178 13860 12796
rect 14252 12796 14420 12852
rect 13804 12126 13806 12178
rect 13858 12126 13860 12178
rect 13804 12114 13860 12126
rect 14084 12180 14140 12190
rect 14084 12086 14140 12124
rect 14140 11844 14196 11854
rect 14028 11396 14084 11406
rect 14028 11302 14084 11340
rect 14140 11394 14196 11788
rect 14140 11342 14142 11394
rect 14194 11342 14196 11394
rect 13748 11284 13804 11294
rect 13748 11190 13804 11228
rect 13468 10546 13524 10556
rect 12572 10210 12628 10220
rect 13916 10386 13972 10398
rect 13916 10334 13918 10386
rect 13970 10334 13972 10386
rect 12964 10164 13020 10174
rect 12964 9940 13020 10108
rect 12964 9846 13020 9884
rect 13804 9826 13860 9838
rect 13804 9774 13806 9826
rect 13858 9774 13860 9826
rect 12796 9716 12852 9726
rect 12460 9044 12516 9054
rect 12236 9042 12516 9044
rect 12236 8990 12462 9042
rect 12514 8990 12516 9042
rect 12236 8988 12516 8990
rect 12460 8978 12516 8988
rect 12796 9042 12852 9660
rect 13524 9716 13580 9726
rect 13524 9622 13580 9660
rect 12796 8990 12798 9042
rect 12850 8990 12852 9042
rect 12796 8978 12852 8990
rect 13562 8484 13618 8494
rect 13804 8484 13860 9774
rect 13562 8482 13860 8484
rect 13562 8430 13564 8482
rect 13616 8430 13860 8482
rect 13562 8428 13860 8430
rect 13916 9826 13972 10334
rect 14140 10276 14196 11342
rect 14252 10610 14308 12796
rect 14588 12740 14644 12750
rect 14364 12292 14420 12302
rect 14364 12178 14420 12236
rect 14364 12126 14366 12178
rect 14418 12126 14420 12178
rect 14364 12114 14420 12126
rect 14588 12178 14644 12684
rect 14588 12126 14590 12178
rect 14642 12126 14644 12178
rect 14588 12114 14644 12126
rect 14700 12738 14756 12750
rect 14700 12686 14702 12738
rect 14754 12686 14756 12738
rect 14700 12404 14756 12686
rect 14700 11844 14756 12348
rect 14924 12180 14980 13804
rect 15708 13860 15764 15822
rect 15708 13794 15764 13804
rect 16492 13746 16548 13758
rect 16492 13694 16494 13746
rect 16546 13694 16548 13746
rect 16156 13524 16212 13534
rect 15820 13522 16212 13524
rect 15820 13470 16158 13522
rect 16210 13470 16212 13522
rect 15820 13468 16212 13470
rect 15036 13412 15092 13422
rect 15036 12962 15092 13356
rect 15198 13356 15462 13366
rect 15254 13300 15302 13356
rect 15358 13300 15406 13356
rect 15198 13290 15462 13300
rect 15820 13074 15876 13468
rect 16156 13458 16212 13468
rect 16492 13300 16548 13694
rect 15820 13022 15822 13074
rect 15874 13022 15876 13074
rect 15820 13010 15876 13022
rect 16044 13244 16548 13300
rect 16716 13300 16772 16380
rect 16940 14532 16996 14542
rect 16940 14438 16996 14476
rect 16716 13244 16996 13300
rect 15036 12910 15038 12962
rect 15090 12910 15092 12962
rect 15036 12852 15092 12910
rect 15036 12414 15092 12796
rect 16044 12740 16100 13244
rect 16940 12740 16996 13244
rect 16044 12684 16268 12740
rect 15036 12404 15148 12414
rect 15036 12402 15316 12404
rect 15036 12350 15094 12402
rect 15146 12350 15316 12402
rect 15036 12348 15316 12350
rect 15092 12338 15148 12348
rect 14924 12124 15092 12180
rect 14700 11778 14756 11788
rect 14588 11508 14644 11518
rect 14588 11414 14644 11452
rect 14252 10558 14254 10610
rect 14306 10558 14308 10610
rect 14252 10388 14308 10558
rect 14364 11284 14420 11294
rect 14364 10610 14420 11228
rect 14364 10558 14366 10610
rect 14418 10558 14420 10610
rect 14364 10546 14420 10558
rect 14252 10332 14924 10388
rect 14140 10220 14476 10276
rect 14420 9938 14476 10220
rect 14420 9886 14422 9938
rect 14474 9886 14476 9938
rect 14420 9874 14476 9886
rect 14868 9938 14924 10332
rect 14868 9886 14870 9938
rect 14922 9886 14924 9938
rect 14868 9874 14924 9886
rect 13916 9774 13918 9826
rect 13970 9774 13972 9826
rect 13562 8418 13618 8428
rect 11788 8206 11790 8258
rect 11842 8206 11844 8258
rect 11788 8194 11844 8206
rect 12012 8260 12068 8270
rect 12460 8260 12516 8270
rect 12012 8258 12180 8260
rect 12012 8206 12014 8258
rect 12066 8206 12180 8258
rect 12012 8204 12180 8206
rect 12012 8194 12068 8204
rect 11060 8036 11116 8046
rect 10536 7868 10800 7878
rect 10592 7812 10640 7868
rect 10696 7812 10744 7868
rect 10536 7802 10800 7812
rect 11060 7812 11116 7980
rect 11060 7700 11116 7756
rect 10780 7698 11116 7700
rect 10780 7646 11062 7698
rect 11114 7646 11116 7698
rect 10780 7644 11116 7646
rect 10220 6860 10612 6916
rect 10108 6692 10164 6702
rect 10388 6692 10444 6702
rect 10108 6690 10444 6692
rect 10108 6638 10110 6690
rect 10162 6638 10390 6690
rect 10442 6638 10444 6690
rect 10108 6636 10444 6638
rect 10108 6626 10164 6636
rect 10388 6626 10444 6636
rect 10108 6468 10164 6478
rect 10556 6468 10612 6860
rect 10668 6692 10724 6702
rect 10668 6598 10724 6636
rect 10780 6690 10836 7644
rect 11060 7634 11116 7644
rect 10780 6638 10782 6690
rect 10834 6638 10836 6690
rect 10780 6626 10836 6638
rect 10892 7476 10948 7486
rect 9660 6076 9828 6132
rect 9996 6132 10052 6142
rect 9660 5684 9716 6076
rect 9996 6074 10052 6076
rect 9996 6022 9998 6074
rect 10050 6022 10052 6074
rect 9996 6010 10052 6022
rect 9940 5908 9996 5918
rect 10108 5908 10164 6412
rect 9940 5906 10164 5908
rect 9940 5854 9942 5906
rect 9994 5854 10164 5906
rect 9940 5852 10164 5854
rect 9940 5842 9996 5852
rect 9660 5628 10052 5684
rect 8316 5142 8372 5180
rect 8988 5170 9044 5180
rect 7980 5070 7982 5122
rect 8034 5070 8036 5122
rect 7980 5058 8036 5070
rect 9100 5124 9156 5134
rect 6300 4900 6356 4910
rect 6972 4900 7028 4910
rect 6300 4898 6580 4900
rect 6300 4846 6302 4898
rect 6354 4846 6580 4898
rect 6300 4844 6580 4846
rect 6300 4834 6356 4844
rect 6188 4620 6356 4676
rect 3500 4338 3556 4508
rect 3500 4286 3502 4338
rect 3554 4286 3556 4338
rect 3500 4274 3556 4286
rect 5852 4365 5908 4377
rect 5852 4313 5854 4365
rect 5906 4313 5908 4365
rect 3164 4116 3220 4126
rect 4844 4116 4900 4126
rect 5852 4116 5908 4313
rect 2940 4114 3220 4116
rect 2940 4062 3166 4114
rect 3218 4062 3220 4114
rect 2940 4060 3220 4062
rect 2940 3780 2996 4060
rect 3164 4050 3220 4060
rect 4732 4114 4900 4116
rect 4732 4062 4846 4114
rect 4898 4062 4900 4114
rect 4732 4060 4900 4062
rect 2828 3724 2996 3780
rect 2828 3526 2884 3724
rect 2828 3474 2830 3526
rect 2882 3474 2884 3526
rect 2828 3462 2884 3474
rect 3500 3666 3556 3678
rect 3500 3614 3502 3666
rect 3554 3614 3556 3666
rect 1932 3378 1988 3388
rect 2940 3444 2996 3454
rect 2940 800 2996 3388
rect 3500 3444 3556 3614
rect 3500 3378 3556 3388
rect 4732 800 4788 4060
rect 4844 4050 4900 4060
rect 5740 4060 5908 4116
rect 5740 3778 5796 4060
rect 5874 3948 6138 3958
rect 5930 3892 5978 3948
rect 6034 3892 6082 3948
rect 5874 3882 6138 3892
rect 5740 3726 5742 3778
rect 5794 3726 5796 3778
rect 5740 3714 5796 3726
rect 6076 3556 6132 3566
rect 6300 3556 6356 4620
rect 6524 4365 6580 4844
rect 6524 4313 6526 4365
rect 6578 4313 6580 4365
rect 6524 4301 6580 4313
rect 6636 4898 7028 4900
rect 6636 4846 6974 4898
rect 7026 4846 7028 4898
rect 6636 4844 7028 4846
rect 6076 3554 6356 3556
rect 6076 3502 6078 3554
rect 6130 3502 6356 3554
rect 6076 3500 6356 3502
rect 6524 4116 6580 4126
rect 6076 3490 6132 3500
rect 6524 800 6580 4060
rect 6636 3526 6692 4844
rect 6972 4834 7028 4844
rect 7644 4900 7700 4910
rect 7644 4806 7700 4844
rect 9100 4228 9156 5068
rect 9100 4172 9604 4228
rect 7532 4116 7588 4126
rect 7532 4022 7588 4060
rect 9548 3778 9604 4172
rect 9548 3726 9550 3778
rect 9602 3726 9604 3778
rect 9548 3714 9604 3726
rect 6636 3474 6638 3526
rect 6690 3474 6692 3526
rect 6636 3462 6692 3474
rect 8316 3554 8372 3566
rect 8316 3502 8318 3554
rect 8370 3502 8372 3554
rect 8316 800 8372 3502
rect 9884 3556 9940 3566
rect 9996 3556 10052 5628
rect 10108 5012 10164 5852
rect 10332 6412 10612 6468
rect 10220 5236 10276 5246
rect 10220 5142 10276 5180
rect 10332 5012 10388 6412
rect 10536 6300 10800 6310
rect 10592 6244 10640 6300
rect 10696 6244 10744 6300
rect 10536 6234 10800 6244
rect 10892 6132 10948 7420
rect 11900 7476 11956 7486
rect 11900 7382 11956 7420
rect 12124 7476 12180 8204
rect 12124 7382 12180 7420
rect 12460 7586 12516 8204
rect 13804 8260 13860 8270
rect 13804 8166 13860 8204
rect 13916 7700 13972 9774
rect 14252 8820 14308 8830
rect 13916 7634 13972 7644
rect 14140 8818 14308 8820
rect 14140 8766 14254 8818
rect 14306 8766 14308 8818
rect 14140 8764 14308 8766
rect 12460 7534 12462 7586
rect 12514 7534 12516 7586
rect 11620 7252 11676 7262
rect 11228 7250 11676 7252
rect 11228 7198 11622 7250
rect 11674 7198 11676 7250
rect 11228 7196 11676 7198
rect 11116 6692 11172 6702
rect 11228 6692 11284 7196
rect 11620 7186 11676 7196
rect 12460 6804 12516 7534
rect 14140 7476 14196 8764
rect 14252 8754 14308 8764
rect 15036 8382 15092 12124
rect 15260 12178 15316 12348
rect 16212 12290 16268 12684
rect 16212 12238 16214 12290
rect 16266 12238 16268 12290
rect 16212 12226 16268 12238
rect 16716 12684 16996 12740
rect 15260 12126 15262 12178
rect 15314 12126 15316 12178
rect 15260 12114 15316 12126
rect 16492 12178 16548 12190
rect 16492 12126 16494 12178
rect 16546 12126 16548 12178
rect 16492 11956 16548 12126
rect 16716 12178 16772 12684
rect 16716 12126 16718 12178
rect 16770 12126 16772 12178
rect 16716 12114 16772 12126
rect 17052 11956 17108 23662
rect 17164 23380 17220 28476
rect 17276 27188 17332 30268
rect 17724 30826 17780 30838
rect 17724 30774 17726 30826
rect 17778 30774 17780 30826
rect 17612 30212 17668 30222
rect 17612 30118 17668 30156
rect 17724 29764 17780 30774
rect 17948 30436 18004 30446
rect 18060 30436 18116 31726
rect 17948 30434 18116 30436
rect 17948 30382 17950 30434
rect 18002 30382 18116 30434
rect 17948 30380 18116 30382
rect 17948 30370 18004 30380
rect 17724 29708 18004 29764
rect 17556 29316 17612 29326
rect 17500 29314 17612 29316
rect 17500 29262 17558 29314
rect 17610 29262 17612 29314
rect 17500 29250 17612 29262
rect 17388 28754 17444 28766
rect 17388 28702 17390 28754
rect 17442 28702 17444 28754
rect 17388 28644 17444 28702
rect 17388 28578 17444 28588
rect 17388 28420 17444 28430
rect 17500 28420 17556 29250
rect 17948 28642 18004 29708
rect 18284 29540 18340 32732
rect 18396 32589 18452 32601
rect 18396 32537 18398 32589
rect 18450 32537 18452 32589
rect 18396 32340 18452 32537
rect 18732 32562 18788 33740
rect 18956 33572 19012 33582
rect 18956 33478 19012 33516
rect 19404 33236 19460 33246
rect 20076 33236 20132 34300
rect 20412 34262 20468 34300
rect 19460 33180 19516 33236
rect 19404 33170 19516 33180
rect 20076 33170 20132 33180
rect 20412 33236 20468 33246
rect 18732 32510 18734 32562
rect 18786 32510 18788 32562
rect 18732 32498 18788 32510
rect 18844 32730 18900 32742
rect 18844 32678 18846 32730
rect 18898 32678 18900 32730
rect 18396 32274 18452 32284
rect 18844 32116 18900 32678
rect 19460 32618 19516 33170
rect 19860 32956 20124 32966
rect 19916 32900 19964 32956
rect 20020 32900 20068 32956
rect 19860 32890 20124 32900
rect 19292 32562 19348 32574
rect 19292 32510 19294 32562
rect 19346 32510 19348 32562
rect 19460 32566 19462 32618
rect 19514 32566 19516 32618
rect 19460 32554 19516 32566
rect 19628 32676 19684 32686
rect 19292 32340 19348 32510
rect 19292 32274 19348 32284
rect 19628 32228 19684 32620
rect 18844 32050 18900 32060
rect 19516 32172 19684 32228
rect 19740 32562 19796 32574
rect 19740 32510 19742 32562
rect 19794 32510 19796 32562
rect 19516 31220 19572 32172
rect 19740 31892 19796 32510
rect 20020 32564 20076 32574
rect 20020 32470 20076 32508
rect 20412 32562 20468 33180
rect 20636 33124 20692 34860
rect 20972 34804 21028 35308
rect 21084 35252 21140 39200
rect 22204 37828 22260 39200
rect 22204 37772 22708 37828
rect 21084 35186 21140 35196
rect 21756 35588 21812 35598
rect 20860 34748 21028 34804
rect 21532 34886 21588 34898
rect 21532 34834 21534 34886
rect 21586 34834 21588 34886
rect 20636 33068 20726 33124
rect 20670 32600 20726 33068
rect 20412 32510 20414 32562
rect 20466 32510 20468 32562
rect 20076 32116 20132 32126
rect 19740 31826 19796 31836
rect 19964 31892 20020 31902
rect 19964 31798 20020 31836
rect 20076 31892 20132 32060
rect 20076 31836 20356 31892
rect 20076 31556 20132 31836
rect 20300 31778 20356 31836
rect 20300 31726 20302 31778
rect 20354 31726 20356 31778
rect 20300 31714 20356 31726
rect 19516 31154 19572 31164
rect 19628 31500 20132 31556
rect 19516 30996 19572 31006
rect 19404 30940 19516 30996
rect 19292 29988 19348 29998
rect 18284 29474 18340 29484
rect 19068 29986 19348 29988
rect 19068 29934 19294 29986
rect 19346 29934 19348 29986
rect 19068 29932 19348 29934
rect 18396 29428 18452 29438
rect 18228 29316 18284 29326
rect 18396 29316 18452 29372
rect 18228 29314 18452 29316
rect 18228 29262 18230 29314
rect 18282 29262 18452 29314
rect 18228 29260 18452 29262
rect 18228 29250 18284 29260
rect 17444 28364 17556 28420
rect 17782 28586 17838 28598
rect 17782 28534 17784 28586
rect 17836 28534 17838 28586
rect 17948 28590 17950 28642
rect 18002 28590 18004 28642
rect 17948 28578 18004 28590
rect 18060 28642 18116 28654
rect 18060 28590 18062 28642
rect 18114 28590 18116 28642
rect 17388 28354 17444 28364
rect 17276 27122 17332 27132
rect 17388 28196 17444 28206
rect 17388 27074 17444 28140
rect 17782 28084 17838 28534
rect 18060 28196 18116 28590
rect 18396 28532 18452 29260
rect 18676 29314 18732 29326
rect 18676 29262 18678 29314
rect 18730 29262 18732 29314
rect 18676 29092 18732 29262
rect 18676 29026 18732 29036
rect 19068 28756 19124 29932
rect 19292 29922 19348 29932
rect 19404 29596 19460 30940
rect 19516 30902 19572 30940
rect 19628 30212 19684 31500
rect 19860 31388 20124 31398
rect 19916 31332 19964 31388
rect 20020 31332 20068 31388
rect 19860 31322 20124 31332
rect 19852 31220 19908 31230
rect 19852 30994 19908 31164
rect 20076 31108 20132 31118
rect 19852 30942 19854 30994
rect 19906 30942 19908 30994
rect 19852 30930 19908 30942
rect 19964 30994 20020 31006
rect 19964 30942 19966 30994
rect 20018 30942 20020 30994
rect 19964 30772 20020 30942
rect 19964 30706 20020 30716
rect 19628 30118 19684 30156
rect 19908 30100 19964 30110
rect 19348 29540 19460 29596
rect 19740 30098 19964 30100
rect 19740 30046 19910 30098
rect 19962 30046 19964 30098
rect 19740 30044 19964 30046
rect 19348 29482 19404 29540
rect 19180 29426 19236 29438
rect 19180 29374 19182 29426
rect 19234 29374 19236 29426
rect 19348 29430 19350 29482
rect 19402 29430 19404 29482
rect 19348 29418 19404 29430
rect 19516 29428 19572 29438
rect 19180 28868 19236 29374
rect 19516 29334 19572 29372
rect 19628 29426 19684 29438
rect 19628 29374 19630 29426
rect 19682 29374 19684 29426
rect 19404 29204 19460 29214
rect 19180 28812 19348 28868
rect 18732 28700 19180 28756
rect 18732 28642 18788 28700
rect 18732 28590 18734 28642
rect 18786 28590 18788 28642
rect 18732 28578 18788 28590
rect 19124 28698 19180 28700
rect 19124 28646 19126 28698
rect 19178 28646 19180 28698
rect 19124 28644 19180 28646
rect 19124 28568 19180 28588
rect 18396 28466 18452 28476
rect 18956 28530 19012 28542
rect 18956 28478 18958 28530
rect 19010 28478 19012 28530
rect 18564 28420 18620 28430
rect 18564 28418 18900 28420
rect 18564 28366 18566 28418
rect 18618 28366 18900 28418
rect 18564 28364 18900 28366
rect 18564 28354 18620 28364
rect 18060 28130 18116 28140
rect 18732 28196 18788 28206
rect 18284 28084 18340 28094
rect 17782 28028 17892 28084
rect 17500 27860 17556 27870
rect 17836 27860 17892 28028
rect 18284 27990 18340 28028
rect 17948 27860 18004 27870
rect 18732 27860 18788 28140
rect 17500 27634 17556 27804
rect 17500 27582 17502 27634
rect 17554 27582 17556 27634
rect 17500 27524 17556 27582
rect 17500 27458 17556 27468
rect 17724 27858 17948 27860
rect 17724 27806 17838 27858
rect 17890 27806 17948 27858
rect 17724 27804 17948 27806
rect 17724 27298 17780 27804
rect 17836 27794 17892 27804
rect 17948 27766 18004 27804
rect 18396 27858 18788 27860
rect 18396 27806 18734 27858
rect 18786 27806 18788 27858
rect 18396 27804 18788 27806
rect 18396 27412 18452 27804
rect 18732 27794 18788 27804
rect 18844 27858 18900 28364
rect 18956 28196 19012 28478
rect 18956 28130 19012 28140
rect 18844 27806 18846 27858
rect 18898 27806 18900 27858
rect 18844 27794 18900 27806
rect 19010 27860 19066 27870
rect 19010 27766 19066 27804
rect 19292 27636 19348 28812
rect 19404 27746 19460 29148
rect 19628 29204 19684 29374
rect 19628 29138 19684 29148
rect 19516 29092 19572 29102
rect 19516 28980 19572 29036
rect 19516 28924 19684 28980
rect 19404 27694 19406 27746
rect 19458 27694 19460 27746
rect 19404 27682 19460 27694
rect 19628 28642 19684 28924
rect 19628 28590 19630 28642
rect 19682 28590 19684 28642
rect 18396 27346 18452 27356
rect 18564 27580 19348 27636
rect 19628 27636 19684 28590
rect 19740 27860 19796 30044
rect 19908 30034 19964 30044
rect 20076 29988 20132 31052
rect 20412 31024 20468 32510
rect 20524 32564 20580 32574
rect 20670 32548 20672 32600
rect 20724 32548 20726 32600
rect 20670 32536 20726 32548
rect 20524 32470 20580 32508
rect 20636 31556 20692 31566
rect 20636 31462 20692 31500
rect 20860 31220 20916 34748
rect 21308 33290 21364 33302
rect 21308 33238 21310 33290
rect 21362 33238 21364 33290
rect 21308 33236 21364 33238
rect 21308 33170 21364 33180
rect 21420 33290 21476 33302
rect 21420 33238 21422 33290
rect 21474 33238 21476 33290
rect 21420 32788 21476 33238
rect 20860 31154 20916 31164
rect 20972 32732 21476 32788
rect 20972 31108 21028 32732
rect 21420 32564 21476 32574
rect 21084 32562 21476 32564
rect 21084 32510 21422 32562
rect 21474 32510 21476 32562
rect 21084 32508 21476 32510
rect 21084 32450 21140 32508
rect 21420 32498 21476 32508
rect 21084 32398 21086 32450
rect 21138 32398 21140 32450
rect 21084 32386 21140 32398
rect 21532 32004 21588 34834
rect 21756 32788 21812 35532
rect 22316 35252 22372 35262
rect 21868 35140 21924 35150
rect 21868 34130 21924 35084
rect 22316 35138 22372 35196
rect 22316 35086 22318 35138
rect 22370 35086 22372 35138
rect 22316 35074 22372 35086
rect 22652 35028 22708 37772
rect 22764 36482 22820 36494
rect 22764 36430 22766 36482
rect 22818 36430 22820 36482
rect 22764 35812 22820 36430
rect 22764 35746 22820 35756
rect 22876 35588 22932 35598
rect 22652 34962 22708 34972
rect 22764 35586 22932 35588
rect 22764 35534 22878 35586
rect 22930 35534 22932 35586
rect 22764 35532 22932 35534
rect 21868 34078 21870 34130
rect 21922 34078 21924 34130
rect 21868 34066 21924 34078
rect 22652 34020 22708 34030
rect 22540 34018 22708 34020
rect 22540 33966 22654 34018
rect 22706 33966 22708 34018
rect 22540 33964 22708 33966
rect 22148 33348 22204 33358
rect 22148 33254 22204 33292
rect 22316 33346 22372 33358
rect 22316 33294 22318 33346
rect 22370 33294 22372 33346
rect 21980 33236 22036 33246
rect 21756 32722 21812 32732
rect 21868 33234 22036 33236
rect 21868 33182 21982 33234
rect 22034 33182 22036 33234
rect 21868 33180 22036 33182
rect 21644 32564 21700 32574
rect 21868 32564 21924 33180
rect 21980 33170 22036 33180
rect 22316 32900 22372 33294
rect 22540 33124 22596 33964
rect 22652 33954 22708 33964
rect 22652 33572 22708 33582
rect 22764 33572 22820 35532
rect 22876 35522 22932 35532
rect 22652 33570 22820 33572
rect 22652 33518 22654 33570
rect 22706 33518 22820 33570
rect 22652 33516 22820 33518
rect 22876 34916 22932 34926
rect 22652 33506 22708 33516
rect 22876 33348 22932 34860
rect 23324 34916 23380 39200
rect 24444 37268 24500 39200
rect 24332 37212 24500 37268
rect 24332 36596 24388 37212
rect 24522 36876 24786 36886
rect 24578 36820 24626 36876
rect 24682 36820 24730 36876
rect 24522 36810 24786 36820
rect 24332 36530 24388 36540
rect 23548 36482 23604 36494
rect 23548 36430 23550 36482
rect 23602 36430 23604 36482
rect 23548 35700 23604 36430
rect 24556 36454 24612 36466
rect 24556 36402 24558 36454
rect 24610 36402 24612 36454
rect 23940 36258 23996 36270
rect 23940 36206 23942 36258
rect 23994 36206 23996 36258
rect 23660 35700 23716 35710
rect 23548 35698 23716 35700
rect 23548 35646 23662 35698
rect 23714 35646 23716 35698
rect 23548 35644 23716 35646
rect 23660 35588 23716 35644
rect 23940 35588 23996 36206
rect 24556 35924 24612 36402
rect 24556 35858 24612 35868
rect 24332 35812 24388 35822
rect 24052 35588 24108 35598
rect 23660 35586 24108 35588
rect 23660 35534 24054 35586
rect 24106 35534 24108 35586
rect 23660 35532 24108 35534
rect 24052 35140 24108 35532
rect 24052 35074 24108 35084
rect 24332 35138 24388 35756
rect 25228 35725 25284 35738
rect 24780 35700 24836 35710
rect 25228 35700 25230 35725
rect 25282 35700 25284 35725
rect 24780 35698 25172 35700
rect 24780 35646 24782 35698
rect 24834 35646 25172 35698
rect 24780 35644 25172 35646
rect 24780 35634 24836 35644
rect 24444 35476 24500 35514
rect 24444 35410 24500 35420
rect 24522 35308 24786 35318
rect 24578 35252 24626 35308
rect 24682 35252 24730 35308
rect 24522 35242 24786 35252
rect 24332 35086 24334 35138
rect 24386 35086 24388 35138
rect 24332 35074 24388 35086
rect 24892 35140 24948 35150
rect 23324 34850 23380 34860
rect 23996 34914 24052 34926
rect 23996 34862 23998 34914
rect 24050 34862 24052 34914
rect 23996 33796 24052 34862
rect 24892 34916 24948 35084
rect 25004 34916 25060 34926
rect 24892 34914 25060 34916
rect 24892 34862 25006 34914
rect 25058 34862 25060 34914
rect 24892 34860 25060 34862
rect 24556 34018 24612 34030
rect 24556 33966 24558 34018
rect 24610 33966 24612 34018
rect 24556 33908 24612 33966
rect 23996 33730 24052 33740
rect 24108 33852 24612 33908
rect 22988 33348 23044 33358
rect 22876 33346 23044 33348
rect 22876 33294 22990 33346
rect 23042 33294 23044 33346
rect 22876 33292 23044 33294
rect 22988 33282 23044 33292
rect 23996 33236 24052 33246
rect 23156 33124 23212 33134
rect 22540 33068 23044 33124
rect 21644 32562 21924 32564
rect 21644 32510 21646 32562
rect 21698 32510 21924 32562
rect 21644 32508 21924 32510
rect 21980 32844 22372 32900
rect 21644 32498 21700 32508
rect 21980 32350 22036 32844
rect 22988 32674 23044 33068
rect 22596 32618 22652 32630
rect 22596 32566 22598 32618
rect 22650 32566 22652 32618
rect 22988 32622 22990 32674
rect 23042 32622 23044 32674
rect 22988 32610 23044 32622
rect 23156 32618 23212 33068
rect 22596 32564 22652 32566
rect 22596 32508 22708 32564
rect 21924 32338 22036 32350
rect 21924 32286 21926 32338
rect 21978 32286 22036 32338
rect 21924 32284 22036 32286
rect 21924 32274 21980 32284
rect 21532 31938 21588 31948
rect 21756 32228 21812 32238
rect 21756 31118 21812 32172
rect 22372 32004 22428 32014
rect 22652 32004 22708 32508
rect 22764 32562 22820 32574
rect 22764 32510 22766 32562
rect 22818 32510 22820 32562
rect 23156 32566 23158 32618
rect 23210 32566 23212 32618
rect 23324 33122 23380 33134
rect 23324 33070 23326 33122
rect 23378 33070 23380 33122
rect 23324 32676 23380 33070
rect 23324 32610 23380 32620
rect 23996 33012 24052 33180
rect 23156 32554 23212 32566
rect 23660 32562 23716 32574
rect 22764 32228 22820 32510
rect 23660 32510 23662 32562
rect 23714 32510 23716 32562
rect 23660 32452 23716 32510
rect 23660 32386 23716 32396
rect 22764 32162 22820 32172
rect 23100 32340 23156 32350
rect 23492 32340 23548 32350
rect 22764 32004 22820 32014
rect 22652 32002 22820 32004
rect 22652 31950 22766 32002
rect 22818 31950 22820 32002
rect 22652 31948 22820 31950
rect 22092 31778 22148 31790
rect 22092 31726 22094 31778
rect 22146 31726 22148 31778
rect 22092 31668 22148 31726
rect 22092 31602 22148 31612
rect 22204 31778 22260 31790
rect 22204 31726 22206 31778
rect 22258 31726 22260 31778
rect 20972 31042 21028 31052
rect 21700 31106 21812 31118
rect 21700 31054 21702 31106
rect 21754 31054 21812 31106
rect 21700 31052 21812 31054
rect 21700 31042 21756 31052
rect 20188 30996 20244 31006
rect 20412 30968 20916 31024
rect 20188 30548 20244 30940
rect 20468 30772 20524 30782
rect 20188 30482 20244 30492
rect 20300 30770 20524 30772
rect 20300 30718 20470 30770
rect 20522 30718 20524 30770
rect 20300 30716 20524 30718
rect 20188 30212 20244 30222
rect 20188 30118 20244 30156
rect 20300 30212 20356 30716
rect 20468 30706 20524 30716
rect 20636 30548 20692 30558
rect 20412 30212 20468 30222
rect 20300 30210 20412 30212
rect 20300 30158 20302 30210
rect 20354 30158 20412 30210
rect 20300 30156 20412 30158
rect 20300 30146 20356 30156
rect 20412 30146 20468 30156
rect 20076 29932 20244 29988
rect 19860 29820 20124 29830
rect 19916 29764 19964 29820
rect 20020 29764 20068 29820
rect 19860 29754 20124 29764
rect 20188 29652 20244 29932
rect 20076 29596 20244 29652
rect 19908 29540 19964 29550
rect 19908 29446 19964 29484
rect 19870 28868 19926 28878
rect 20076 28868 20132 29596
rect 20524 29428 20580 29438
rect 19870 28866 20132 28868
rect 19870 28814 19872 28866
rect 19924 28814 20132 28866
rect 19870 28812 20132 28814
rect 20412 29426 20580 29428
rect 20412 29374 20526 29426
rect 20578 29374 20580 29426
rect 20412 29372 20580 29374
rect 19870 28802 19926 28812
rect 20412 28644 20468 29372
rect 20524 29362 20580 29372
rect 20412 28550 20468 28588
rect 20524 28810 20580 28822
rect 20524 28758 20526 28810
rect 20578 28758 20580 28810
rect 19860 28252 20124 28262
rect 19916 28196 19964 28252
rect 20020 28196 20068 28252
rect 19860 28186 20124 28196
rect 19740 27794 19796 27804
rect 20076 27972 20132 27982
rect 20076 27858 20132 27916
rect 20334 27895 20390 27907
rect 20076 27806 20078 27858
rect 20130 27806 20132 27858
rect 17724 27246 17726 27298
rect 17778 27246 17780 27298
rect 17724 27234 17780 27246
rect 18564 27298 18620 27580
rect 19628 27570 19684 27580
rect 18564 27246 18566 27298
rect 18618 27246 18620 27298
rect 18564 27234 18620 27246
rect 19292 27412 19348 27422
rect 17388 27022 17390 27074
rect 17442 27022 17444 27074
rect 17388 26964 17444 27022
rect 18844 27076 18900 27086
rect 18844 26982 18900 27020
rect 19068 27074 19124 27086
rect 19068 27022 19070 27074
rect 19122 27022 19124 27074
rect 17388 26898 17444 26908
rect 17948 26964 18004 26974
rect 17276 26292 17332 26302
rect 17276 26198 17332 26236
rect 17612 26068 17668 26078
rect 17388 26066 17668 26068
rect 17388 26014 17614 26066
rect 17666 26014 17668 26066
rect 17388 26012 17668 26014
rect 17388 23940 17444 26012
rect 17612 26002 17668 26012
rect 17612 25844 17668 25854
rect 17612 24766 17668 25788
rect 17612 24714 17614 24766
rect 17666 24714 17668 24766
rect 17612 24702 17668 24714
rect 17836 24724 17892 24734
rect 17500 24612 17556 24622
rect 17500 24610 17724 24612
rect 17500 24558 17502 24610
rect 17554 24558 17724 24610
rect 17500 24556 17724 24558
rect 17500 24546 17556 24556
rect 17668 23994 17724 24556
rect 17500 23940 17556 23950
rect 17388 23884 17500 23940
rect 17668 23942 17670 23994
rect 17722 23942 17724 23994
rect 17668 23930 17724 23942
rect 17500 23846 17556 23884
rect 17836 23716 17892 24668
rect 17836 23650 17892 23660
rect 17164 23314 17220 23324
rect 17948 23380 18004 26908
rect 19068 26964 19124 27022
rect 19292 27074 19348 27356
rect 19964 27188 20020 27198
rect 19852 27186 20020 27188
rect 19852 27134 19966 27186
rect 20018 27134 20020 27186
rect 19852 27132 20020 27134
rect 19292 27022 19294 27074
rect 19346 27022 19348 27074
rect 19292 27010 19348 27022
rect 19404 27074 19460 27086
rect 19404 27022 19406 27074
rect 19458 27022 19460 27074
rect 19404 26908 19460 27022
rect 19516 27076 19628 27132
rect 19572 27074 19628 27076
rect 19624 27022 19628 27074
rect 19572 27020 19628 27022
rect 19516 27010 19626 27020
rect 19068 26898 19124 26908
rect 19180 26852 19236 26862
rect 18732 26292 18788 26302
rect 18620 25508 18676 25518
rect 18620 25414 18676 25452
rect 18116 25282 18172 25294
rect 18116 25230 18118 25282
rect 18170 25230 18172 25282
rect 18116 24724 18172 25230
rect 18452 25284 18508 25294
rect 18452 25190 18508 25228
rect 18732 24948 18788 26236
rect 19180 25956 19236 26796
rect 19180 25890 19236 25900
rect 19292 26852 19460 26908
rect 19852 26852 19908 27132
rect 19964 27122 20020 27132
rect 19292 25732 19348 26852
rect 19740 26796 19908 26852
rect 20076 26852 20132 27806
rect 20188 27860 20244 27870
rect 20188 27766 20244 27804
rect 20334 27843 20336 27895
rect 20388 27843 20390 27895
rect 20334 27412 20390 27843
rect 20300 27356 20390 27412
rect 20076 26796 20244 26852
rect 19572 26628 19628 26638
rect 19572 26346 19628 26572
rect 19404 26290 19460 26302
rect 19404 26238 19406 26290
rect 19458 26238 19460 26290
rect 19572 26294 19574 26346
rect 19626 26294 19628 26346
rect 19572 26282 19628 26294
rect 19404 26180 19460 26238
rect 19404 26124 19684 26180
rect 19516 25956 19572 25966
rect 19292 25666 19348 25676
rect 19404 25844 19460 25854
rect 18956 25620 19012 25630
rect 18508 24892 18788 24948
rect 18844 25618 19012 25620
rect 18844 25566 18958 25618
rect 19010 25566 19012 25618
rect 18844 25564 19012 25566
rect 18284 24836 18340 24846
rect 18284 24778 18340 24780
rect 18284 24726 18286 24778
rect 18338 24726 18340 24778
rect 18284 24714 18340 24726
rect 18396 24750 18452 24762
rect 18116 24658 18172 24668
rect 18396 24698 18398 24750
rect 18450 24698 18452 24750
rect 18396 24174 18452 24698
rect 18508 24276 18564 24892
rect 18844 24778 18900 25564
rect 18956 25554 19012 25564
rect 19404 25518 19460 25788
rect 19350 25506 19460 25518
rect 19350 25454 19352 25506
rect 19404 25454 19460 25506
rect 19350 25452 19460 25454
rect 19516 25506 19572 25900
rect 19516 25454 19518 25506
rect 19570 25454 19572 25506
rect 19350 25442 19406 25452
rect 19516 25442 19572 25454
rect 19628 25506 19684 26124
rect 19628 25454 19630 25506
rect 19682 25454 19684 25506
rect 18676 24757 18732 24769
rect 18676 24705 18678 24757
rect 18730 24724 18732 24757
rect 18844 24726 18846 24778
rect 18898 24726 18900 24778
rect 18730 24705 18788 24724
rect 18844 24714 18900 24726
rect 18956 25284 19012 25294
rect 18676 24668 18788 24705
rect 18508 24220 18676 24276
rect 18396 24162 18470 24174
rect 18396 24110 18416 24162
rect 18468 24110 18470 24162
rect 18396 24108 18470 24110
rect 18414 24098 18470 24108
rect 17948 23314 18004 23324
rect 18172 23938 18228 23950
rect 18172 23886 18174 23938
rect 18226 23886 18228 23938
rect 18060 23268 18116 23278
rect 17948 23154 18004 23166
rect 17948 23102 17950 23154
rect 18002 23102 18004 23154
rect 17164 19348 17220 19358
rect 17164 19254 17220 19292
rect 17500 19236 17556 19246
rect 17276 18450 17332 18462
rect 17276 18398 17278 18450
rect 17330 18398 17332 18450
rect 17276 16436 17332 18398
rect 17500 17118 17556 19180
rect 17780 19236 17836 19246
rect 17780 19142 17836 19180
rect 17948 18452 18004 23102
rect 18060 23154 18116 23212
rect 18060 23102 18062 23154
rect 18114 23102 18116 23154
rect 18060 23090 18116 23102
rect 18172 21812 18228 23886
rect 18340 23604 18396 23614
rect 18340 23266 18396 23548
rect 18340 23214 18342 23266
rect 18394 23214 18396 23266
rect 18340 23202 18396 23214
rect 18620 22372 18676 24220
rect 18732 23278 18788 24668
rect 18956 24612 19012 25228
rect 19292 25284 19348 25294
rect 18956 24556 19068 24612
rect 19012 23994 19068 24556
rect 19124 24500 19180 24510
rect 19124 24406 19180 24444
rect 18844 23938 18900 23950
rect 18844 23886 18846 23938
rect 18898 23886 18900 23938
rect 19012 23942 19014 23994
rect 19066 23942 19068 23994
rect 19012 23930 19068 23942
rect 19180 23940 19236 23950
rect 18844 23604 18900 23886
rect 19180 23846 19236 23884
rect 19292 23938 19348 25228
rect 19628 25060 19684 25454
rect 19292 23886 19294 23938
rect 19346 23886 19348 23938
rect 19292 23874 19348 23886
rect 19404 25004 19684 25060
rect 19404 23940 19460 25004
rect 19740 24948 19796 26796
rect 19860 26684 20124 26694
rect 19916 26628 19964 26684
rect 20020 26628 20068 26684
rect 19860 26618 20124 26628
rect 19852 26404 19908 26414
rect 19852 25284 19908 26348
rect 20076 26292 20132 26302
rect 20076 26198 20132 26236
rect 20076 25732 20132 25742
rect 20188 25732 20244 26796
rect 20300 26628 20356 27356
rect 20524 26852 20580 28758
rect 20636 28642 20692 30492
rect 20748 30436 20804 30446
rect 20748 29482 20804 30380
rect 20748 29430 20750 29482
rect 20802 29430 20804 29482
rect 20860 29540 20916 30968
rect 21196 30994 21252 31006
rect 21196 30942 21198 30994
rect 21250 30942 21252 30994
rect 21028 30882 21084 30894
rect 21028 30830 21030 30882
rect 21082 30830 21084 30882
rect 21028 30772 21084 30830
rect 21028 30706 21084 30716
rect 21196 29876 21252 30942
rect 21420 30994 21476 31006
rect 21420 30942 21422 30994
rect 21474 30942 21476 30994
rect 21420 30660 21476 30942
rect 21420 30594 21476 30604
rect 21532 30548 21588 30558
rect 20860 29474 20916 29484
rect 20972 29820 21196 29876
rect 20748 29418 20804 29430
rect 20860 29316 20916 29326
rect 20860 29222 20916 29260
rect 20636 28590 20638 28642
rect 20690 28590 20692 28642
rect 20636 28578 20692 28590
rect 20972 28084 21028 29820
rect 21196 29810 21252 29820
rect 21308 30210 21364 30222
rect 21308 30158 21310 30210
rect 21362 30158 21364 30210
rect 20972 28018 21028 28028
rect 21084 29540 21140 29550
rect 21084 28756 21140 29484
rect 21196 29428 21252 29438
rect 21196 29334 21252 29372
rect 20524 26786 20580 26796
rect 20636 27860 20692 27870
rect 20300 26562 20356 26572
rect 20318 26404 20374 26414
rect 20524 26404 20580 26414
rect 20318 26402 20524 26404
rect 20318 26350 20320 26402
rect 20372 26350 20524 26402
rect 20318 26348 20524 26350
rect 20318 26338 20374 26348
rect 20524 26338 20580 26348
rect 20636 26180 20692 27804
rect 21084 27860 21140 28700
rect 21308 27972 21364 30158
rect 21420 30212 21476 30222
rect 21420 30118 21476 30156
rect 21532 29428 21588 30492
rect 22204 30446 22260 31726
rect 22372 31778 22428 31948
rect 22764 31938 22820 31948
rect 22372 31726 22374 31778
rect 22426 31726 22428 31778
rect 22372 31714 22428 31726
rect 22652 31780 22708 31790
rect 21700 30436 21756 30446
rect 21700 30210 21756 30380
rect 22148 30434 22260 30446
rect 22148 30382 22150 30434
rect 22202 30382 22260 30434
rect 22148 30380 22260 30382
rect 22316 31556 22372 31566
rect 22316 30994 22372 31500
rect 22652 30996 22708 31724
rect 22876 31033 22932 31045
rect 22876 31024 22878 31033
rect 22316 30942 22318 30994
rect 22370 30942 22372 30994
rect 22148 30370 22204 30380
rect 21700 30158 21702 30210
rect 21754 30158 21756 30210
rect 21700 30146 21756 30158
rect 22316 30212 22372 30942
rect 22540 30994 22708 30996
rect 22540 30942 22654 30994
rect 22706 30942 22708 30994
rect 22540 30940 22708 30942
rect 22540 30436 22596 30940
rect 22652 30930 22708 30940
rect 22764 30996 22878 31024
rect 22930 30996 22932 31033
rect 22764 30968 22876 30996
rect 22428 30212 22484 30222
rect 22316 30210 22484 30212
rect 22316 30158 22430 30210
rect 22482 30158 22484 30210
rect 22316 30156 22484 30158
rect 21644 29428 21700 29438
rect 21532 29426 21700 29428
rect 21532 29374 21646 29426
rect 21698 29374 21700 29426
rect 21532 29372 21700 29374
rect 21644 29362 21700 29372
rect 22316 29426 22372 30156
rect 22428 30146 22484 30156
rect 22540 30210 22596 30380
rect 22540 30158 22542 30210
rect 22594 30158 22596 30210
rect 22764 30166 22820 30968
rect 22876 30892 22932 30940
rect 22988 30882 23044 30894
rect 22988 30830 22990 30882
rect 23042 30830 23044 30882
rect 22988 30324 23044 30830
rect 22988 30258 23044 30268
rect 22540 30146 22596 30158
rect 22708 30154 22820 30166
rect 22708 30102 22710 30154
rect 22762 30102 22820 30154
rect 22708 29988 22820 30102
rect 22876 30210 22932 30222
rect 22876 30158 22878 30210
rect 22930 30158 22932 30210
rect 22876 30100 22932 30158
rect 23100 30100 23156 32284
rect 23324 32338 23548 32340
rect 23324 32286 23494 32338
rect 23546 32286 23548 32338
rect 23324 32284 23548 32286
rect 23324 32004 23380 32284
rect 23492 32274 23548 32284
rect 23324 30994 23380 31948
rect 23996 32004 24052 32956
rect 24108 32452 24164 33852
rect 24522 33740 24786 33750
rect 24578 33684 24626 33740
rect 24682 33684 24730 33740
rect 24522 33674 24786 33684
rect 24276 33236 24332 33246
rect 24276 33142 24332 33180
rect 24724 33124 24780 33134
rect 24892 33124 24948 34860
rect 25004 34850 25060 34860
rect 25116 33796 25172 35644
rect 25228 35634 25284 35644
rect 25564 35140 25620 39200
rect 25900 36258 25956 36270
rect 25900 36206 25902 36258
rect 25954 36206 25956 36258
rect 25788 35476 25844 35486
rect 25564 35074 25620 35084
rect 25676 35252 25732 35262
rect 25116 33730 25172 33740
rect 25564 34018 25620 34030
rect 25564 33966 25566 34018
rect 25618 33966 25620 34018
rect 25116 33460 25172 33470
rect 24444 33122 24948 33124
rect 24444 33070 24726 33122
rect 24778 33070 24948 33122
rect 24444 33068 24948 33070
rect 24444 32900 24500 33068
rect 24724 33058 24780 33068
rect 24276 32844 24500 32900
rect 24276 32786 24332 32844
rect 24276 32734 24278 32786
rect 24330 32734 24332 32786
rect 24276 32722 24332 32734
rect 24612 32730 24668 32742
rect 24612 32678 24614 32730
rect 24666 32678 24668 32730
rect 24612 32564 24668 32678
rect 24612 32498 24668 32508
rect 24780 32676 24836 32686
rect 24780 32562 24836 32620
rect 24780 32510 24782 32562
rect 24834 32510 24836 32562
rect 24780 32498 24836 32510
rect 24108 32386 24164 32396
rect 24332 32452 24388 32462
rect 23996 31938 24052 31948
rect 24220 31890 24276 31902
rect 24220 31838 24222 31890
rect 24274 31838 24276 31890
rect 23436 31778 23492 31790
rect 23436 31726 23438 31778
rect 23490 31726 23492 31778
rect 23436 31556 23492 31726
rect 23772 31780 23828 31790
rect 23772 31686 23828 31724
rect 24108 31722 24164 31734
rect 23436 31490 23492 31500
rect 24108 31670 24110 31722
rect 24162 31670 24164 31722
rect 23324 30942 23326 30994
rect 23378 30942 23380 30994
rect 23324 30930 23380 30942
rect 23660 31108 23716 31118
rect 22876 30044 23268 30100
rect 22708 29932 22932 29988
rect 22316 29374 22318 29426
rect 22370 29374 22372 29426
rect 22316 29362 22372 29374
rect 22708 29428 22764 29438
rect 21532 29258 21588 29270
rect 21532 29206 21534 29258
rect 21586 29206 21588 29258
rect 21532 28868 21588 29206
rect 22708 29258 22764 29372
rect 22708 29206 22710 29258
rect 22762 29206 22764 29258
rect 22708 29194 22764 29206
rect 22876 29426 22932 29932
rect 22876 29374 22878 29426
rect 22930 29374 22932 29426
rect 22876 29092 22932 29374
rect 21532 28802 21588 28812
rect 21700 29036 22932 29092
rect 21700 28698 21756 29036
rect 23100 28980 23156 28990
rect 22260 28868 22316 28878
rect 22260 28774 22316 28812
rect 21532 28644 21588 28654
rect 21308 27906 21364 27916
rect 21420 28642 21588 28644
rect 21420 28590 21534 28642
rect 21586 28590 21588 28642
rect 21700 28646 21702 28698
rect 21754 28646 21756 28698
rect 22764 28756 22820 28766
rect 22764 28662 22820 28700
rect 21700 28634 21756 28646
rect 21980 28642 22036 28654
rect 21420 28588 21588 28590
rect 21196 27860 21252 27870
rect 21084 27858 21252 27860
rect 21084 27806 21198 27858
rect 21250 27806 21252 27858
rect 21084 27804 21252 27806
rect 20748 27748 20804 27758
rect 20748 27654 20804 27692
rect 21084 27188 21140 27804
rect 21196 27794 21252 27804
rect 21420 27412 21476 28588
rect 21532 28578 21588 28588
rect 21980 28590 21982 28642
rect 22034 28590 22036 28642
rect 21868 28532 21924 28542
rect 21868 28438 21924 28476
rect 21980 28308 22036 28590
rect 23100 28642 23156 28924
rect 23100 28590 23102 28642
rect 23154 28590 23156 28642
rect 21644 28252 22036 28308
rect 22148 28420 22204 28430
rect 21532 27858 21588 27870
rect 21532 27806 21534 27858
rect 21586 27806 21588 27858
rect 21532 27748 21588 27806
rect 21532 27682 21588 27692
rect 21644 27690 21700 28252
rect 21644 27638 21646 27690
rect 21698 27638 21700 27690
rect 21644 27626 21700 27638
rect 21756 28084 21812 28094
rect 21084 27122 21140 27132
rect 21196 27356 21476 27412
rect 21644 27524 21700 27534
rect 20804 27076 20860 27086
rect 20804 26982 20860 27020
rect 21196 26458 21252 27356
rect 20748 26404 20804 26414
rect 21196 26406 21198 26458
rect 21250 26406 21252 26458
rect 21196 26394 21252 26406
rect 21308 27242 21364 27254
rect 21308 27190 21310 27242
rect 21362 27190 21364 27242
rect 20748 26292 20804 26348
rect 21028 26319 21084 26331
rect 21028 26292 21030 26319
rect 20748 26267 21030 26292
rect 21082 26267 21084 26319
rect 20748 26236 21084 26267
rect 21308 26290 21364 27190
rect 21420 27188 21476 27198
rect 21420 27074 21476 27132
rect 21420 27022 21422 27074
rect 21474 27022 21476 27074
rect 21420 27010 21476 27022
rect 21644 27076 21700 27468
rect 21308 26238 21310 26290
rect 21362 26238 21364 26290
rect 21308 26226 21364 26238
rect 20076 25730 20244 25732
rect 20076 25678 20078 25730
rect 20130 25678 20244 25730
rect 20076 25676 20244 25678
rect 20076 25508 20132 25676
rect 20076 25442 20132 25452
rect 19852 25218 19908 25228
rect 19860 25116 20124 25126
rect 19916 25060 19964 25116
rect 20020 25060 20068 25116
rect 19860 25050 20124 25060
rect 19740 24892 20132 24948
rect 19516 24836 19572 24846
rect 19516 24778 19572 24780
rect 19516 24726 19518 24778
rect 19570 24726 19572 24778
rect 20076 24778 20132 24892
rect 19516 24714 19572 24726
rect 19628 24750 19684 24762
rect 19628 24698 19630 24750
rect 19682 24698 19684 24750
rect 19908 24757 19964 24769
rect 19628 24174 19684 24698
rect 19572 24162 19684 24174
rect 19572 24110 19574 24162
rect 19626 24110 19684 24162
rect 19572 24108 19684 24110
rect 19740 24724 19796 24734
rect 19908 24705 19910 24757
rect 19962 24724 19964 24757
rect 20076 24726 20078 24778
rect 20130 24726 20132 24778
rect 19962 24705 20020 24724
rect 20076 24714 20132 24726
rect 19908 24668 20020 24705
rect 19572 24098 19628 24108
rect 19404 23874 19460 23884
rect 18844 23538 18900 23548
rect 18956 23828 19012 23838
rect 18732 23266 18844 23278
rect 18732 23214 18790 23266
rect 18842 23214 18844 23266
rect 18732 23212 18844 23214
rect 18788 23202 18844 23212
rect 18732 22484 18788 22494
rect 18732 22390 18788 22428
rect 18060 21756 18228 21812
rect 18340 22316 18676 22372
rect 18340 21810 18396 22316
rect 18340 21758 18342 21810
rect 18394 21758 18396 21810
rect 18060 18564 18116 21756
rect 18340 21746 18396 21758
rect 18172 21586 18228 21598
rect 18172 21534 18174 21586
rect 18226 21534 18228 21586
rect 18172 19348 18228 21534
rect 18956 20132 19012 23772
rect 19292 23716 19348 23726
rect 19068 23156 19124 23166
rect 19068 21810 19124 23100
rect 19292 23156 19348 23660
rect 19740 23380 19796 24668
rect 19964 24174 20020 24668
rect 20188 24500 20244 25676
rect 20524 26124 20692 26180
rect 20412 25506 20468 25518
rect 20412 25454 20414 25506
rect 20466 25454 20468 25506
rect 20412 25284 20468 25454
rect 20524 25506 20580 26124
rect 20692 25732 20748 25742
rect 20692 25638 20748 25676
rect 20524 25454 20526 25506
rect 20578 25454 20580 25506
rect 20524 25396 20580 25454
rect 20524 25330 20580 25340
rect 20412 25218 20468 25228
rect 21476 25284 21532 25294
rect 21476 25190 21532 25228
rect 20356 24724 20412 24734
rect 20636 24724 20692 24734
rect 20356 24722 20692 24724
rect 20356 24670 20358 24722
rect 20410 24670 20638 24722
rect 20690 24670 20692 24722
rect 20356 24668 20692 24670
rect 20356 24658 20412 24668
rect 20636 24658 20692 24668
rect 21308 24724 21364 24734
rect 20972 24612 21028 24622
rect 20972 24518 21028 24556
rect 20524 24500 20580 24510
rect 20188 24444 20468 24500
rect 19964 24162 20076 24174
rect 19964 24110 20022 24162
rect 20074 24110 20076 24162
rect 19964 24108 20076 24110
rect 20020 24098 20076 24108
rect 20300 23938 20356 23950
rect 20300 23886 20302 23938
rect 20354 23886 20356 23938
rect 19860 23548 20124 23558
rect 19916 23492 19964 23548
rect 20020 23492 20068 23548
rect 19860 23482 20124 23492
rect 19740 23324 20020 23380
rect 19292 23154 19460 23156
rect 19292 23102 19294 23154
rect 19346 23102 19460 23154
rect 19292 23100 19460 23102
rect 19292 23090 19348 23100
rect 19404 22494 19460 23100
rect 19740 23154 19796 23166
rect 19740 23102 19742 23154
rect 19794 23102 19796 23154
rect 19404 22482 19516 22494
rect 19404 22430 19462 22482
rect 19514 22430 19516 22482
rect 19404 22428 19516 22430
rect 19460 22418 19516 22428
rect 19068 21758 19070 21810
rect 19122 21758 19124 21810
rect 19068 21746 19124 21758
rect 19628 22372 19684 22382
rect 19740 22372 19796 23102
rect 19964 22594 20020 23324
rect 20076 23268 20132 23278
rect 20076 23174 20132 23212
rect 20300 23156 20356 23886
rect 20412 23938 20468 24444
rect 20412 23886 20414 23938
rect 20466 23886 20468 23938
rect 20412 23874 20468 23886
rect 20300 23090 20356 23100
rect 20412 23156 20468 23166
rect 20524 23156 20580 24444
rect 20748 23940 20804 23950
rect 20748 23378 20804 23884
rect 21196 23940 21252 23950
rect 21308 23940 21364 24668
rect 21196 23938 21364 23940
rect 21196 23886 21198 23938
rect 21250 23886 21364 23938
rect 21196 23884 21364 23886
rect 21196 23874 21252 23884
rect 20748 23326 20750 23378
rect 20802 23326 20804 23378
rect 20748 23314 20804 23326
rect 20412 23154 20580 23156
rect 20412 23102 20414 23154
rect 20466 23102 20580 23154
rect 20412 23100 20580 23102
rect 20412 23090 20468 23100
rect 19964 22542 19966 22594
rect 20018 22542 20020 22594
rect 19964 22530 20020 22542
rect 19628 22370 19796 22372
rect 19628 22318 19630 22370
rect 19682 22318 19796 22370
rect 19628 22316 19796 22318
rect 19404 21588 19460 21598
rect 19292 21532 19404 21588
rect 19068 20804 19124 20814
rect 19068 20802 19236 20804
rect 19068 20750 19070 20802
rect 19122 20750 19236 20802
rect 19068 20748 19236 20750
rect 19068 20738 19124 20748
rect 18956 20066 19012 20076
rect 18172 19282 18228 19292
rect 18844 19234 18900 19246
rect 18844 19182 18846 19234
rect 18898 19182 18900 19234
rect 18844 18676 18900 19182
rect 18844 18610 18900 18620
rect 19068 19178 19124 19190
rect 19068 19126 19070 19178
rect 19122 19126 19124 19178
rect 19068 18676 19124 19126
rect 19068 18610 19124 18620
rect 18060 18508 18228 18564
rect 17724 18396 18004 18452
rect 17500 17106 17612 17118
rect 17500 17054 17558 17106
rect 17610 17054 17612 17106
rect 17500 17052 17612 17054
rect 17556 17042 17612 17052
rect 17724 16996 17780 18396
rect 18060 18340 18116 18350
rect 17836 18338 18116 18340
rect 17836 18286 18062 18338
rect 18114 18286 18116 18338
rect 17836 18284 18116 18286
rect 17836 17890 17892 18284
rect 18060 18274 18116 18284
rect 17836 17838 17838 17890
rect 17890 17838 17892 17890
rect 17836 17826 17892 17838
rect 18172 17892 18228 18508
rect 19180 18340 19236 20748
rect 19180 18274 19236 18284
rect 19292 18116 19348 21532
rect 19404 21494 19460 21532
rect 19404 21028 19460 21038
rect 19404 20934 19460 20972
rect 19516 19236 19572 19246
rect 19516 19142 19572 19180
rect 19404 19066 19460 19078
rect 19404 19014 19406 19066
rect 19458 19014 19460 19066
rect 19404 19012 19460 19014
rect 19628 19012 19684 22316
rect 19860 21980 20124 21990
rect 19916 21924 19964 21980
rect 20020 21924 20068 21980
rect 19860 21914 20124 21924
rect 21644 21812 21700 27020
rect 21756 25284 21812 28028
rect 22148 28082 22204 28364
rect 23100 28420 23156 28590
rect 23100 28354 23156 28364
rect 22148 28030 22150 28082
rect 22202 28030 22204 28082
rect 22148 28018 22204 28030
rect 23212 26628 23268 30044
rect 23548 29988 23604 29998
rect 23436 29426 23492 29438
rect 23436 29374 23438 29426
rect 23490 29374 23492 29426
rect 23436 28868 23492 29374
rect 23436 28802 23492 28812
rect 23548 28644 23604 29932
rect 23548 28578 23604 28588
rect 23660 28756 23716 31052
rect 23772 30996 23828 31006
rect 23772 30902 23828 30940
rect 24108 30996 24164 31670
rect 24108 30902 24164 30940
rect 23996 30772 24052 30782
rect 23772 30212 23828 30222
rect 23772 30118 23828 30156
rect 23772 29652 23828 29662
rect 23772 29558 23828 29596
rect 23492 28420 23548 28430
rect 23492 28326 23548 28364
rect 23660 27860 23716 28700
rect 23884 27860 23940 27870
rect 21756 25218 21812 25228
rect 22204 26068 22260 26078
rect 22092 24612 22148 24622
rect 22092 24518 22148 24556
rect 21980 23940 22036 23950
rect 21980 23846 22036 23884
rect 21532 21756 21700 21812
rect 19796 21588 19852 21598
rect 19796 21494 19852 21532
rect 21532 21028 21588 21756
rect 21644 21588 21700 21598
rect 21644 21494 21700 21532
rect 21980 21364 22036 21374
rect 21980 21270 22036 21308
rect 21532 20962 21588 20972
rect 22092 21028 22148 21038
rect 22204 21028 22260 26012
rect 22316 23380 22372 23390
rect 22316 22986 22372 23324
rect 23212 23268 23268 26572
rect 23548 27858 23940 27860
rect 23548 27806 23886 27858
rect 23938 27806 23940 27858
rect 23548 27804 23940 27806
rect 23548 25620 23604 27804
rect 23884 27794 23940 27804
rect 23996 27636 24052 30716
rect 24220 30660 24276 31838
rect 24332 31778 24388 32396
rect 24522 32172 24786 32182
rect 24578 32116 24626 32172
rect 24682 32116 24730 32172
rect 24522 32106 24786 32116
rect 24332 31726 24334 31778
rect 24386 31726 24388 31778
rect 24332 31714 24388 31726
rect 24724 30884 24780 30894
rect 24724 30790 24780 30828
rect 24220 30594 24276 30604
rect 24522 30604 24786 30614
rect 24578 30548 24626 30604
rect 24682 30548 24730 30604
rect 24522 30538 24786 30548
rect 24892 30548 24948 33068
rect 25004 33346 25060 33358
rect 25004 33294 25006 33346
rect 25058 33294 25060 33346
rect 25004 32340 25060 33294
rect 25116 33346 25172 33404
rect 25116 33294 25118 33346
rect 25170 33294 25172 33346
rect 25116 32676 25172 33294
rect 25282 33348 25338 33358
rect 25282 33254 25338 33292
rect 25116 32610 25172 32620
rect 25228 33124 25284 33134
rect 25004 32274 25060 32284
rect 25228 32002 25284 33068
rect 25564 32340 25620 33966
rect 25676 33570 25732 35196
rect 25788 35026 25844 35420
rect 25788 34974 25790 35026
rect 25842 34974 25844 35026
rect 25788 34962 25844 34974
rect 25900 35028 25956 36206
rect 26236 35474 26292 35486
rect 26236 35422 26238 35474
rect 26290 35422 26292 35474
rect 26236 35364 26292 35422
rect 25900 34962 25956 34972
rect 26012 35308 26292 35364
rect 26684 35364 26740 39200
rect 26012 34916 26068 35308
rect 26684 35298 26740 35308
rect 27244 36482 27300 36494
rect 27244 36430 27246 36482
rect 27298 36430 27300 36482
rect 27244 35252 27300 36430
rect 27244 35186 27300 35196
rect 27580 36258 27636 36270
rect 27580 36206 27582 36258
rect 27634 36206 27636 36258
rect 26012 34850 26068 34860
rect 27468 34132 27524 34142
rect 27580 34132 27636 36206
rect 27804 35252 27860 39200
rect 28588 36596 28644 36606
rect 28588 36482 28644 36540
rect 28588 36430 28590 36482
rect 28642 36430 28644 36482
rect 28588 36418 28644 36430
rect 28028 35725 28084 35737
rect 28028 35673 28030 35725
rect 28082 35673 28084 35725
rect 28028 35588 28084 35673
rect 28028 35522 28084 35532
rect 27804 35186 27860 35196
rect 28140 35476 28196 35486
rect 28028 34914 28084 34926
rect 28028 34862 28030 34914
rect 28082 34862 28084 34914
rect 27468 34130 27636 34132
rect 27468 34078 27470 34130
rect 27522 34078 27636 34130
rect 27468 34076 27636 34078
rect 27692 34802 27748 34814
rect 27692 34750 27694 34802
rect 27746 34750 27748 34802
rect 27468 34066 27524 34076
rect 25676 33518 25678 33570
rect 25730 33518 25732 33570
rect 25676 33506 25732 33518
rect 27244 33796 27300 33806
rect 26460 33318 26516 33330
rect 26460 33266 26462 33318
rect 26514 33266 26516 33318
rect 26292 33124 26348 33134
rect 26292 32676 26348 33068
rect 26292 32618 26348 32620
rect 25564 32274 25620 32284
rect 25676 32590 25732 32602
rect 25676 32538 25678 32590
rect 25730 32538 25732 32590
rect 25228 31950 25230 32002
rect 25282 31950 25284 32002
rect 25228 31938 25284 31950
rect 25564 31778 25620 31790
rect 25564 31726 25566 31778
rect 25618 31726 25620 31778
rect 25452 31108 25508 31118
rect 25452 30994 25508 31052
rect 25452 30942 25454 30994
rect 25506 30942 25508 30994
rect 25452 30930 25508 30942
rect 25564 30884 25620 31726
rect 25676 31780 25732 32538
rect 25900 32562 25956 32574
rect 25900 32510 25902 32562
rect 25954 32510 25956 32562
rect 26292 32566 26294 32618
rect 26346 32566 26348 32618
rect 26292 32554 26348 32566
rect 25676 31724 25844 31780
rect 25564 30818 25620 30828
rect 25676 30994 25732 31006
rect 25676 30942 25678 30994
rect 25730 30942 25732 30994
rect 24892 30482 24948 30492
rect 24668 30436 24724 30446
rect 24724 30380 24836 30436
rect 24668 30370 24724 30380
rect 23548 25554 23604 25564
rect 23660 27580 24052 27636
rect 24332 30212 24388 30222
rect 23212 23202 23268 23212
rect 23548 25396 23604 25406
rect 22428 23156 22484 23166
rect 22428 23062 22484 23100
rect 22764 23154 22820 23166
rect 22764 23102 22766 23154
rect 22818 23102 22820 23154
rect 22316 22934 22318 22986
rect 22370 22934 22372 22986
rect 22316 22922 22372 22934
rect 22652 21588 22708 21598
rect 22092 21026 22260 21028
rect 22092 20974 22094 21026
rect 22146 20974 22260 21026
rect 22092 20972 22260 20974
rect 22092 20962 22148 20972
rect 20188 20916 20244 20954
rect 20188 20850 20244 20860
rect 19852 20804 19908 20814
rect 19740 20802 19908 20804
rect 19740 20750 19854 20802
rect 19906 20750 19908 20802
rect 20524 20802 20580 20814
rect 19740 20748 19908 20750
rect 19740 20188 19796 20748
rect 19852 20738 19908 20748
rect 20300 20746 20356 20758
rect 20188 20692 20244 20702
rect 19860 20412 20124 20422
rect 19916 20356 19964 20412
rect 20020 20356 20068 20412
rect 19860 20346 20124 20356
rect 19908 20188 19964 20198
rect 19740 20186 19964 20188
rect 19740 20134 19910 20186
rect 19962 20134 19964 20186
rect 19740 20132 19964 20134
rect 19908 20066 19964 20076
rect 20076 20018 20132 20030
rect 20076 19966 20078 20018
rect 20130 19966 20132 20018
rect 19964 19236 20020 19246
rect 20076 19236 20132 19966
rect 20188 20020 20244 20636
rect 20300 20694 20302 20746
rect 20354 20694 20356 20746
rect 20300 20580 20356 20694
rect 20300 20514 20356 20524
rect 20524 20750 20526 20802
rect 20578 20750 20580 20802
rect 20188 19954 20244 19964
rect 20300 20053 20356 20065
rect 20300 20001 20302 20053
rect 20354 20001 20356 20053
rect 20300 19460 20356 20001
rect 20300 19394 20356 19404
rect 20412 20046 20468 20058
rect 20412 19994 20414 20046
rect 20466 19994 20468 20046
rect 20412 19236 20468 19994
rect 20524 19572 20580 20750
rect 21756 20804 21812 20814
rect 21420 20580 21476 20590
rect 20524 19506 20580 19516
rect 20636 20046 20692 20058
rect 20636 19994 20638 20046
rect 20690 19994 20692 20046
rect 19964 19234 20132 19236
rect 19964 19182 19966 19234
rect 20018 19182 20132 19234
rect 19964 19180 20132 19182
rect 20188 19180 20468 19236
rect 20524 19236 20580 19246
rect 20636 19236 20692 19994
rect 20910 20046 20966 20058
rect 20910 19994 20912 20046
rect 20964 20020 20966 20046
rect 21420 20020 21476 20524
rect 20964 19994 21364 20020
rect 20910 19964 21364 19994
rect 21140 19796 21196 19806
rect 21140 19702 21196 19740
rect 21308 19470 21364 19964
rect 21420 20018 21700 20020
rect 21420 19966 21422 20018
rect 21474 19966 21700 20018
rect 21420 19964 21700 19966
rect 21420 19954 21476 19964
rect 21308 19458 21420 19470
rect 21308 19406 21366 19458
rect 21418 19406 21420 19458
rect 21308 19404 21420 19406
rect 21364 19394 21420 19404
rect 20524 19234 20692 19236
rect 20524 19182 20526 19234
rect 20578 19182 20692 19234
rect 20524 19180 20692 19182
rect 21532 19234 21588 19246
rect 21532 19182 21534 19234
rect 21586 19182 21588 19234
rect 19404 18956 19684 19012
rect 19740 19124 19796 19134
rect 18172 17826 18228 17836
rect 19180 18060 19348 18116
rect 19404 18676 19460 18686
rect 18172 17668 18228 17678
rect 18172 17574 18228 17612
rect 17724 16930 17780 16940
rect 18396 17108 18452 17118
rect 17276 16370 17332 16380
rect 18060 16660 18116 16670
rect 18060 16100 18116 16604
rect 18396 16322 18452 17052
rect 18788 16882 18844 16894
rect 18788 16830 18790 16882
rect 18842 16830 18844 16882
rect 18788 16660 18844 16830
rect 18788 16594 18844 16604
rect 18396 16270 18398 16322
rect 18450 16270 18452 16322
rect 18396 16258 18452 16270
rect 17948 16098 18116 16100
rect 17948 16046 18062 16098
rect 18114 16046 18116 16098
rect 17948 16044 18116 16046
rect 17276 15314 17332 15326
rect 17276 15262 17278 15314
rect 17330 15262 17332 15314
rect 17276 13412 17332 15262
rect 17948 15148 18004 16044
rect 18060 16034 18116 16044
rect 18844 16212 18900 16222
rect 18844 16098 18900 16156
rect 18844 16046 18846 16098
rect 18898 16046 18900 16098
rect 18844 16034 18900 16046
rect 18060 15316 18116 15326
rect 18060 15222 18116 15260
rect 17724 15092 18004 15148
rect 17724 14644 17780 15092
rect 17724 14642 18004 14644
rect 17724 14590 17726 14642
rect 17778 14590 18004 14642
rect 17724 14588 18004 14590
rect 17724 14578 17780 14588
rect 17948 13982 18004 14588
rect 17948 13970 18060 13982
rect 17948 13918 18006 13970
rect 18058 13918 18060 13970
rect 17948 13916 18060 13918
rect 18004 13906 18060 13916
rect 17276 13346 17332 13356
rect 18172 13746 18228 13758
rect 18172 13694 18174 13746
rect 18226 13694 18228 13746
rect 18172 13412 18228 13694
rect 17724 12964 17780 12974
rect 17724 12870 17780 12908
rect 16492 11900 17108 11956
rect 15198 11788 15462 11798
rect 15254 11732 15302 11788
rect 15358 11732 15406 11788
rect 15198 11722 15462 11732
rect 16492 11396 16548 11406
rect 16268 11394 16548 11396
rect 16268 11342 16494 11394
rect 16546 11342 16548 11394
rect 16268 11340 16548 11342
rect 16268 10948 16324 11340
rect 16492 11330 16548 11340
rect 15820 10892 16324 10948
rect 15820 10834 15876 10892
rect 15820 10782 15822 10834
rect 15874 10782 15876 10834
rect 15820 10770 15876 10782
rect 15198 10220 15462 10230
rect 15254 10164 15302 10220
rect 15358 10164 15406 10220
rect 15198 10154 15462 10164
rect 15484 9940 15540 9950
rect 15484 9798 15540 9884
rect 15484 9746 15486 9798
rect 15538 9746 15540 9798
rect 15484 9268 15540 9746
rect 15484 9202 15540 9212
rect 15820 8818 15876 8830
rect 15820 8766 15822 8818
rect 15874 8766 15876 8818
rect 15198 8652 15462 8662
rect 15254 8596 15302 8652
rect 15358 8596 15406 8652
rect 15198 8586 15462 8596
rect 14980 8372 15092 8382
rect 14308 8370 15092 8372
rect 14308 8318 14982 8370
rect 15034 8318 15092 8370
rect 14308 8316 15092 8318
rect 14308 8314 14364 8316
rect 14308 8262 14310 8314
rect 14362 8262 14364 8314
rect 14980 8306 15036 8316
rect 14308 8250 14364 8262
rect 14476 8146 14532 8158
rect 14476 8094 14478 8146
rect 14530 8094 14532 8146
rect 14364 7476 14420 7486
rect 14140 7474 14420 7476
rect 14140 7422 14366 7474
rect 14418 7422 14420 7474
rect 14140 7420 14420 7422
rect 14364 7410 14420 7420
rect 12460 6738 12516 6748
rect 11116 6690 11284 6692
rect 11116 6638 11118 6690
rect 11170 6638 11284 6690
rect 11116 6636 11284 6638
rect 13804 6690 13860 6702
rect 13804 6638 13806 6690
rect 13858 6638 13860 6690
rect 11116 6626 11172 6636
rect 13562 6578 13618 6590
rect 13562 6526 13564 6578
rect 13616 6526 13618 6578
rect 12236 6468 12292 6478
rect 10686 6076 10948 6132
rect 11788 6466 12292 6468
rect 11788 6414 12238 6466
rect 12290 6414 12292 6466
rect 11788 6412 12292 6414
rect 10444 6020 10500 6030
rect 10444 5906 10500 5964
rect 10686 6018 10742 6076
rect 10686 5966 10688 6018
rect 10740 5966 10742 6018
rect 10686 5954 10742 5966
rect 10444 5854 10446 5906
rect 10498 5854 10500 5906
rect 10444 5842 10500 5854
rect 11004 5908 11060 5918
rect 11004 5124 11060 5852
rect 11788 5906 11844 6412
rect 12236 6402 12292 6412
rect 13562 6244 13618 6526
rect 11788 5854 11790 5906
rect 11842 5854 11844 5906
rect 11788 5842 11844 5854
rect 13468 6188 13618 6244
rect 11004 5030 11060 5068
rect 12572 5124 12628 5134
rect 10108 4956 10276 5012
rect 10108 4788 10164 4798
rect 10108 4365 10164 4732
rect 10108 4313 10110 4365
rect 10162 4313 10164 4365
rect 10108 4301 10164 4313
rect 9884 3554 10052 3556
rect 9884 3502 9886 3554
rect 9938 3502 10052 3554
rect 9884 3500 10052 3502
rect 10220 3526 10276 4956
rect 10332 4946 10388 4956
rect 11900 4898 11956 4910
rect 11900 4846 11902 4898
rect 11954 4846 11956 4898
rect 10536 4732 10800 4742
rect 10592 4676 10640 4732
rect 10696 4676 10744 4732
rect 10536 4666 10800 4676
rect 11900 4340 11956 4846
rect 11900 4274 11956 4284
rect 12572 4338 12628 5068
rect 13020 5124 13076 5134
rect 13020 5122 13188 5124
rect 13020 5070 13022 5122
rect 13074 5070 13188 5122
rect 13020 5068 13188 5070
rect 13020 5058 13076 5068
rect 12572 4286 12574 4338
rect 12626 4286 12628 4338
rect 12572 4274 12628 4286
rect 9884 3490 9940 3500
rect 10220 3474 10222 3526
rect 10274 3474 10276 3526
rect 10220 3462 10276 3474
rect 10892 4114 10948 4126
rect 10892 4062 10894 4114
rect 10946 4062 10948 4114
rect 10536 3164 10800 3174
rect 10592 3108 10640 3164
rect 10696 3108 10744 3164
rect 10536 3098 10800 3108
rect 10108 868 10164 878
rect 10108 800 10164 812
rect 10892 868 10948 4062
rect 13132 3790 13188 5068
rect 13356 4340 13412 4350
rect 13356 4246 13412 4284
rect 13132 3778 13244 3790
rect 13132 3726 13190 3778
rect 13242 3726 13244 3778
rect 13132 3724 13244 3726
rect 13188 3714 13244 3724
rect 13468 3554 13524 6188
rect 13692 6020 13748 6030
rect 13692 5926 13748 5964
rect 13580 5684 13636 5694
rect 13580 3780 13636 5628
rect 13804 4564 13860 6638
rect 14308 6634 14364 6646
rect 14308 6582 14310 6634
rect 14362 6582 14364 6634
rect 14308 6132 14364 6582
rect 14252 6076 14364 6132
rect 14476 6578 14532 8094
rect 14476 6526 14478 6578
rect 14530 6526 14532 6578
rect 14476 6132 14532 6526
rect 14140 6020 14196 6030
rect 14252 6020 14308 6076
rect 14476 6066 14532 6076
rect 14588 7476 14644 7486
rect 14196 5964 14308 6020
rect 14140 5933 14196 5964
rect 14140 5881 14142 5933
rect 14194 5881 14196 5933
rect 14140 5869 14196 5881
rect 14252 5236 14308 5246
rect 14252 5142 14308 5180
rect 13804 4498 13860 4508
rect 13916 4004 13972 4014
rect 13580 3724 13748 3780
rect 13468 3502 13470 3554
rect 13522 3502 13524 3554
rect 13468 3490 13524 3502
rect 13580 3556 13636 3566
rect 13580 3462 13636 3500
rect 11788 3332 11844 3342
rect 11788 3330 11956 3332
rect 11788 3278 11790 3330
rect 11842 3278 11956 3330
rect 11788 3276 11956 3278
rect 11788 3266 11844 3276
rect 10892 802 10948 812
rect 11900 800 11956 3276
rect 13692 800 13748 3724
rect 13916 3526 13972 3948
rect 13916 3474 13918 3526
rect 13970 3474 13972 3526
rect 14588 3556 14644 7420
rect 15148 7476 15204 7486
rect 15148 7382 15204 7420
rect 15540 7476 15596 7486
rect 15540 7362 15596 7420
rect 15540 7310 15542 7362
rect 15594 7310 15596 7362
rect 15198 7084 15462 7094
rect 15254 7028 15302 7084
rect 15358 7028 15406 7084
rect 15198 7018 15462 7028
rect 15354 6916 15410 6926
rect 15540 6916 15596 7310
rect 15354 6822 15410 6860
rect 15484 6860 15596 6916
rect 15484 6468 15540 6860
rect 15596 6692 15652 6702
rect 15596 6598 15652 6636
rect 15484 6412 15652 6468
rect 15148 5684 15204 5722
rect 15148 5618 15204 5628
rect 15198 5516 15462 5526
rect 15254 5460 15302 5516
rect 15358 5460 15406 5516
rect 15198 5450 15462 5460
rect 15372 5122 15428 5134
rect 15372 5070 15374 5122
rect 15426 5070 15428 5122
rect 15372 4452 15428 5070
rect 15484 5124 15540 5134
rect 15596 5124 15652 6412
rect 15540 5068 15652 5124
rect 15820 6132 15876 8766
rect 16604 7812 16660 11900
rect 17052 11508 17108 11900
rect 17052 11442 17108 11452
rect 17276 12852 17332 12862
rect 17276 11396 17332 12796
rect 18060 12292 18116 12302
rect 18172 12292 18228 13356
rect 19180 13300 19236 18060
rect 19292 17556 19348 17566
rect 19292 16882 19348 17500
rect 19404 16996 19460 18620
rect 19740 18564 19796 19068
rect 19964 19124 20020 19180
rect 19964 19058 20020 19068
rect 20188 19178 20244 19180
rect 20188 19126 20190 19178
rect 20242 19126 20244 19178
rect 19860 18844 20124 18854
rect 19916 18788 19964 18844
rect 20020 18788 20068 18844
rect 19860 18778 20124 18788
rect 19964 18564 20020 18574
rect 19740 18562 20020 18564
rect 19740 18510 19966 18562
rect 20018 18510 20020 18562
rect 19740 18508 20020 18510
rect 19964 18498 20020 18508
rect 20188 18340 20244 19126
rect 20020 17556 20076 17566
rect 20020 17462 20076 17500
rect 19860 17276 20124 17286
rect 19916 17220 19964 17276
rect 20020 17220 20068 17276
rect 19860 17210 20124 17220
rect 20188 17108 20244 18284
rect 20300 18452 20356 18462
rect 20300 18338 20356 18396
rect 20300 18286 20302 18338
rect 20354 18286 20356 18338
rect 20300 18274 20356 18286
rect 20412 18450 20468 18462
rect 20412 18398 20414 18450
rect 20466 18398 20468 18450
rect 20412 18116 20468 18398
rect 20524 18228 20580 19180
rect 20636 19066 20692 19078
rect 20636 19014 20638 19066
rect 20690 19014 20692 19066
rect 20636 18900 20692 19014
rect 20636 18834 20692 18844
rect 20748 18450 20804 18462
rect 21196 18452 21252 18462
rect 20748 18398 20750 18450
rect 20802 18398 20804 18450
rect 20748 18340 20804 18398
rect 20748 18274 20804 18284
rect 21084 18450 21252 18452
rect 21084 18398 21198 18450
rect 21250 18398 21252 18450
rect 21084 18396 21252 18398
rect 20524 18162 20580 18172
rect 21084 18228 21140 18396
rect 21196 18386 21252 18396
rect 21532 18452 21588 19182
rect 20412 17780 20468 18060
rect 20412 17724 20580 17780
rect 20412 17444 20468 17454
rect 20076 17052 20244 17108
rect 20300 17332 20356 17342
rect 20076 17050 20132 17052
rect 20076 16998 20078 17050
rect 20130 16998 20132 17050
rect 20076 16986 20132 16998
rect 19404 16930 19460 16940
rect 19292 16830 19294 16882
rect 19346 16830 19348 16882
rect 19292 15316 19348 16830
rect 19628 16884 19684 16894
rect 19628 16266 19684 16828
rect 19628 16214 19630 16266
rect 19682 16214 19684 16266
rect 19628 16202 19684 16214
rect 19964 16882 20020 16894
rect 19964 16830 19966 16882
rect 20018 16830 20020 16882
rect 19516 16100 19572 16110
rect 19964 16100 20020 16830
rect 20300 16772 20356 17276
rect 20412 16938 20468 17388
rect 20524 17108 20580 17724
rect 20748 17668 20804 17678
rect 20524 17042 20580 17052
rect 20636 17666 20804 17668
rect 20636 17614 20750 17666
rect 20802 17614 20804 17666
rect 20636 17612 20804 17614
rect 20412 16886 20414 16938
rect 20466 16886 20468 16938
rect 20412 16874 20468 16886
rect 20524 16910 20580 16922
rect 20524 16884 20526 16910
rect 20578 16884 20580 16910
rect 20524 16818 20580 16828
rect 20300 16716 20468 16772
rect 19516 16098 19796 16100
rect 19516 16046 19518 16098
rect 19570 16046 19796 16098
rect 19516 16044 19796 16046
rect 19516 16034 19572 16044
rect 19292 15250 19348 15260
rect 19628 15876 19684 15886
rect 19628 14642 19684 15820
rect 19740 15428 19796 16044
rect 20412 16098 20468 16716
rect 20636 16548 20692 17612
rect 20748 17602 20804 17612
rect 20972 17108 21028 17118
rect 20748 16940 20916 16996
rect 20748 16938 20804 16940
rect 20748 16886 20750 16938
rect 20802 16886 20804 16938
rect 20748 16874 20804 16886
rect 19964 16034 20020 16044
rect 20244 16042 20300 16054
rect 20244 15990 20246 16042
rect 20298 15990 20300 16042
rect 20412 16046 20414 16098
rect 20466 16046 20468 16098
rect 20412 16034 20468 16046
rect 20524 16492 20692 16548
rect 20748 16772 20804 16782
rect 20244 15988 20300 15990
rect 20244 15932 20356 15988
rect 19860 15708 20124 15718
rect 19916 15652 19964 15708
rect 20020 15652 20068 15708
rect 19860 15642 20124 15652
rect 20300 15540 20356 15932
rect 20524 15876 20580 16492
rect 20636 16212 20692 16222
rect 20748 16212 20804 16716
rect 20860 16548 20916 16940
rect 20972 16938 21028 17052
rect 20972 16886 20974 16938
rect 21026 16886 21028 16938
rect 20972 16874 21028 16886
rect 21084 16772 21140 18172
rect 21532 17444 21588 18396
rect 21532 17378 21588 17388
rect 21644 17220 21700 19964
rect 21756 19796 21812 20748
rect 21756 19730 21812 19740
rect 21812 19460 21868 19470
rect 21812 19366 21868 19404
rect 21980 19236 22036 19246
rect 21868 19234 22036 19236
rect 21868 19182 21982 19234
rect 22034 19182 22036 19234
rect 21868 19180 22036 19182
rect 21868 18676 21924 19180
rect 21980 19170 22036 19180
rect 21868 18620 22036 18676
rect 21868 18116 21924 18620
rect 21980 18506 22036 18620
rect 21980 18454 21982 18506
rect 22034 18454 22036 18506
rect 21980 18442 22036 18454
rect 22092 18564 22148 18574
rect 22092 18478 22148 18508
rect 22092 18426 22094 18478
rect 22146 18426 22148 18478
rect 22092 18414 22148 18426
rect 21868 18050 21924 18060
rect 21532 17164 21700 17220
rect 21756 17556 21812 17566
rect 21252 16884 21308 16894
rect 21252 16790 21308 16828
rect 20860 16482 20916 16492
rect 20972 16716 21140 16772
rect 20636 16210 20804 16212
rect 20636 16158 20638 16210
rect 20690 16158 20804 16210
rect 20636 16156 20804 16158
rect 20636 16146 20692 16156
rect 20524 15810 20580 15820
rect 20804 16042 20860 16054
rect 20804 15990 20806 16042
rect 20858 15990 20860 16042
rect 20804 15540 20860 15990
rect 20300 15484 20468 15540
rect 19964 15428 20020 15438
rect 19740 15426 20020 15428
rect 19740 15374 19966 15426
rect 20018 15374 20020 15426
rect 19740 15372 20020 15374
rect 19964 15092 20020 15372
rect 20412 15092 20468 15484
rect 20804 15474 20860 15484
rect 20748 15316 20804 15326
rect 20748 15202 20804 15260
rect 20748 15150 20750 15202
rect 20802 15150 20804 15202
rect 20748 15138 20804 15150
rect 19964 15036 20356 15092
rect 19628 14590 19630 14642
rect 19682 14590 19684 14642
rect 19628 14578 19684 14590
rect 18956 13244 19236 13300
rect 19404 14532 19460 14542
rect 20076 14532 20132 14542
rect 19404 13972 19460 14476
rect 18340 12852 18396 12862
rect 18340 12758 18396 12796
rect 18060 12290 18228 12292
rect 18060 12238 18062 12290
rect 18114 12238 18228 12290
rect 18060 12236 18228 12238
rect 18060 12180 18116 12236
rect 17668 11508 17724 11518
rect 17668 11414 17724 11452
rect 17948 11396 18004 11406
rect 18060 11396 18116 12124
rect 17276 11394 17612 11396
rect 17276 11342 17278 11394
rect 17330 11342 17612 11394
rect 17276 11340 17612 11342
rect 17276 11330 17332 11340
rect 17556 10836 17612 11340
rect 17948 11394 18116 11396
rect 17948 11342 17950 11394
rect 18002 11342 18116 11394
rect 17948 11340 18116 11342
rect 18732 11396 18788 11406
rect 17948 11330 18004 11340
rect 18732 11302 18788 11340
rect 18956 10846 19012 13244
rect 19404 13188 19460 13916
rect 19740 14476 20076 14532
rect 19628 13860 19684 13870
rect 19740 13860 19796 14476
rect 20076 14438 20132 14476
rect 20300 14530 20356 15036
rect 20412 15026 20468 15036
rect 20580 14756 20636 14766
rect 20972 14756 21028 16716
rect 21532 16548 21588 17164
rect 21756 17108 21812 17500
rect 21756 16926 21812 17052
rect 22204 16996 22260 20972
rect 22316 21364 22372 21374
rect 22316 19012 22372 21308
rect 22428 19460 22484 19470
rect 22428 19234 22484 19404
rect 22428 19182 22430 19234
rect 22482 19182 22484 19234
rect 22428 19170 22484 19182
rect 22316 18956 22484 19012
rect 22316 18478 22372 18490
rect 22316 18426 22318 18478
rect 22370 18426 22372 18478
rect 22316 18228 22372 18426
rect 22316 18162 22372 18172
rect 22428 18004 22484 18956
rect 22540 18478 22596 18490
rect 22540 18452 22542 18478
rect 22594 18452 22596 18478
rect 22540 18386 22596 18396
rect 21756 16874 21758 16926
rect 21810 16874 21812 16926
rect 22117 16940 22260 16996
rect 22316 17948 22484 18004
rect 22316 17332 22372 17948
rect 22652 17724 22708 21532
rect 22764 21364 22820 23102
rect 23436 23156 23492 23166
rect 23212 22370 23268 22382
rect 23212 22318 23214 22370
rect 23266 22318 23268 22370
rect 23212 21588 23268 22318
rect 23436 22370 23492 23100
rect 23548 22484 23604 25340
rect 23660 24164 23716 27580
rect 24050 27412 24106 27422
rect 23772 27074 23828 27086
rect 23772 27022 23774 27074
rect 23826 27022 23828 27074
rect 23772 26180 23828 27022
rect 23884 27076 23940 27086
rect 23884 26982 23940 27020
rect 24050 27074 24106 27356
rect 24050 27022 24052 27074
rect 24104 27022 24106 27074
rect 24050 27010 24106 27022
rect 24220 26964 24276 26974
rect 24220 26290 24276 26908
rect 24220 26238 24222 26290
rect 24274 26238 24276 26290
rect 24220 26226 24276 26238
rect 23772 26114 23828 26124
rect 23660 23716 23716 24108
rect 23660 23650 23716 23660
rect 23772 25620 23828 25630
rect 23772 22820 23828 25564
rect 24220 25508 24276 25518
rect 24220 25414 24276 25452
rect 24108 25338 24164 25350
rect 23884 25284 23940 25294
rect 23884 24836 23940 25228
rect 24108 25286 24110 25338
rect 24162 25286 24164 25338
rect 23996 24836 24052 24846
rect 23884 24834 24052 24836
rect 23884 24782 23998 24834
rect 24050 24782 24052 24834
rect 23884 24780 24052 24782
rect 23996 24770 24052 24780
rect 23884 24164 23940 24174
rect 23884 24050 23940 24108
rect 23884 23998 23886 24050
rect 23938 23998 23940 24050
rect 23884 23986 23940 23998
rect 24108 24052 24164 25286
rect 24332 25060 24388 30156
rect 24556 30210 24612 30222
rect 24556 30158 24558 30210
rect 24610 30158 24612 30210
rect 24556 29652 24612 30158
rect 24556 29586 24612 29596
rect 24780 29540 24836 30380
rect 25004 29876 25060 29886
rect 25676 29876 25732 30942
rect 25788 30826 25844 31724
rect 25788 30774 25790 30826
rect 25842 30774 25844 30826
rect 25788 30762 25844 30774
rect 24780 29484 24948 29540
rect 24724 29316 24780 29326
rect 24724 29222 24780 29260
rect 24522 29036 24786 29046
rect 24578 28980 24626 29036
rect 24682 28980 24730 29036
rect 24522 28970 24786 28980
rect 24668 28868 24724 28878
rect 24500 28756 24556 28766
rect 24500 28662 24556 28700
rect 24668 28308 24724 28812
rect 24780 28756 24836 28766
rect 24780 28642 24836 28700
rect 24780 28590 24782 28642
rect 24834 28590 24836 28642
rect 24780 28578 24836 28590
rect 24892 28642 24948 29484
rect 24892 28590 24894 28642
rect 24946 28590 24948 28642
rect 24892 28420 24948 28590
rect 25004 28654 25060 29820
rect 25340 29820 25732 29876
rect 25340 28868 25396 29820
rect 25508 29540 25564 29550
rect 25508 29446 25564 29484
rect 25676 29540 25732 29550
rect 25452 28868 25508 28878
rect 25340 28866 25508 28868
rect 25340 28814 25454 28866
rect 25506 28814 25508 28866
rect 25340 28812 25508 28814
rect 25452 28802 25508 28812
rect 25004 28642 25114 28654
rect 25004 28590 25060 28642
rect 25112 28590 25114 28642
rect 25004 28588 25114 28590
rect 25058 28578 25114 28588
rect 25116 28420 25172 28430
rect 24892 28364 25060 28420
rect 24668 28252 24948 28308
rect 24668 28026 24724 28038
rect 24668 27974 24670 28026
rect 24722 27974 24724 28026
rect 24668 27972 24724 27974
rect 24668 27906 24724 27916
rect 24556 27860 24612 27870
rect 24556 27766 24612 27804
rect 24522 27468 24786 27478
rect 24578 27412 24626 27468
rect 24682 27412 24730 27468
rect 24522 27402 24786 27412
rect 24444 27300 24500 27310
rect 24892 27300 24948 28252
rect 24444 27298 24948 27300
rect 24444 27246 24446 27298
rect 24498 27246 24948 27298
rect 24444 27244 24948 27246
rect 25004 27860 25060 28364
rect 25004 27300 25060 27804
rect 24444 27234 24500 27244
rect 25004 27234 25060 27244
rect 25676 28420 25732 29484
rect 25788 29204 25844 29214
rect 25788 28642 25844 29148
rect 25900 28868 25956 32510
rect 26124 32450 26180 32462
rect 26124 32398 26126 32450
rect 26178 32398 26180 32450
rect 26012 31750 26068 31762
rect 26012 31698 26014 31750
rect 26066 31698 26068 31750
rect 26012 30994 26068 31698
rect 26124 31220 26180 32398
rect 26460 31556 26516 33266
rect 26842 32676 26898 32686
rect 26842 32612 26898 32620
rect 26572 32562 26628 32574
rect 26572 32510 26574 32562
rect 26626 32510 26628 32562
rect 26572 32340 26628 32510
rect 26684 32564 26740 32574
rect 26842 32560 26844 32612
rect 26896 32560 26898 32612
rect 26842 32548 26898 32560
rect 26684 32470 26740 32508
rect 27244 32450 27300 33740
rect 27692 33460 27748 34750
rect 27692 32788 27748 33404
rect 27804 33348 27860 33358
rect 27804 33254 27860 33292
rect 28028 33236 28084 34862
rect 28140 33460 28196 35420
rect 28252 34916 28308 34926
rect 28532 34916 28588 34926
rect 28252 34914 28420 34916
rect 28252 34862 28254 34914
rect 28306 34862 28420 34914
rect 28252 34860 28420 34862
rect 28252 34850 28308 34860
rect 28252 34130 28308 34142
rect 28252 34078 28254 34130
rect 28306 34078 28308 34130
rect 28252 33684 28308 34078
rect 28252 33618 28308 33628
rect 28364 33460 28420 34860
rect 28532 34822 28588 34860
rect 28924 34468 28980 39200
rect 29184 36092 29448 36102
rect 29240 36036 29288 36092
rect 29344 36036 29392 36092
rect 29184 36026 29448 36036
rect 29036 35474 29092 35486
rect 29036 35422 29038 35474
rect 29090 35422 29092 35474
rect 29036 35140 29092 35422
rect 29036 35074 29092 35084
rect 29708 35252 29764 35262
rect 29036 34916 29092 34926
rect 29036 34822 29092 34860
rect 28140 33404 28308 33460
rect 27692 32722 27748 32732
rect 27916 33180 28028 33236
rect 27244 32398 27246 32450
rect 27298 32398 27300 32450
rect 27244 32386 27300 32398
rect 26572 32274 26628 32284
rect 26460 31500 26740 31556
rect 26124 31154 26180 31164
rect 26012 30942 26014 30994
rect 26066 30942 26068 30994
rect 26012 30212 26068 30942
rect 26012 29204 26068 30156
rect 26460 30996 26516 31006
rect 26460 30324 26516 30940
rect 26460 30210 26516 30268
rect 26460 30158 26462 30210
rect 26514 30158 26516 30210
rect 26460 30146 26516 30158
rect 26124 30100 26180 30110
rect 26124 29540 26180 30044
rect 26124 29453 26180 29484
rect 26124 29401 26126 29453
rect 26178 29401 26180 29453
rect 26124 29389 26180 29401
rect 26012 29138 26068 29148
rect 25900 28802 25956 28812
rect 25788 28590 25790 28642
rect 25842 28590 25844 28642
rect 25788 28578 25844 28590
rect 26572 28642 26628 28654
rect 26572 28590 26574 28642
rect 26626 28590 26628 28642
rect 25676 28364 25844 28420
rect 25116 27412 25172 28364
rect 25583 27972 25639 27982
rect 25583 27914 25639 27916
rect 25340 27860 25396 27870
rect 25583 27862 25585 27914
rect 25637 27862 25639 27914
rect 25583 27850 25639 27862
rect 25340 27766 25396 27804
rect 25116 27074 25172 27356
rect 25676 27748 25732 27758
rect 25116 27022 25118 27074
rect 25170 27022 25172 27074
rect 25564 27188 25620 27198
rect 25116 27010 25172 27022
rect 25340 27018 25396 27030
rect 25004 26964 25060 26974
rect 25340 26966 25342 27018
rect 25394 26966 25396 27018
rect 24892 26852 24948 26862
rect 25004 26852 25172 26908
rect 24556 26180 24612 26190
rect 24556 26086 24612 26124
rect 24522 25900 24786 25910
rect 24578 25844 24626 25900
rect 24682 25844 24730 25900
rect 24522 25834 24786 25844
rect 24780 25732 24836 25742
rect 24780 25506 24836 25676
rect 24780 25454 24782 25506
rect 24834 25454 24836 25506
rect 24780 25396 24836 25454
rect 24780 25330 24836 25340
rect 24332 25004 24668 25060
rect 24332 24724 24388 25004
rect 24612 24946 24668 25004
rect 24612 24894 24614 24946
rect 24666 24894 24668 24946
rect 24612 24882 24668 24894
rect 24332 24164 24388 24668
rect 24522 24332 24786 24342
rect 24578 24276 24626 24332
rect 24682 24276 24730 24332
rect 24522 24266 24786 24276
rect 24332 24108 24556 24164
rect 24108 23986 24164 23996
rect 24500 24050 24556 24108
rect 24500 23998 24502 24050
rect 24554 23998 24556 24050
rect 24500 23986 24556 23998
rect 23772 22764 24276 22820
rect 23548 22418 23604 22428
rect 23436 22318 23438 22370
rect 23490 22318 23492 22370
rect 23436 22260 23492 22318
rect 23716 22372 23772 22382
rect 23716 22278 23772 22316
rect 23436 22194 23492 22204
rect 23212 21522 23268 21532
rect 22764 21298 22820 21308
rect 24052 21474 24108 21486
rect 24052 21422 24054 21474
rect 24106 21422 24108 21474
rect 24052 21140 24108 21422
rect 23772 21084 24108 21140
rect 23772 20774 23828 21084
rect 24220 21028 24276 22764
rect 24522 22764 24786 22774
rect 24578 22708 24626 22764
rect 24682 22708 24730 22764
rect 24522 22698 24786 22708
rect 24522 21196 24786 21206
rect 24578 21140 24626 21196
rect 24682 21140 24730 21196
rect 24522 21130 24786 21140
rect 24892 21038 24948 26796
rect 25004 26516 25060 26526
rect 25004 25508 25060 26460
rect 25116 25742 25172 26852
rect 25228 26906 25284 26918
rect 25228 26854 25230 26906
rect 25282 26854 25284 26906
rect 25228 26290 25284 26854
rect 25340 26516 25396 26966
rect 25564 26964 25620 27132
rect 25676 27074 25732 27692
rect 25676 27022 25678 27074
rect 25730 27022 25732 27074
rect 25676 27010 25732 27022
rect 25564 26898 25620 26908
rect 25340 26450 25396 26460
rect 25676 26628 25732 26638
rect 25228 26238 25230 26290
rect 25282 26238 25284 26290
rect 25564 26290 25620 26302
rect 25228 26226 25284 26238
rect 25396 26234 25452 26246
rect 25396 26182 25398 26234
rect 25450 26182 25452 26234
rect 25396 25844 25452 26182
rect 25340 25788 25452 25844
rect 25564 26238 25566 26290
rect 25618 26238 25620 26290
rect 25116 25730 25228 25742
rect 25116 25678 25174 25730
rect 25226 25678 25228 25730
rect 25116 25676 25228 25678
rect 25172 25666 25228 25676
rect 25340 25732 25396 25788
rect 25564 25732 25620 26238
rect 25676 26290 25732 26572
rect 25676 26238 25678 26290
rect 25730 26238 25732 26290
rect 25676 26226 25732 26238
rect 25788 26068 25844 28364
rect 26572 28084 26628 28590
rect 26572 28018 26628 28028
rect 26460 27860 26516 27898
rect 26460 27794 26516 27804
rect 26348 27412 26404 27422
rect 26012 27300 26068 27310
rect 26012 27074 26068 27244
rect 26012 27022 26014 27074
rect 26066 27022 26068 27074
rect 26012 27010 26068 27022
rect 26236 27188 26292 27198
rect 26236 27074 26292 27132
rect 26236 27022 26238 27074
rect 26290 27022 26292 27074
rect 26236 27010 26292 27022
rect 25900 26964 25956 26974
rect 26348 26908 26404 27356
rect 26516 27076 26572 27114
rect 26516 27010 26572 27020
rect 25900 26852 26012 26908
rect 26348 26852 26628 26908
rect 25956 26402 26012 26852
rect 26572 26514 26628 26852
rect 26572 26462 26574 26514
rect 26626 26462 26628 26514
rect 26572 26450 26628 26462
rect 25956 26350 25958 26402
rect 26010 26350 26012 26402
rect 25956 26338 26012 26350
rect 25788 26002 25844 26012
rect 26236 26290 26292 26302
rect 26236 26238 26238 26290
rect 26290 26238 26292 26290
rect 25340 25666 25396 25676
rect 25452 25676 25620 25732
rect 25452 25508 25508 25676
rect 25004 25442 25060 25452
rect 25340 25506 25508 25508
rect 25340 25454 25454 25506
rect 25506 25454 25508 25506
rect 25340 25452 25508 25454
rect 25340 24498 25396 25452
rect 25452 25442 25508 25452
rect 25676 25508 25732 25518
rect 26068 25508 26124 25518
rect 25676 25506 25844 25508
rect 25676 25454 25678 25506
rect 25730 25454 25844 25506
rect 25676 25452 25844 25454
rect 25676 25442 25732 25452
rect 25340 24446 25342 24498
rect 25394 24446 25396 24498
rect 25340 24162 25396 24446
rect 25340 24110 25342 24162
rect 25394 24110 25396 24162
rect 25340 24098 25396 24110
rect 25788 25172 25844 25452
rect 26068 25414 26124 25452
rect 25676 23938 25732 23950
rect 25676 23886 25678 23938
rect 25730 23886 25732 23938
rect 25564 23154 25620 23166
rect 25564 23102 25566 23154
rect 25618 23102 25620 23154
rect 25340 23042 25396 23054
rect 25340 22990 25342 23042
rect 25394 22990 25396 23042
rect 25340 21812 25396 22990
rect 25564 22484 25620 23102
rect 25564 22418 25620 22428
rect 25676 22932 25732 23886
rect 25676 22372 25732 22876
rect 25676 22278 25732 22316
rect 25340 21746 25396 21756
rect 25788 21700 25844 25116
rect 26236 24498 26292 26238
rect 26516 25282 26572 25294
rect 26516 25230 26518 25282
rect 26570 25230 26572 25282
rect 26516 25172 26572 25230
rect 26516 24724 26572 25116
rect 26516 24658 26572 24668
rect 26236 24446 26238 24498
rect 26290 24446 26292 24498
rect 26236 24434 26292 24446
rect 26572 24498 26628 24510
rect 26572 24446 26574 24498
rect 26626 24446 26628 24498
rect 26572 23938 26628 24446
rect 26572 23886 26574 23938
rect 26626 23886 26628 23938
rect 26572 23874 26628 23886
rect 26684 23716 26740 31500
rect 26796 31220 26852 31230
rect 26796 30994 26852 31164
rect 26796 30942 26798 30994
rect 26850 30942 26852 30994
rect 26796 30930 26852 30942
rect 27020 31108 27076 31118
rect 27020 30670 27076 31052
rect 27916 30996 27972 33180
rect 28028 33170 28084 33180
rect 28028 32589 28084 32601
rect 28028 32537 28030 32589
rect 28082 32537 28084 32589
rect 28028 32452 28084 32537
rect 28028 32386 28084 32396
rect 27020 30660 27132 30670
rect 27916 30660 27972 30940
rect 28140 32116 28196 32126
rect 27020 30604 27076 30660
rect 27076 30210 27132 30604
rect 27076 30158 27078 30210
rect 27130 30158 27132 30210
rect 27076 30146 27132 30158
rect 27692 30604 27972 30660
rect 28028 30884 28084 30894
rect 27692 30210 27748 30604
rect 27692 30158 27694 30210
rect 27746 30158 27748 30210
rect 27692 30146 27748 30158
rect 28028 30210 28084 30828
rect 28028 30158 28030 30210
rect 28082 30158 28084 30210
rect 28028 29652 28084 30158
rect 28028 29586 28084 29596
rect 28140 30210 28196 32060
rect 28140 30158 28142 30210
rect 28194 30158 28196 30210
rect 27916 29316 27972 29326
rect 26796 29204 26852 29214
rect 26796 29110 26852 29148
rect 26964 28420 27020 28430
rect 26964 27914 27020 28364
rect 26796 27858 26852 27870
rect 26796 27806 26798 27858
rect 26850 27806 26852 27858
rect 26964 27862 26966 27914
rect 27018 27862 27020 27914
rect 27132 27972 27188 27982
rect 27132 27878 27188 27916
rect 26964 27850 27020 27862
rect 27244 27858 27300 27870
rect 26796 27300 26852 27806
rect 27244 27806 27246 27858
rect 27298 27806 27300 27858
rect 26964 27300 27020 27310
rect 27244 27300 27300 27806
rect 27524 27860 27580 27870
rect 27804 27860 27860 27870
rect 27524 27858 27860 27860
rect 27524 27806 27526 27858
rect 27578 27806 27806 27858
rect 27858 27806 27860 27858
rect 27524 27804 27860 27806
rect 27524 27794 27580 27804
rect 27804 27794 27860 27804
rect 26796 27298 27020 27300
rect 26796 27246 26966 27298
rect 27018 27246 27020 27298
rect 26796 27244 27020 27246
rect 26964 27234 27020 27244
rect 27132 27244 27300 27300
rect 27356 27636 27412 27646
rect 27916 27636 27972 29260
rect 28140 29316 28196 30158
rect 28140 29250 28196 29260
rect 28140 28084 28196 28094
rect 28140 27990 28196 28028
rect 28252 27860 28308 33404
rect 28364 33394 28420 33404
rect 28588 34412 28980 34468
rect 29184 34524 29448 34534
rect 29240 34468 29288 34524
rect 29344 34468 29392 34524
rect 29184 34458 29448 34468
rect 28476 29986 28532 29998
rect 28476 29934 28478 29986
rect 28530 29934 28532 29986
rect 28364 29652 28420 29662
rect 28364 28532 28420 29596
rect 28476 29316 28532 29934
rect 28476 29250 28532 29260
rect 28476 29092 28532 29102
rect 28476 28754 28532 29036
rect 28476 28702 28478 28754
rect 28530 28702 28532 28754
rect 28476 28690 28532 28702
rect 28364 28476 28532 28532
rect 27132 26908 27188 27244
rect 27020 26852 27188 26908
rect 27244 27074 27300 27086
rect 27244 27022 27246 27074
rect 27298 27022 27300 27074
rect 27244 26964 27300 27022
rect 27356 27076 27412 27580
rect 27356 26982 27412 27020
rect 27468 27580 27972 27636
rect 28140 27804 28308 27860
rect 27244 26898 27300 26908
rect 27020 26180 27076 26852
rect 27188 26516 27244 26526
rect 27188 26422 27244 26460
rect 27020 26114 27076 26124
rect 27132 24498 27188 24510
rect 27132 24446 27134 24498
rect 27186 24446 27188 24498
rect 26908 24052 26964 24062
rect 27132 24052 27188 24446
rect 26908 24050 27188 24052
rect 26908 23998 26910 24050
rect 26962 23998 27188 24050
rect 26908 23996 27188 23998
rect 26908 23986 26964 23996
rect 27244 23938 27300 23950
rect 25788 21634 25844 21644
rect 25900 23660 26740 23716
rect 27020 23882 27076 23894
rect 27020 23830 27022 23882
rect 27074 23830 27076 23882
rect 25508 21615 25564 21627
rect 25228 21586 25284 21598
rect 25508 21588 25510 21615
rect 25228 21534 25230 21586
rect 25282 21534 25284 21586
rect 25228 21364 25284 21534
rect 25228 21298 25284 21308
rect 25340 21563 25510 21588
rect 25562 21563 25564 21615
rect 25340 21532 25564 21563
rect 23772 20722 23774 20774
rect 23826 20722 23828 20774
rect 23436 20132 23492 20142
rect 22876 20020 22932 20030
rect 22876 19926 22932 19964
rect 23436 20018 23492 20076
rect 23436 19966 23438 20018
rect 23490 19966 23492 20018
rect 23436 19954 23492 19966
rect 23772 20020 23828 20722
rect 24108 20972 24276 21028
rect 24836 21026 24948 21038
rect 24836 20974 24838 21026
rect 24890 20974 24948 21026
rect 24836 20972 24948 20974
rect 24108 20802 24164 20972
rect 24836 20962 24892 20972
rect 24108 20750 24110 20802
rect 24162 20750 24164 20802
rect 24556 20802 24612 20814
rect 24108 20580 24164 20750
rect 24108 20514 24164 20524
rect 24276 20746 24332 20758
rect 24276 20694 24278 20746
rect 24330 20694 24332 20746
rect 24556 20750 24558 20802
rect 24610 20750 24612 20802
rect 23996 20132 24052 20142
rect 24276 20132 24332 20694
rect 24444 20690 24500 20702
rect 24444 20638 24446 20690
rect 24498 20638 24500 20690
rect 24276 20076 24388 20132
rect 23772 19964 23940 20020
rect 23436 19796 23492 19806
rect 22988 19572 23044 19582
rect 22764 19234 22820 19246
rect 22764 19182 22766 19234
rect 22818 19182 22820 19234
rect 22764 18564 22820 19182
rect 22764 18498 22820 18508
rect 22988 19236 23044 19516
rect 22988 19143 22990 19180
rect 23042 19143 23044 19180
rect 22820 18340 22876 18350
rect 22988 18340 23044 19143
rect 23100 19346 23156 19358
rect 23100 19294 23102 19346
rect 23154 19294 23156 19346
rect 23100 19012 23156 19294
rect 23436 19234 23492 19740
rect 23772 19796 23828 19806
rect 23772 19702 23828 19740
rect 23772 19572 23828 19582
rect 23772 19236 23828 19516
rect 23436 19182 23438 19234
rect 23490 19182 23492 19234
rect 23436 19170 23492 19182
rect 23548 19234 23828 19236
rect 23548 19182 23774 19234
rect 23826 19182 23828 19234
rect 23548 19180 23828 19182
rect 23100 18946 23156 18956
rect 23380 18564 23436 18574
rect 23380 18470 23436 18508
rect 22820 18338 23044 18340
rect 22820 18286 22822 18338
rect 22874 18286 23044 18338
rect 22820 18284 23044 18286
rect 22820 18274 22876 18284
rect 22876 18116 22932 18126
rect 22652 17668 22820 17724
rect 21980 16884 22036 16894
rect 21756 16862 21812 16874
rect 21868 16882 22036 16884
rect 21868 16830 21982 16882
rect 22034 16830 22036 16882
rect 21868 16828 22036 16830
rect 21644 16770 21700 16782
rect 21644 16718 21646 16770
rect 21698 16718 21700 16770
rect 21644 16660 21700 16718
rect 21868 16772 21924 16828
rect 21980 16818 22036 16828
rect 22117 16772 22173 16940
rect 22316 16882 22372 17276
rect 22652 17556 22708 17566
rect 22316 16830 22318 16882
rect 22370 16830 22372 16882
rect 22316 16818 22372 16830
rect 22484 17050 22540 17062
rect 22484 16998 22486 17050
rect 22538 16998 22540 17050
rect 21644 16604 21812 16660
rect 21756 16548 21812 16604
rect 21532 16492 21700 16548
rect 21308 16100 21364 16110
rect 21308 16006 21364 16044
rect 21476 16042 21532 16054
rect 21476 15990 21478 16042
rect 21530 15990 21532 16042
rect 21476 15876 21532 15990
rect 21476 15810 21532 15820
rect 21122 15540 21178 15550
rect 21122 15352 21178 15484
rect 21122 15300 21124 15352
rect 21176 15300 21178 15352
rect 21122 15148 21178 15300
rect 21308 15314 21364 15326
rect 21308 15262 21310 15314
rect 21362 15262 21364 15314
rect 21122 15092 21198 15148
rect 21142 14980 21198 15092
rect 21308 15092 21364 15262
rect 21308 15026 21364 15036
rect 21420 15314 21476 15326
rect 21420 15262 21422 15314
rect 21474 15262 21476 15314
rect 21142 14914 21198 14924
rect 21420 14756 21476 15262
rect 21644 15316 21700 16492
rect 21756 16482 21812 16492
rect 21868 16212 21924 16716
rect 22092 16716 22173 16772
rect 21868 16146 21924 16156
rect 21980 16660 22036 16670
rect 21756 16100 21812 16110
rect 21756 15426 21812 16044
rect 21980 16098 22036 16604
rect 21980 16046 21982 16098
rect 22034 16046 22036 16098
rect 21980 15876 22036 16046
rect 21980 15810 22036 15820
rect 21756 15374 21758 15426
rect 21810 15374 21812 15426
rect 21756 15362 21812 15374
rect 21644 15250 21700 15260
rect 21924 15258 21980 15270
rect 21924 15206 21926 15258
rect 21978 15206 21980 15258
rect 20580 14754 21028 14756
rect 20580 14702 20582 14754
rect 20634 14702 21028 14754
rect 20580 14700 21028 14702
rect 21308 14700 21476 14756
rect 21644 15092 21700 15102
rect 20580 14690 20636 14700
rect 20300 14478 20302 14530
rect 20354 14478 20356 14530
rect 20300 14466 20356 14478
rect 21308 14532 21364 14700
rect 21308 14438 21364 14476
rect 21476 14474 21532 14486
rect 21476 14422 21478 14474
rect 21530 14422 21532 14474
rect 19860 14140 20124 14150
rect 19916 14084 19964 14140
rect 20020 14084 20068 14140
rect 19860 14074 20124 14084
rect 20860 14084 20916 14094
rect 19628 13858 19796 13860
rect 19628 13806 19630 13858
rect 19682 13806 19796 13858
rect 19628 13804 19796 13806
rect 19628 13794 19684 13804
rect 19180 13186 19460 13188
rect 19180 13134 19406 13186
rect 19458 13134 19460 13186
rect 19180 13132 19460 13134
rect 19180 12178 19236 13132
rect 19404 13122 19460 13132
rect 20188 13746 20244 13758
rect 20188 13694 20190 13746
rect 20242 13694 20244 13746
rect 20188 12964 20244 13694
rect 19860 12572 20124 12582
rect 19916 12516 19964 12572
rect 20020 12516 20068 12572
rect 19860 12506 20124 12516
rect 19180 12126 19182 12178
rect 19234 12126 19236 12178
rect 19180 12114 19236 12126
rect 19628 12180 19684 12190
rect 19628 12086 19684 12124
rect 20188 12180 20244 12908
rect 20524 12964 20580 12974
rect 20188 12114 20244 12124
rect 20412 12852 20468 12862
rect 20412 12178 20468 12796
rect 20412 12126 20414 12178
rect 20466 12126 20468 12178
rect 20412 12114 20468 12126
rect 20524 11396 20580 12908
rect 20860 12962 20916 14028
rect 21308 14084 21364 14094
rect 21308 13858 21364 14028
rect 21308 13806 21310 13858
rect 21362 13806 21364 13858
rect 21308 13794 21364 13806
rect 21476 13860 21532 14422
rect 21476 13804 21588 13860
rect 21532 13412 21588 13804
rect 21644 13524 21700 15036
rect 21924 14756 21980 15206
rect 21644 13458 21700 13468
rect 21868 14700 21980 14756
rect 21868 13412 21924 14700
rect 21980 14530 22036 14542
rect 21980 14478 21982 14530
rect 22034 14478 22036 14530
rect 21980 14420 22036 14478
rect 21980 14354 22036 14364
rect 21980 13412 22036 13422
rect 21868 13356 21980 13412
rect 21532 13346 21588 13356
rect 21980 13346 22036 13356
rect 22092 13076 22148 16716
rect 22222 16660 22278 16670
rect 22222 16322 22278 16604
rect 22484 16436 22540 16998
rect 22540 16380 22596 16436
rect 22484 16370 22596 16380
rect 22222 16270 22224 16322
rect 22276 16270 22278 16322
rect 22222 16258 22278 16270
rect 22316 15988 22372 15998
rect 22204 15876 22260 15886
rect 22204 14756 22260 15820
rect 22204 14690 22260 14700
rect 22316 14644 22372 15932
rect 22428 15316 22484 15326
rect 22428 15222 22484 15260
rect 22316 14588 22398 14644
rect 22222 14532 22278 14542
rect 22342 14532 22398 14588
rect 22222 14530 22398 14532
rect 22222 14478 22224 14530
rect 22276 14478 22398 14530
rect 22222 14476 22398 14478
rect 22222 14466 22278 14476
rect 22316 13860 22372 13870
rect 22540 13860 22596 16370
rect 22652 15438 22708 17500
rect 22764 16772 22820 17668
rect 22764 16322 22820 16716
rect 22764 16270 22766 16322
rect 22818 16270 22820 16322
rect 22764 16258 22820 16270
rect 22876 15988 22932 18060
rect 23548 17332 23604 19180
rect 23772 19170 23828 19180
rect 23772 18564 23828 18574
rect 23660 18450 23716 18462
rect 23660 18398 23662 18450
rect 23714 18398 23716 18450
rect 23660 17556 23716 18398
rect 23772 18450 23828 18508
rect 23772 18398 23774 18450
rect 23826 18398 23828 18450
rect 23772 18386 23828 18398
rect 23884 18228 23940 19964
rect 23996 19236 24052 20076
rect 23996 19142 24052 19180
rect 24108 20018 24164 20030
rect 24108 19966 24110 20018
rect 24162 19966 24164 20018
rect 24108 19796 24164 19966
rect 24108 18564 24164 19740
rect 24332 19796 24388 20076
rect 24444 20020 24500 20638
rect 24556 20132 24612 20750
rect 25340 20244 25396 21532
rect 25676 21476 25732 21486
rect 25900 21476 25956 23660
rect 26348 23154 26404 23166
rect 26348 23102 26350 23154
rect 26402 23102 26404 23154
rect 26348 22708 26404 23102
rect 26348 22642 26404 22652
rect 26460 23156 26516 23166
rect 26012 22484 26068 22522
rect 26012 22418 26068 22428
rect 26348 22372 26404 22382
rect 26460 22372 26516 23100
rect 27020 22932 27076 23830
rect 27244 23886 27246 23938
rect 27298 23886 27300 23938
rect 27132 23156 27188 23166
rect 27244 23156 27300 23886
rect 27468 23380 27524 27580
rect 27860 27412 27916 27422
rect 27860 27186 27916 27356
rect 27860 27134 27862 27186
rect 27914 27134 27916 27186
rect 27860 27122 27916 27134
rect 28140 26516 28196 27804
rect 28252 27076 28308 27086
rect 28252 26908 28308 27020
rect 28252 26852 28364 26908
rect 28308 26850 28364 26852
rect 28308 26798 28310 26850
rect 28362 26798 28364 26850
rect 28308 26786 28364 26798
rect 28140 26450 28196 26460
rect 28196 26292 28252 26302
rect 28196 26198 28252 26236
rect 28476 26292 28532 28476
rect 28588 28084 28644 34412
rect 28924 34244 28980 34254
rect 28924 34150 28980 34188
rect 29316 33290 29372 33302
rect 29148 33236 29204 33246
rect 28924 33234 29204 33236
rect 28924 33182 29150 33234
rect 29202 33182 29204 33234
rect 28924 33180 29204 33182
rect 28700 30882 28756 30894
rect 28700 30830 28702 30882
rect 28754 30830 28756 30882
rect 28700 30772 28756 30830
rect 28700 30706 28756 30716
rect 28756 29314 28812 29326
rect 28756 29262 28758 29314
rect 28810 29262 28812 29314
rect 28756 29204 28812 29262
rect 28756 29138 28812 29148
rect 28588 28018 28644 28028
rect 28812 28980 28868 28990
rect 28644 27860 28700 27870
rect 28644 27690 28700 27804
rect 28812 27858 28868 28924
rect 28812 27806 28814 27858
rect 28866 27806 28868 27858
rect 28812 27794 28868 27806
rect 28644 27638 28646 27690
rect 28698 27638 28700 27690
rect 28644 27626 28700 27638
rect 28924 26908 28980 33180
rect 29148 33170 29204 33180
rect 29316 33238 29318 33290
rect 29370 33238 29372 33290
rect 29316 33124 29372 33238
rect 29316 33058 29372 33068
rect 29184 32956 29448 32966
rect 29240 32900 29288 32956
rect 29344 32900 29392 32956
rect 29184 32890 29448 32900
rect 29260 32788 29316 32798
rect 29148 31892 29204 31902
rect 29036 31890 29204 31892
rect 29036 31838 29150 31890
rect 29202 31838 29204 31890
rect 29036 31836 29204 31838
rect 29036 31220 29092 31836
rect 29148 31826 29204 31836
rect 29260 31763 29316 32732
rect 29708 32786 29764 35196
rect 30044 34468 30100 39200
rect 31052 36482 31108 36494
rect 30716 36454 30772 36466
rect 30716 36402 30718 36454
rect 30770 36402 30772 36454
rect 30716 36372 30772 36402
rect 30492 34916 30548 34926
rect 30492 34822 30548 34860
rect 30044 34402 30100 34412
rect 29820 33796 29876 33806
rect 29820 33346 29876 33740
rect 30586 33460 30642 33470
rect 30586 33366 30642 33404
rect 29820 33294 29822 33346
rect 29874 33294 29876 33346
rect 29820 33282 29876 33294
rect 30062 33236 30118 33246
rect 29708 32734 29710 32786
rect 29762 32734 29764 32786
rect 29708 32722 29764 32734
rect 29932 33234 30118 33236
rect 29932 33182 30064 33234
rect 30116 33182 30118 33234
rect 29932 33180 30118 33182
rect 29260 31711 29262 31763
rect 29314 31711 29316 31763
rect 29484 32340 29540 32350
rect 29484 31778 29540 32284
rect 29484 31726 29486 31778
rect 29538 31726 29540 31778
rect 29484 31714 29540 31726
rect 29260 31699 29316 31711
rect 29184 31388 29448 31398
rect 29240 31332 29288 31388
rect 29344 31332 29392 31388
rect 29184 31322 29448 31332
rect 29036 31164 29204 31220
rect 29036 30996 29092 31006
rect 29036 30902 29092 30940
rect 29148 29988 29204 31164
rect 29932 31108 29988 33180
rect 30062 33170 30118 33180
rect 30156 33012 30212 33022
rect 29260 31052 29988 31108
rect 30044 32788 30100 32798
rect 29260 30994 29316 31052
rect 30044 30996 30100 32732
rect 29260 30942 29262 30994
rect 29314 30942 29316 30994
rect 29260 30930 29316 30942
rect 29540 30940 30100 30996
rect 29540 30882 29596 30940
rect 29540 30830 29542 30882
rect 29594 30830 29596 30882
rect 29540 30818 29596 30830
rect 30156 30772 30212 32956
rect 29708 30716 30212 30772
rect 30380 32004 30436 32014
rect 30380 31021 30436 31948
rect 30716 31108 30772 36316
rect 31052 36430 31054 36482
rect 31106 36430 31108 36482
rect 30940 35924 30996 35934
rect 31052 35924 31108 36430
rect 30940 35922 31108 35924
rect 30940 35870 30942 35922
rect 30994 35870 31108 35922
rect 30940 35868 31108 35870
rect 30940 35858 30996 35868
rect 30940 35700 30996 35710
rect 30828 34020 30884 34030
rect 30828 33926 30884 33964
rect 30828 33460 30884 33470
rect 30828 33346 30884 33404
rect 30828 33294 30830 33346
rect 30882 33294 30884 33346
rect 30828 32116 30884 33294
rect 30940 32900 30996 35644
rect 31164 35140 31220 39200
rect 31388 36260 31444 36270
rect 31388 36166 31444 36204
rect 31276 35700 31332 35710
rect 31276 35606 31332 35644
rect 31724 35698 31780 35710
rect 32284 35700 32340 39200
rect 33180 36594 33236 36606
rect 33180 36542 33182 36594
rect 33234 36542 33236 36594
rect 31724 35646 31726 35698
rect 31778 35646 31780 35698
rect 31164 35074 31220 35084
rect 31052 34914 31108 34926
rect 31052 34862 31054 34914
rect 31106 34862 31108 34914
rect 31052 33572 31108 34862
rect 31724 34356 31780 35646
rect 31948 35644 32340 35700
rect 32508 36454 32564 36466
rect 32508 36402 32510 36454
rect 32562 36402 32564 36454
rect 31836 34916 31892 34926
rect 31836 34822 31892 34860
rect 31724 34300 31892 34356
rect 31052 33506 31108 33516
rect 31164 34132 31220 34142
rect 30940 32834 30996 32844
rect 31164 32788 31220 34076
rect 31612 34130 31668 34142
rect 31612 34078 31614 34130
rect 31666 34078 31668 34130
rect 31332 33908 31388 33918
rect 31332 33402 31388 33852
rect 31332 33350 31334 33402
rect 31386 33350 31388 33402
rect 31332 33338 31388 33350
rect 31612 33572 31668 34078
rect 31724 34132 31780 34142
rect 31724 34038 31780 34076
rect 31612 33348 31668 33516
rect 31724 33348 31780 33358
rect 31612 33346 31780 33348
rect 31612 33294 31726 33346
rect 31778 33294 31780 33346
rect 31612 33292 31780 33294
rect 31500 33236 31556 33246
rect 31500 33234 31668 33236
rect 31500 33182 31502 33234
rect 31554 33182 31668 33234
rect 31500 33180 31668 33182
rect 31500 33170 31556 33180
rect 31164 32722 31220 32732
rect 31444 32676 31500 32686
rect 31444 32582 31500 32620
rect 30828 32050 30884 32060
rect 30940 32562 30996 32574
rect 30940 32510 30942 32562
rect 30994 32510 30996 32562
rect 30940 32340 30996 32510
rect 31164 32564 31220 32574
rect 31164 32562 31332 32564
rect 31164 32510 31166 32562
rect 31218 32510 31332 32562
rect 31164 32508 31332 32510
rect 31164 32498 31220 32508
rect 30716 31042 30772 31052
rect 30380 30969 30382 31021
rect 30434 30969 30436 31021
rect 29484 30212 29540 30222
rect 29484 30118 29540 30156
rect 29596 30212 29652 30222
rect 29708 30212 29764 30716
rect 29596 30210 29764 30212
rect 29596 30158 29598 30210
rect 29650 30158 29764 30210
rect 29596 30156 29764 30158
rect 29876 30212 29932 30222
rect 29596 30146 29652 30156
rect 29876 30118 29932 30156
rect 29148 29932 29876 29988
rect 29184 29820 29448 29830
rect 29240 29764 29288 29820
rect 29344 29764 29392 29820
rect 29184 29754 29448 29764
rect 29092 29652 29148 29662
rect 29092 29558 29148 29596
rect 29260 29540 29316 29550
rect 29260 29482 29316 29484
rect 29260 29430 29262 29482
rect 29314 29430 29316 29482
rect 29260 29418 29316 29430
rect 29372 29428 29428 29466
rect 29372 29362 29428 29372
rect 29036 29204 29092 29214
rect 29036 28084 29092 29148
rect 29372 29204 29428 29214
rect 29260 28644 29316 28654
rect 29372 28644 29428 29148
rect 29260 28642 29428 28644
rect 29260 28590 29262 28642
rect 29314 28590 29428 28642
rect 29260 28588 29428 28590
rect 29596 28644 29652 28654
rect 29260 28578 29316 28588
rect 29596 28550 29652 28588
rect 29184 28252 29448 28262
rect 29240 28196 29288 28252
rect 29344 28196 29392 28252
rect 29184 28186 29448 28196
rect 29204 28084 29260 28094
rect 29036 28082 29316 28084
rect 29036 28030 29206 28082
rect 29258 28030 29316 28082
rect 29036 28028 29316 28030
rect 29204 28018 29316 28028
rect 29260 27198 29316 28018
rect 29652 27748 29708 27758
rect 29596 27692 29652 27748
rect 29596 27654 29708 27692
rect 29260 27186 29372 27198
rect 29260 27134 29318 27186
rect 29370 27134 29372 27186
rect 29260 27132 29372 27134
rect 29316 27122 29372 27132
rect 29596 26908 29652 27654
rect 28476 26226 28532 26236
rect 28588 26852 28980 26908
rect 29036 26852 29652 26908
rect 29820 26908 29876 29932
rect 30380 29428 30436 30969
rect 30940 29652 30996 32284
rect 30940 29586 30996 29596
rect 30380 29362 30436 29372
rect 30156 29316 30212 29326
rect 29932 29314 30212 29316
rect 29932 29262 30158 29314
rect 30210 29262 30212 29314
rect 29932 29260 30212 29262
rect 29932 28084 29988 29260
rect 30156 29250 30212 29260
rect 30604 28980 30660 28990
rect 30212 28644 30268 28654
rect 30156 28642 30268 28644
rect 30156 28590 30214 28642
rect 30266 28590 30268 28642
rect 30156 28578 30268 28590
rect 30044 28084 30100 28094
rect 29932 28082 30100 28084
rect 29932 28030 30046 28082
rect 30098 28030 30100 28082
rect 29932 28028 30100 28030
rect 30044 28018 30100 28028
rect 30156 27748 30212 28578
rect 30380 28532 30436 28542
rect 30156 27682 30212 27692
rect 30268 28474 30324 28486
rect 30268 28422 30270 28474
rect 30322 28422 30324 28474
rect 30268 26908 30324 28422
rect 30380 27858 30436 28476
rect 30380 27806 30382 27858
rect 30434 27806 30436 27858
rect 30380 27794 30436 27806
rect 30492 27860 30548 27870
rect 30604 27860 30660 28924
rect 30958 28868 31014 28878
rect 31276 28868 31332 32508
rect 30958 28866 31332 28868
rect 30958 28814 30960 28866
rect 31012 28814 31332 28866
rect 30958 28812 31332 28814
rect 31388 32452 31444 32462
rect 30958 28802 31014 28812
rect 31388 28756 31444 32396
rect 31500 31890 31556 31902
rect 31500 31838 31502 31890
rect 31554 31838 31556 31890
rect 31500 31780 31556 31838
rect 31500 31714 31556 31724
rect 31612 30100 31668 33180
rect 31724 32004 31780 33292
rect 31836 32676 31892 34300
rect 31948 32788 32004 35644
rect 32060 35474 32116 35486
rect 32060 35422 32062 35474
rect 32114 35422 32116 35474
rect 32060 34356 32116 35422
rect 32508 35252 32564 36402
rect 33068 36260 33124 36270
rect 33068 35725 33124 36204
rect 33068 35673 33070 35725
rect 33122 35673 33124 35725
rect 33068 35661 33124 35673
rect 32508 35196 33012 35252
rect 32956 34356 33012 35196
rect 33180 35028 33236 36542
rect 33180 34962 33236 34972
rect 32060 34300 32564 34356
rect 32172 34132 32228 34142
rect 32060 34020 32116 34030
rect 32060 33926 32116 33964
rect 32172 33460 32228 34076
rect 32172 33394 32228 33404
rect 32508 33458 32564 34300
rect 32508 33406 32510 33458
rect 32562 33406 32564 33458
rect 32508 33394 32564 33406
rect 32620 34300 33012 34356
rect 31948 32732 32116 32788
rect 31836 32610 31892 32620
rect 31948 32562 32004 32574
rect 31948 32510 31950 32562
rect 32002 32510 32004 32562
rect 31948 32340 32004 32510
rect 31948 32274 32004 32284
rect 31724 30434 31780 31948
rect 31724 30382 31726 30434
rect 31778 30382 31780 30434
rect 31724 30370 31780 30382
rect 31612 30044 31892 30100
rect 31276 28700 31444 28756
rect 30716 28644 30772 28654
rect 31276 28644 31332 28700
rect 30716 28642 31332 28644
rect 30716 28590 30718 28642
rect 30770 28590 31332 28642
rect 30716 28588 31332 28590
rect 30716 28578 30772 28588
rect 31556 28586 31612 28598
rect 31388 28532 31444 28542
rect 30828 28530 31444 28532
rect 30828 28478 31390 28530
rect 31442 28478 31444 28530
rect 30828 28476 31444 28478
rect 30716 27860 30772 27870
rect 30604 27858 30772 27860
rect 30604 27806 30718 27858
rect 30770 27806 30772 27858
rect 30604 27804 30772 27806
rect 30492 27298 30548 27804
rect 30716 27794 30772 27804
rect 30828 27748 30884 28476
rect 31388 28466 31444 28476
rect 31556 28534 31558 28586
rect 31610 28534 31612 28586
rect 31556 28196 31612 28534
rect 30996 28140 31612 28196
rect 30996 27970 31052 28140
rect 30996 27918 30998 27970
rect 31050 27918 31052 27970
rect 30996 27906 31052 27918
rect 31500 27860 31556 27870
rect 31388 27858 31556 27860
rect 31388 27806 31502 27858
rect 31554 27806 31556 27858
rect 31388 27804 31556 27806
rect 30828 27692 30996 27748
rect 30492 27246 30494 27298
rect 30546 27246 30548 27298
rect 30492 27234 30548 27246
rect 30716 27636 30772 27646
rect 30716 26908 30772 27580
rect 30828 27076 30884 27114
rect 30828 27010 30884 27020
rect 29820 26852 30100 26908
rect 30268 26852 30548 26908
rect 30716 26852 30884 26908
rect 28364 26180 28420 26190
rect 27916 25620 27972 25630
rect 27692 25506 27748 25518
rect 27692 25454 27694 25506
rect 27746 25454 27748 25506
rect 27692 24498 27748 25454
rect 27916 25338 27972 25564
rect 28364 25506 28420 26124
rect 28588 25620 28644 26852
rect 28588 25554 28644 25564
rect 28364 25454 28366 25506
rect 28418 25454 28420 25506
rect 28364 25442 28420 25454
rect 27916 25286 27918 25338
rect 27970 25286 27972 25338
rect 27916 25274 27972 25286
rect 28028 25284 28084 25294
rect 28028 25172 28084 25228
rect 27692 24446 27694 24498
rect 27746 24446 27748 24498
rect 27692 24434 27748 24446
rect 27916 25116 28084 25172
rect 27580 23940 27636 23950
rect 27580 23846 27636 23884
rect 27804 23380 27860 23390
rect 27468 23324 27636 23380
rect 27188 23100 27300 23156
rect 27468 23154 27524 23166
rect 27468 23102 27470 23154
rect 27522 23102 27524 23154
rect 27132 23062 27188 23100
rect 27468 22932 27524 23102
rect 27580 23044 27636 23324
rect 27804 23210 27860 23324
rect 27804 23158 27806 23210
rect 27858 23158 27860 23210
rect 27804 23146 27860 23158
rect 27580 22988 27748 23044
rect 27020 22876 27524 22932
rect 26348 22370 26516 22372
rect 26124 22314 26180 22326
rect 25676 21474 25956 21476
rect 25676 21422 25678 21474
rect 25730 21422 25956 21474
rect 25676 21420 25956 21422
rect 26012 22260 26068 22270
rect 25676 21410 25732 21420
rect 26012 21252 26068 22204
rect 25564 21196 26068 21252
rect 26124 22262 26126 22314
rect 26178 22262 26180 22314
rect 26124 21586 26180 22262
rect 26348 22318 26350 22370
rect 26402 22318 26516 22370
rect 26348 22316 26516 22318
rect 26348 21700 26404 22316
rect 26796 21700 26852 21710
rect 26348 21644 26628 21700
rect 26124 21534 26126 21586
rect 26178 21534 26180 21586
rect 25564 20802 25620 21196
rect 25788 21028 25844 21038
rect 25564 20750 25566 20802
rect 25618 20750 25620 20802
rect 25564 20738 25620 20750
rect 25676 20970 25732 20982
rect 25676 20918 25678 20970
rect 25730 20918 25732 20970
rect 24556 20066 24612 20076
rect 25228 20188 25396 20244
rect 25228 20020 25284 20188
rect 24444 19954 24500 19964
rect 25004 19964 25284 20020
rect 25452 20018 25508 20030
rect 25452 19966 25454 20018
rect 25506 19966 25508 20018
rect 24444 19796 24500 19806
rect 24332 19794 24500 19796
rect 24332 19742 24446 19794
rect 24498 19742 24500 19794
rect 24332 19740 24500 19742
rect 24332 19572 24388 19740
rect 24444 19730 24500 19740
rect 24522 19628 24786 19638
rect 24578 19572 24626 19628
rect 24682 19572 24730 19628
rect 24522 19562 24786 19572
rect 24332 19506 24388 19516
rect 25004 19346 25060 19964
rect 25284 19794 25340 19806
rect 25284 19742 25286 19794
rect 25338 19742 25340 19794
rect 25284 19460 25340 19742
rect 25284 19394 25340 19404
rect 25004 19294 25006 19346
rect 25058 19294 25060 19346
rect 25004 19282 25060 19294
rect 24780 19234 24836 19246
rect 25340 19236 25396 19246
rect 24780 19182 24782 19234
rect 24834 19182 24836 19234
rect 25228 19234 25396 19236
rect 24276 19124 24332 19134
rect 24780 19124 24836 19182
rect 24276 19122 24836 19124
rect 24276 19070 24278 19122
rect 24330 19070 24836 19122
rect 24276 19068 24836 19070
rect 24276 19058 24332 19068
rect 24108 18450 24164 18508
rect 24108 18398 24110 18450
rect 24162 18398 24164 18450
rect 24108 18386 24164 18398
rect 24332 18450 24388 18462
rect 24332 18398 24334 18450
rect 24386 18398 24388 18450
rect 23884 18172 24164 18228
rect 23660 17490 23716 17500
rect 23884 17666 23940 17678
rect 23884 17614 23886 17666
rect 23938 17614 23940 17666
rect 23884 17332 23940 17614
rect 23548 17276 23940 17332
rect 23044 17108 23100 17118
rect 23044 17014 23100 17052
rect 23548 16882 23604 17276
rect 23772 17108 23828 17118
rect 23548 16830 23550 16882
rect 23602 16830 23604 16882
rect 23548 16818 23604 16830
rect 23660 16996 23716 17006
rect 23660 16882 23716 16940
rect 23660 16830 23662 16882
rect 23714 16830 23716 16882
rect 23660 16818 23716 16830
rect 23100 16100 23156 16110
rect 23156 16044 23380 16100
rect 23100 16006 23156 16044
rect 22876 15922 22932 15932
rect 23324 15538 23380 16044
rect 23492 15876 23548 15886
rect 23772 15876 23828 17052
rect 23940 16658 23996 16670
rect 23940 16606 23942 16658
rect 23994 16606 23996 16658
rect 23940 16100 23996 16606
rect 23940 16034 23996 16044
rect 23772 15820 23996 15876
rect 23492 15782 23548 15820
rect 23324 15486 23326 15538
rect 23378 15486 23380 15538
rect 23324 15474 23380 15486
rect 23940 15538 23996 15820
rect 23940 15486 23942 15538
rect 23994 15486 23996 15538
rect 23940 15474 23996 15486
rect 22652 15426 22726 15438
rect 22652 15374 22672 15426
rect 22724 15374 22726 15426
rect 22652 15372 22726 15374
rect 22670 15362 22726 15372
rect 22988 15314 23044 15326
rect 22988 15262 22990 15314
rect 23042 15262 23044 15314
rect 22988 15148 23044 15262
rect 22876 15092 23044 15148
rect 23436 15316 23492 15326
rect 22764 14980 22820 14990
rect 22652 14532 22708 14542
rect 22652 14438 22708 14476
rect 22764 14362 22820 14924
rect 22764 14310 22766 14362
rect 22818 14310 22820 14362
rect 22764 14298 22820 14310
rect 22876 13972 22932 15092
rect 23324 14532 23380 14542
rect 23436 14532 23492 15260
rect 24108 15148 24164 18172
rect 24332 18116 24388 18398
rect 24612 18452 24668 18462
rect 24612 18358 24668 18396
rect 24780 18228 24836 19068
rect 25004 19178 25060 19190
rect 25004 19126 25006 19178
rect 25058 19126 25060 19178
rect 25004 18676 25060 19126
rect 25004 18610 25060 18620
rect 25228 19182 25342 19234
rect 25394 19182 25396 19234
rect 25228 19180 25396 19182
rect 25228 18340 25284 19180
rect 25340 19170 25396 19180
rect 25452 19236 25508 19966
rect 25452 19170 25508 19180
rect 25564 18676 25620 18686
rect 25564 18450 25620 18620
rect 25564 18398 25566 18450
rect 25618 18398 25620 18450
rect 25564 18386 25620 18398
rect 25228 18274 25284 18284
rect 24780 18162 24836 18172
rect 25564 18228 25620 18238
rect 24332 18050 24388 18060
rect 24522 18060 24786 18070
rect 24578 18004 24626 18060
rect 24682 18004 24730 18060
rect 24522 17994 24786 18004
rect 24332 17892 24388 17912
rect 24332 17834 24388 17836
rect 24332 17782 24334 17834
rect 24386 17782 24388 17834
rect 24220 17666 24276 17678
rect 24220 17614 24222 17666
rect 24274 17614 24276 17666
rect 24220 17556 24276 17614
rect 24220 17490 24276 17500
rect 24332 16996 24388 17782
rect 25172 17668 25228 17678
rect 25172 17574 25228 17612
rect 25452 17668 25508 17678
rect 25452 17574 25508 17612
rect 25564 17666 25620 18172
rect 25676 18116 25732 20918
rect 25788 20802 25844 20972
rect 25788 20750 25790 20802
rect 25842 20750 25844 20802
rect 25788 20254 25844 20750
rect 26124 20804 26180 21534
rect 26572 21625 26628 21644
rect 26572 21573 26574 21625
rect 26626 21588 26628 21625
rect 26626 21573 26740 21588
rect 26572 21532 26740 21573
rect 26124 20710 26180 20748
rect 26236 21474 26292 21486
rect 26236 21422 26238 21474
rect 26290 21422 26292 21474
rect 26236 20692 26292 21422
rect 26236 20626 26292 20636
rect 26460 21028 26516 21038
rect 26460 20578 26516 20972
rect 26460 20526 26462 20578
rect 26514 20526 26516 20578
rect 25788 20242 25900 20254
rect 25788 20190 25846 20242
rect 25898 20190 25900 20242
rect 25788 20188 25900 20190
rect 25844 20178 25900 20188
rect 26460 20020 26516 20526
rect 26236 19964 26516 20020
rect 25900 19234 25956 19246
rect 25900 19182 25902 19234
rect 25954 19182 25956 19234
rect 25900 19124 25956 19182
rect 25900 19058 25956 19068
rect 25788 18508 25956 18564
rect 25788 18340 25844 18508
rect 25900 18506 25956 18508
rect 25900 18454 25902 18506
rect 25954 18454 25956 18506
rect 25900 18442 25956 18454
rect 26236 18450 26292 19964
rect 26572 19236 26628 19246
rect 26236 18398 26238 18450
rect 26290 18398 26292 18450
rect 26236 18386 26292 18398
rect 26348 19178 26404 19190
rect 26348 19126 26350 19178
rect 26402 19126 26404 19178
rect 25788 18274 25844 18284
rect 25900 18340 25956 18350
rect 25900 18338 26180 18340
rect 25900 18286 25902 18338
rect 25954 18286 26180 18338
rect 25900 18284 26180 18286
rect 25900 18274 25956 18284
rect 25676 18060 25956 18116
rect 25564 17614 25566 17666
rect 25618 17614 25620 17666
rect 25900 17666 25956 18060
rect 25564 17602 25620 17614
rect 25732 17610 25788 17622
rect 25732 17558 25734 17610
rect 25786 17558 25788 17610
rect 25732 17220 25788 17558
rect 25900 17614 25902 17666
rect 25954 17614 25956 17666
rect 25900 17444 25956 17614
rect 25900 17378 25956 17388
rect 26012 17780 26068 17790
rect 26012 17220 26068 17724
rect 25732 17154 25788 17164
rect 25900 17164 26068 17220
rect 24332 16930 24388 16940
rect 25564 16996 25620 17006
rect 25564 16882 25620 16940
rect 25564 16830 25566 16882
rect 25618 16830 25620 16882
rect 25732 16996 25788 17006
rect 25732 16938 25788 16940
rect 25732 16886 25734 16938
rect 25786 16886 25788 16938
rect 25900 16994 25956 17164
rect 25900 16942 25902 16994
rect 25954 16942 25956 16994
rect 25900 16930 25956 16942
rect 25732 16874 25788 16886
rect 26012 16884 26068 16894
rect 25564 16818 25620 16830
rect 26012 16790 26068 16828
rect 24522 16492 24786 16502
rect 24578 16436 24626 16492
rect 24682 16436 24730 16492
rect 24522 16426 24786 16436
rect 24575 16100 24631 16110
rect 24575 16006 24631 16044
rect 25452 16100 25508 16110
rect 25452 16006 25508 16044
rect 24332 15988 24388 15998
rect 24332 15986 24500 15988
rect 24332 15934 24334 15986
rect 24386 15934 24500 15986
rect 24332 15932 24500 15934
rect 24332 15922 24388 15932
rect 24444 15540 24500 15932
rect 25508 15540 25564 15550
rect 26012 15540 26068 15550
rect 24444 15484 25172 15540
rect 24388 15316 24444 15326
rect 24388 15202 24444 15260
rect 24388 15150 24390 15202
rect 24442 15150 24444 15202
rect 24108 15092 24276 15148
rect 23324 14530 23492 14532
rect 22876 13906 22932 13916
rect 23100 14474 23156 14486
rect 23100 14422 23102 14474
rect 23154 14422 23156 14474
rect 23324 14478 23326 14530
rect 23378 14478 23492 14530
rect 23324 14476 23492 14478
rect 23324 14466 23380 14476
rect 23100 14420 23156 14422
rect 22316 13858 22596 13860
rect 22316 13806 22318 13858
rect 22370 13806 22596 13858
rect 22316 13804 22596 13806
rect 22316 13794 22372 13804
rect 22988 13748 23044 13758
rect 22652 13746 23044 13748
rect 22484 13690 22540 13702
rect 22484 13638 22486 13690
rect 22538 13638 22540 13690
rect 21980 13020 22148 13076
rect 22316 13412 22372 13422
rect 20860 12910 20862 12962
rect 20914 12910 20916 12962
rect 20860 12898 20916 12910
rect 21308 12964 21364 12974
rect 21308 12870 21364 12908
rect 21084 11844 21140 11854
rect 19860 11004 20124 11014
rect 19916 10948 19964 11004
rect 20020 10948 20068 11004
rect 19860 10938 20124 10948
rect 17500 10834 17612 10836
rect 17500 10782 17558 10834
rect 17610 10782 17612 10834
rect 17500 10770 17612 10782
rect 18900 10836 19012 10846
rect 20524 10836 20580 11340
rect 20636 11396 20692 11406
rect 21084 11396 21140 11788
rect 21980 11508 22036 13020
rect 22184 12906 22240 12918
rect 22184 12854 22186 12906
rect 22238 12854 22240 12906
rect 22184 12852 22240 12854
rect 22184 12786 22240 12796
rect 22316 12292 22372 13356
rect 22484 13198 22540 13638
rect 22428 13186 22540 13198
rect 22428 13134 22430 13186
rect 22482 13134 22540 13186
rect 22428 13132 22540 13134
rect 22652 13694 22990 13746
rect 23042 13694 23044 13746
rect 22652 13692 23044 13694
rect 22428 13122 22484 13132
rect 21308 11396 21364 11406
rect 20636 11394 21364 11396
rect 20636 11342 20638 11394
rect 20690 11342 21310 11394
rect 21362 11342 21364 11394
rect 20636 11340 21364 11342
rect 20636 11330 20692 11340
rect 21308 11330 21364 11340
rect 18900 10834 19684 10836
rect 18900 10782 18902 10834
rect 18954 10782 19684 10834
rect 18900 10780 19684 10782
rect 18900 10770 18956 10780
rect 17500 9828 17556 10770
rect 19292 10612 19348 10622
rect 19292 10518 19348 10556
rect 19628 10610 19684 10780
rect 20524 10770 20580 10780
rect 21028 10836 21084 10846
rect 21028 10742 21084 10780
rect 19628 10558 19630 10610
rect 19682 10558 19684 10610
rect 19628 9940 19684 10558
rect 19740 10612 19796 10622
rect 19740 10518 19796 10556
rect 20076 10386 20132 10398
rect 20076 10334 20078 10386
rect 20130 10334 20132 10386
rect 20076 10052 20132 10334
rect 20076 9996 20244 10052
rect 19628 9884 19796 9940
rect 17164 9826 17556 9828
rect 17164 9774 17502 9826
rect 17554 9774 17556 9826
rect 17164 9772 17556 9774
rect 16940 9604 16996 9614
rect 16940 9042 16996 9548
rect 16940 8990 16942 9042
rect 16994 8990 16996 9042
rect 16940 8978 16996 8990
rect 17164 8046 17220 9772
rect 17500 9762 17556 9772
rect 17556 9604 17612 9614
rect 17556 9266 17612 9548
rect 18956 9602 19012 9614
rect 18956 9550 18958 9602
rect 19010 9550 19012 9602
rect 17556 9214 17558 9266
rect 17610 9214 17612 9266
rect 17556 9202 17612 9214
rect 18228 9268 18284 9278
rect 18228 9174 18284 9212
rect 18732 8820 18788 8830
rect 18732 8370 18788 8764
rect 18732 8318 18734 8370
rect 18786 8318 18788 8370
rect 18732 8306 18788 8318
rect 17948 8258 18004 8270
rect 17948 8206 17950 8258
rect 18002 8206 18004 8258
rect 16604 7746 16660 7756
rect 17108 8036 17220 8046
rect 17108 8034 17164 8036
rect 17108 7982 17110 8034
rect 17162 7982 17164 8034
rect 17108 7980 17164 7982
rect 17108 7942 17220 7980
rect 17780 8036 17836 8046
rect 17948 8036 18004 8206
rect 17836 7980 18004 8036
rect 17780 7942 17836 7980
rect 16716 7474 16772 7486
rect 16716 7422 16718 7474
rect 16770 7422 16772 7474
rect 16436 7252 16492 7262
rect 16436 7250 16548 7252
rect 16436 7198 16438 7250
rect 16490 7198 16548 7250
rect 16436 7186 16548 7198
rect 16268 6692 16324 6702
rect 15484 5030 15540 5068
rect 15372 4386 15428 4396
rect 15820 4450 15876 6076
rect 16100 6634 16156 6646
rect 16100 6582 16102 6634
rect 16154 6582 16156 6634
rect 16268 6598 16324 6636
rect 16492 6690 16548 7186
rect 16716 6916 16772 7422
rect 16716 6850 16772 6860
rect 16940 7474 16996 7486
rect 16940 7422 16942 7474
rect 16994 7422 16996 7474
rect 16492 6638 16494 6690
rect 16546 6638 16548 6690
rect 16492 6626 16548 6638
rect 16100 6132 16156 6582
rect 16940 6468 16996 7422
rect 17108 7476 17164 7942
rect 18956 7700 19012 9550
rect 19740 9268 19796 9884
rect 20076 9826 20132 9838
rect 20076 9774 20078 9826
rect 20130 9774 20132 9826
rect 20076 9604 20132 9774
rect 20076 9538 20132 9548
rect 19860 9436 20124 9446
rect 19916 9380 19964 9436
rect 20020 9380 20068 9436
rect 19860 9370 20124 9380
rect 20188 9268 20244 9996
rect 20468 9940 20524 9950
rect 20468 9604 20524 9884
rect 20468 9538 20524 9548
rect 21868 9828 21924 9838
rect 19740 9212 20020 9268
rect 19180 8820 19236 8830
rect 19180 8726 19236 8764
rect 19964 8036 20020 9212
rect 20076 9212 20244 9268
rect 20076 8260 20132 9212
rect 20636 9042 20692 9054
rect 20636 8990 20638 9042
rect 20690 8990 20692 9042
rect 20636 8428 20692 8990
rect 20076 8194 20132 8204
rect 20524 8372 20692 8428
rect 21868 8484 21924 9772
rect 21980 9268 22036 11452
rect 22204 12290 22372 12292
rect 22204 12238 22318 12290
rect 22370 12238 22372 12290
rect 22204 12236 22372 12238
rect 22204 11406 22260 12236
rect 22316 12226 22372 12236
rect 22428 11620 22484 11630
rect 22652 11620 22708 13692
rect 22988 13682 23044 13692
rect 22876 13524 22932 13534
rect 22876 13074 22932 13468
rect 22876 13022 22878 13074
rect 22930 13022 22932 13074
rect 22876 13010 22932 13022
rect 22988 13412 23044 13422
rect 22988 12947 23044 13356
rect 22988 12895 22990 12947
rect 23042 12895 23044 12947
rect 23100 13188 23156 14364
rect 23230 13748 23286 13758
rect 23230 13654 23286 13692
rect 23100 12964 23156 13132
rect 23100 12898 23156 12908
rect 23212 13300 23268 13310
rect 23212 12962 23268 13244
rect 23212 12910 23214 12962
rect 23266 12910 23268 12962
rect 22988 12883 23044 12895
rect 22428 11618 22708 11620
rect 22428 11566 22430 11618
rect 22482 11566 22708 11618
rect 22428 11564 22708 11566
rect 22764 12852 22820 12862
rect 22764 12404 22820 12796
rect 22932 12404 22988 12414
rect 22764 12402 22988 12404
rect 22764 12350 22934 12402
rect 22986 12350 22988 12402
rect 22764 12348 22988 12350
rect 22428 11554 22484 11564
rect 22184 11394 22260 11406
rect 22184 11342 22186 11394
rect 22238 11342 22260 11394
rect 22184 11340 22260 11342
rect 22764 11508 22820 12348
rect 22932 12338 22988 12348
rect 23212 11844 23268 12910
rect 23324 13188 23380 13198
rect 23324 12414 23380 13132
rect 23436 12852 23492 14476
rect 24052 14308 24108 14318
rect 24052 14306 24164 14308
rect 24052 14254 24054 14306
rect 24106 14254 24164 14306
rect 24052 14242 24164 14254
rect 23548 14084 23604 14094
rect 23548 12962 23604 14028
rect 23940 13972 23996 13982
rect 23940 13878 23996 13916
rect 23772 13748 23828 13758
rect 23772 13654 23828 13692
rect 24108 13188 24164 14242
rect 24108 13122 24164 13132
rect 23548 12910 23550 12962
rect 23602 12910 23604 12962
rect 23548 12898 23604 12910
rect 23436 12786 23492 12796
rect 24220 12740 24276 15092
rect 24388 14644 24444 15150
rect 24522 14924 24786 14934
rect 24578 14868 24626 14924
rect 24682 14868 24730 14924
rect 24522 14858 24786 14868
rect 24500 14644 24556 14654
rect 24388 14642 24556 14644
rect 24388 14590 24502 14642
rect 24554 14590 24556 14642
rect 24388 14588 24556 14590
rect 24500 14578 24556 14588
rect 25116 14530 25172 15484
rect 25508 15538 26068 15540
rect 25508 15486 25510 15538
rect 25562 15486 26014 15538
rect 26066 15486 26068 15538
rect 25508 15484 26068 15486
rect 25508 15474 25564 15484
rect 26012 15474 26068 15484
rect 25116 14478 25118 14530
rect 25170 14478 25172 14530
rect 25116 14466 25172 14478
rect 25340 15314 25396 15326
rect 25340 15262 25342 15314
rect 25394 15262 25396 15314
rect 25340 14532 25396 15262
rect 26124 15148 26180 18284
rect 26348 17332 26404 19126
rect 26460 18228 26516 18238
rect 26460 17638 26516 18172
rect 26572 17780 26628 19180
rect 26684 19066 26740 21532
rect 26796 21586 26852 21644
rect 26796 21534 26798 21586
rect 26850 21534 26852 21586
rect 26796 21522 26852 21534
rect 27132 21588 27188 21598
rect 27132 21494 27188 21532
rect 26908 21028 26964 21038
rect 26908 19236 26964 20972
rect 27468 21028 27524 22876
rect 27580 22484 27636 22494
rect 27580 22370 27636 22428
rect 27580 22318 27582 22370
rect 27634 22318 27636 22370
rect 27580 21586 27636 22318
rect 27580 21534 27582 21586
rect 27634 21534 27636 21586
rect 27580 21522 27636 21534
rect 27692 21364 27748 22988
rect 27916 23042 27972 25116
rect 29036 24948 29092 26852
rect 29184 26684 29448 26694
rect 29240 26628 29288 26684
rect 29344 26628 29392 26684
rect 29184 26618 29448 26628
rect 29596 25564 29876 25620
rect 29428 25508 29484 25518
rect 29428 25338 29484 25452
rect 29596 25506 29652 25564
rect 29596 25454 29598 25506
rect 29650 25454 29652 25506
rect 29596 25442 29652 25454
rect 29428 25286 29430 25338
rect 29482 25286 29484 25338
rect 29428 25284 29484 25286
rect 29428 25228 29652 25284
rect 29184 25116 29448 25126
rect 29240 25060 29288 25116
rect 29344 25060 29392 25116
rect 29184 25050 29448 25060
rect 29596 24948 29652 25228
rect 29820 25060 29876 25564
rect 29932 25508 29988 25518
rect 29932 25414 29988 25452
rect 29820 24994 29876 25004
rect 29036 24882 29092 24892
rect 29260 24892 29652 24948
rect 29260 24766 29316 24892
rect 29036 24722 29092 24734
rect 29036 24670 29038 24722
rect 29090 24670 29092 24722
rect 29260 24714 29262 24766
rect 29314 24714 29316 24766
rect 29260 24702 29316 24714
rect 29820 24724 29876 24734
rect 29036 24164 29092 24670
rect 29820 24630 29876 24668
rect 28140 24106 28196 24118
rect 28140 24054 28142 24106
rect 28194 24054 28196 24106
rect 28028 23492 28084 23502
rect 28028 23154 28084 23436
rect 28028 23102 28030 23154
rect 28082 23102 28084 23154
rect 28028 23090 28084 23102
rect 27916 22990 27918 23042
rect 27970 22990 27972 23042
rect 27916 22978 27972 22990
rect 28140 22820 28196 24054
rect 28924 24108 29036 24164
rect 28252 23940 28308 23950
rect 28252 23846 28308 23884
rect 28588 23940 28644 23950
rect 28588 23938 28868 23940
rect 28588 23886 28590 23938
rect 28642 23886 28868 23938
rect 28588 23884 28868 23886
rect 28588 23874 28644 23884
rect 28644 23492 28700 23502
rect 28644 23378 28700 23436
rect 28644 23326 28646 23378
rect 28698 23326 28700 23378
rect 28644 23314 28700 23326
rect 28812 22820 28868 23884
rect 28924 23492 28980 24108
rect 29036 24098 29092 24108
rect 29372 24610 29428 24622
rect 29372 24558 29374 24610
rect 29426 24558 29428 24610
rect 28924 23426 28980 23436
rect 29036 23940 29092 23950
rect 29036 23380 29092 23884
rect 29372 23940 29428 24558
rect 29652 24164 29708 24174
rect 29652 24050 29708 24108
rect 29652 23998 29654 24050
rect 29706 23998 29708 24050
rect 29652 23986 29708 23998
rect 29820 24052 29876 24062
rect 29372 23874 29428 23884
rect 29184 23548 29448 23558
rect 29240 23492 29288 23548
rect 29344 23492 29392 23548
rect 29184 23482 29448 23492
rect 29036 23324 29316 23380
rect 29036 23156 29092 23166
rect 29036 23154 29204 23156
rect 29036 23102 29038 23154
rect 29090 23102 29204 23154
rect 29036 23100 29204 23102
rect 29036 23090 29092 23100
rect 27804 22764 28196 22820
rect 28700 22764 28868 22820
rect 29036 22986 29092 22998
rect 29036 22934 29038 22986
rect 29090 22934 29092 22986
rect 27804 21586 27860 22764
rect 27804 21534 27806 21586
rect 27858 21534 27860 21586
rect 27804 21522 27860 21534
rect 27916 22482 27972 22494
rect 27916 22430 27918 22482
rect 27970 22430 27972 22482
rect 27692 21308 27860 21364
rect 27468 20962 27524 20972
rect 27076 20580 27132 20590
rect 27076 20486 27132 20524
rect 27020 19236 27076 19246
rect 26908 19234 27076 19236
rect 26908 19182 27022 19234
rect 27074 19182 27076 19234
rect 26908 19180 27076 19182
rect 27020 19170 27076 19180
rect 27244 19234 27300 19246
rect 27244 19182 27246 19234
rect 27298 19182 27300 19234
rect 26684 19014 26686 19066
rect 26738 19014 26740 19066
rect 26684 19002 26740 19014
rect 26684 18450 26740 18462
rect 26684 18398 26686 18450
rect 26738 18398 26740 18450
rect 26684 17892 26740 18398
rect 26908 18450 26964 18462
rect 26908 18398 26910 18450
rect 26962 18398 26964 18450
rect 26908 18340 26964 18398
rect 26908 18274 26964 18284
rect 27244 18238 27300 19182
rect 27524 19124 27580 19134
rect 27524 19122 27636 19124
rect 27524 19070 27526 19122
rect 27578 19070 27636 19122
rect 27524 19058 27636 19070
rect 27188 18226 27300 18238
rect 27188 18174 27190 18226
rect 27242 18174 27300 18226
rect 27188 18172 27300 18174
rect 26684 17826 26740 17836
rect 27076 17892 27132 17902
rect 26572 17714 26628 17724
rect 27076 17722 27132 17836
rect 26460 17586 26462 17638
rect 26514 17586 26516 17638
rect 26460 17574 26516 17586
rect 26684 17666 26740 17678
rect 26684 17614 26686 17666
rect 26738 17614 26740 17666
rect 27076 17670 27078 17722
rect 27130 17670 27132 17722
rect 27188 17780 27244 18172
rect 27188 17714 27244 17724
rect 27076 17658 27132 17670
rect 26684 17556 26740 17614
rect 26348 17276 26516 17332
rect 26292 16884 26348 16894
rect 26292 16790 26348 16828
rect 26348 15540 26404 15550
rect 26460 15540 26516 17276
rect 26684 17220 26740 17500
rect 26908 17556 26964 17566
rect 26908 17554 27524 17556
rect 26908 17502 26910 17554
rect 26962 17502 27524 17554
rect 26908 17500 27524 17502
rect 26908 17490 26964 17500
rect 27468 17442 27524 17500
rect 27468 17390 27470 17442
rect 27522 17390 27524 17442
rect 27468 17378 27524 17390
rect 26684 17154 26740 17164
rect 27412 16436 27468 16446
rect 27412 16212 27468 16380
rect 26348 15538 26516 15540
rect 26348 15486 26350 15538
rect 26402 15486 26516 15538
rect 26348 15484 26516 15486
rect 27132 16210 27468 16212
rect 27132 16158 27414 16210
rect 27466 16158 27468 16210
rect 27132 16156 27468 16158
rect 26348 15474 26404 15484
rect 27132 15204 27188 16156
rect 27412 16146 27468 16156
rect 27580 15652 27636 19058
rect 27692 18340 27748 18350
rect 27692 18246 27748 18284
rect 27804 18116 27860 21308
rect 27916 18228 27972 22430
rect 28140 22370 28196 22382
rect 28140 22318 28142 22370
rect 28194 22318 28196 22370
rect 28140 21924 28196 22318
rect 28140 21868 28532 21924
rect 28084 21476 28140 21486
rect 28084 21382 28140 21420
rect 28476 21418 28532 21868
rect 28700 21700 28756 22764
rect 29036 22484 29092 22934
rect 29148 22932 29204 23100
rect 29260 23154 29316 23324
rect 29260 23102 29262 23154
rect 29314 23102 29316 23154
rect 29820 23198 29876 23996
rect 29820 23146 29822 23198
rect 29874 23146 29876 23198
rect 29820 23134 29876 23146
rect 29260 23090 29316 23102
rect 29708 23042 29764 23054
rect 29708 22990 29710 23042
rect 29762 22990 29764 23042
rect 29708 22932 29764 22990
rect 29148 22876 29764 22932
rect 28700 21634 28756 21644
rect 28812 22428 29092 22484
rect 29148 22708 29204 22718
rect 29148 22538 29204 22652
rect 29148 22486 29150 22538
rect 29202 22486 29204 22538
rect 29148 22474 29204 22486
rect 28588 21588 28644 21598
rect 28588 21494 28644 21532
rect 28476 21366 28478 21418
rect 28530 21366 28532 21418
rect 28476 21354 28532 21366
rect 28812 20244 28868 22428
rect 29260 22372 29316 22382
rect 29036 22370 29316 22372
rect 29036 22318 29262 22370
rect 29314 22318 29316 22370
rect 29036 22316 29316 22318
rect 28924 21700 28980 21710
rect 28924 21586 28980 21644
rect 28924 21534 28926 21586
rect 28978 21534 28980 21586
rect 28924 21522 28980 21534
rect 29036 21588 29092 22316
rect 29260 22306 29316 22316
rect 29484 22370 29540 22876
rect 29484 22318 29486 22370
rect 29538 22318 29540 22370
rect 29484 22306 29540 22318
rect 30044 22260 30100 26852
rect 30324 26404 30380 26414
rect 30324 26310 30380 26348
rect 30492 26068 30548 26852
rect 30604 26740 30660 26750
rect 30604 26290 30660 26684
rect 30604 26238 30606 26290
rect 30658 26238 30660 26290
rect 30604 26226 30660 26238
rect 30716 26290 30772 26302
rect 30716 26238 30718 26290
rect 30770 26238 30772 26290
rect 30492 26012 30660 26068
rect 30492 25506 30548 25518
rect 30268 25450 30324 25462
rect 30268 25398 30270 25450
rect 30322 25398 30324 25450
rect 30268 25284 30324 25398
rect 30492 25454 30494 25506
rect 30546 25454 30548 25506
rect 30380 25284 30436 25294
rect 30268 25228 30380 25284
rect 30156 24836 30212 24846
rect 30156 24742 30212 24780
rect 30268 24724 30324 24734
rect 30380 24724 30436 25228
rect 30492 24948 30548 25454
rect 30604 25338 30660 26012
rect 30604 25286 30606 25338
rect 30658 25286 30660 25338
rect 30604 25274 30660 25286
rect 30716 25172 30772 26238
rect 30828 26068 30884 26852
rect 30940 26404 30996 27692
rect 31164 27300 31220 27310
rect 30940 26338 30996 26348
rect 31052 26964 31108 26974
rect 31052 26290 31108 26908
rect 31052 26238 31054 26290
rect 31106 26238 31108 26290
rect 31052 26226 31108 26238
rect 31164 26178 31220 27244
rect 31276 27188 31332 27198
rect 31276 27074 31332 27132
rect 31276 27022 31278 27074
rect 31330 27022 31332 27074
rect 31276 27010 31332 27022
rect 31276 26852 31332 26862
rect 31276 26404 31332 26796
rect 31388 26516 31444 27804
rect 31500 27794 31556 27804
rect 31668 27860 31724 27870
rect 31668 27766 31724 27804
rect 31612 27186 31668 27198
rect 31612 27134 31614 27186
rect 31666 27134 31668 27186
rect 31500 27076 31556 27086
rect 31500 27018 31556 27020
rect 31500 26966 31502 27018
rect 31554 26966 31556 27018
rect 31500 26852 31556 26966
rect 31500 26786 31556 26796
rect 31612 26740 31668 27134
rect 31612 26674 31668 26684
rect 31388 26460 31556 26516
rect 31276 26348 31444 26404
rect 31164 26126 31166 26178
rect 31218 26126 31220 26178
rect 31164 26114 31220 26126
rect 31388 26317 31444 26348
rect 31388 26265 31390 26317
rect 31442 26265 31444 26317
rect 30828 26012 31108 26068
rect 30828 25172 30884 25182
rect 30716 25116 30828 25172
rect 30492 24892 30660 24948
rect 30492 24724 30548 24734
rect 30380 24722 30548 24724
rect 30380 24670 30494 24722
rect 30546 24670 30548 24722
rect 30380 24668 30548 24670
rect 30268 24062 30324 24668
rect 30492 24658 30548 24668
rect 30604 24276 30660 24892
rect 30828 24946 30884 25116
rect 30828 24894 30830 24946
rect 30882 24894 30884 24946
rect 30828 24882 30884 24894
rect 30604 24220 30884 24276
rect 30828 24106 30884 24220
rect 30268 24050 30380 24062
rect 30268 23998 30326 24050
rect 30378 23998 30380 24050
rect 30268 23996 30380 23998
rect 30324 23986 30380 23996
rect 30716 24052 30772 24062
rect 30716 23938 30772 23996
rect 30716 23886 30718 23938
rect 30770 23886 30772 23938
rect 30716 23874 30772 23886
rect 30828 24054 30830 24106
rect 30882 24054 30884 24106
rect 30380 23380 30436 23390
rect 30156 23268 30212 23278
rect 30156 23154 30212 23212
rect 30156 23102 30158 23154
rect 30210 23102 30212 23154
rect 30156 23090 30212 23102
rect 30044 22194 30100 22204
rect 30156 22146 30212 22158
rect 30156 22094 30158 22146
rect 30210 22094 30212 22146
rect 29184 21980 29448 21990
rect 29240 21924 29288 21980
rect 29344 21924 29392 21980
rect 29184 21914 29448 21924
rect 29036 21522 29092 21532
rect 30156 21588 30212 22094
rect 30380 21642 30436 23324
rect 30492 23268 30548 23278
rect 30492 23154 30548 23212
rect 30492 23102 30494 23154
rect 30546 23102 30548 23154
rect 30492 23090 30548 23102
rect 30828 22820 30884 24054
rect 30940 23940 30996 23950
rect 30940 23846 30996 23884
rect 31052 23716 31108 26012
rect 30712 22764 30884 22820
rect 30940 23660 31108 23716
rect 31164 25956 31220 25966
rect 30492 22372 30548 22382
rect 30492 22278 30548 22316
rect 30712 22332 30768 22764
rect 30940 22708 30996 23660
rect 30712 22280 30714 22332
rect 30766 22280 30768 22332
rect 30712 22268 30768 22280
rect 30828 22652 30996 22708
rect 31052 23156 31108 23166
rect 30716 22148 30772 22158
rect 30380 21590 30382 21642
rect 30434 21590 30436 21642
rect 30380 21578 30436 21590
rect 30492 22036 30548 22046
rect 30156 21494 30212 21532
rect 30492 21028 30548 21980
rect 30716 21586 30772 22092
rect 30716 21534 30718 21586
rect 30770 21534 30772 21586
rect 30716 21522 30772 21534
rect 30604 21474 30660 21486
rect 30604 21422 30606 21474
rect 30658 21422 30660 21474
rect 30604 21252 30660 21422
rect 30604 21186 30660 21196
rect 30492 20972 30772 21028
rect 30324 20804 30380 20814
rect 30044 20802 30380 20804
rect 30044 20750 30326 20802
rect 30378 20750 30380 20802
rect 30044 20748 30380 20750
rect 29184 20412 29448 20422
rect 29240 20356 29288 20412
rect 29344 20356 29392 20412
rect 29184 20346 29448 20356
rect 28812 20178 28868 20188
rect 29036 20020 29092 20030
rect 29036 19926 29092 19964
rect 29260 20018 29316 20030
rect 29260 19966 29262 20018
rect 29314 19966 29316 20018
rect 29260 19572 29316 19966
rect 29540 20020 29596 20030
rect 29540 19926 29596 19964
rect 29932 20018 29988 20030
rect 29932 19966 29934 20018
rect 29986 19966 29988 20018
rect 29932 19908 29988 19966
rect 29932 19842 29988 19852
rect 29260 19506 29316 19516
rect 29484 19796 29540 19806
rect 29484 19460 29540 19740
rect 29820 19796 29876 19806
rect 29820 19572 29876 19740
rect 29484 19458 29652 19460
rect 29484 19406 29486 19458
rect 29538 19406 29652 19458
rect 29484 19404 29652 19406
rect 29484 19394 29540 19404
rect 29148 19236 29204 19246
rect 29036 19180 29148 19236
rect 29036 18900 29092 19180
rect 29148 19142 29204 19180
rect 29036 18834 29092 18844
rect 29184 18844 29448 18854
rect 29240 18788 29288 18844
rect 29344 18788 29392 18844
rect 29184 18778 29448 18788
rect 29596 18676 29652 19404
rect 29820 19236 29876 19516
rect 30044 19470 30100 20748
rect 30324 20738 30380 20748
rect 30268 20132 30324 20142
rect 29988 19458 30100 19470
rect 29988 19406 29990 19458
rect 30042 19406 30100 19458
rect 29988 19404 30100 19406
rect 30156 20076 30268 20132
rect 30156 19460 30212 20076
rect 30268 20074 30324 20076
rect 30268 20022 30270 20074
rect 30322 20022 30324 20074
rect 30268 20010 30324 20022
rect 30604 20018 30660 20030
rect 30604 19966 30606 20018
rect 30658 19966 30660 20018
rect 30268 19906 30324 19918
rect 30268 19854 30270 19906
rect 30322 19854 30324 19906
rect 30268 19572 30324 19854
rect 30604 19796 30660 19966
rect 30604 19730 30660 19740
rect 30492 19572 30548 19582
rect 30268 19516 30492 19572
rect 30492 19506 30548 19516
rect 30156 19404 30436 19460
rect 29988 19394 30044 19404
rect 30268 19236 30324 19246
rect 29820 19234 30324 19236
rect 29820 19182 30270 19234
rect 30322 19182 30324 19234
rect 29820 19180 30324 19182
rect 30268 18788 30324 19180
rect 30380 19234 30436 19404
rect 30380 19182 30382 19234
rect 30434 19182 30436 19234
rect 30380 19170 30436 19182
rect 30548 19236 30604 19246
rect 30548 19142 30604 19180
rect 30716 19234 30772 20972
rect 30716 19182 30718 19234
rect 30770 19182 30772 19234
rect 30716 19170 30772 19182
rect 30828 19068 30884 22652
rect 31052 22148 31108 23100
rect 31052 22082 31108 22092
rect 31164 21476 31220 25900
rect 31276 25506 31332 25518
rect 31276 25454 31278 25506
rect 31330 25454 31332 25506
rect 31276 25284 31332 25454
rect 31276 25218 31332 25228
rect 31388 24948 31444 26265
rect 31500 26068 31556 26460
rect 31724 26290 31780 26302
rect 31724 26238 31726 26290
rect 31778 26238 31780 26290
rect 31724 26180 31780 26238
rect 31724 26114 31780 26124
rect 31500 26002 31556 26012
rect 31836 25956 31892 30044
rect 32060 29988 32116 32732
rect 32172 32562 32228 32574
rect 32172 32510 32174 32562
rect 32226 32510 32228 32562
rect 32172 31220 32228 32510
rect 32284 32340 32340 32350
rect 32452 32340 32508 32350
rect 32284 31750 32340 32284
rect 32284 31698 32286 31750
rect 32338 31698 32340 31750
rect 32284 31686 32340 31698
rect 32396 32338 32508 32340
rect 32396 32286 32454 32338
rect 32506 32286 32508 32338
rect 32396 32274 32508 32286
rect 32172 31154 32228 31164
rect 32284 31108 32340 31118
rect 32396 31108 32452 32274
rect 32340 31052 32452 31108
rect 32284 31042 32340 31052
rect 32620 30324 32676 34300
rect 32956 34130 33012 34142
rect 32956 34078 32958 34130
rect 33010 34078 33012 34130
rect 32732 34020 32788 34030
rect 32732 31892 32788 33964
rect 32956 33684 33012 34078
rect 33404 33684 33460 39200
rect 33846 36876 34110 36886
rect 33902 36820 33950 36876
rect 34006 36820 34054 36876
rect 33846 36810 34110 36820
rect 34412 35474 34468 35486
rect 34412 35422 34414 35474
rect 34466 35422 34468 35474
rect 33846 35308 34110 35318
rect 33902 35252 33950 35308
rect 34006 35252 34054 35308
rect 33846 35242 34110 35252
rect 34412 35140 34468 35422
rect 34412 35074 34468 35084
rect 33740 34916 33796 34926
rect 33740 34804 33796 34860
rect 33628 34802 33796 34804
rect 33628 34750 33742 34802
rect 33794 34750 33796 34802
rect 33628 34748 33796 34750
rect 33628 33908 33684 34748
rect 33740 34738 33796 34748
rect 34300 34692 34356 34702
rect 33852 34690 34356 34692
rect 33852 34638 34302 34690
rect 34354 34638 34356 34690
rect 33852 34636 34356 34638
rect 33740 34132 33796 34142
rect 33852 34132 33908 34636
rect 34300 34626 34356 34636
rect 33740 34130 33908 34132
rect 33740 34078 33742 34130
rect 33794 34078 33908 34130
rect 33740 34076 33908 34078
rect 33964 34468 34020 34478
rect 33740 34066 33796 34076
rect 33628 33842 33684 33852
rect 33964 33908 34020 34412
rect 34524 34356 34580 39200
rect 35420 36484 35476 36494
rect 35420 36482 35588 36484
rect 35420 36430 35422 36482
rect 35474 36430 35588 36482
rect 35420 36428 35588 36430
rect 35420 36418 35476 36428
rect 35084 36260 35140 36270
rect 35084 36166 35140 36204
rect 35532 35028 35588 36428
rect 35532 34962 35588 34972
rect 34636 34916 34692 34926
rect 34636 34914 34804 34916
rect 34636 34862 34638 34914
rect 34690 34862 34804 34914
rect 34636 34860 34804 34862
rect 34636 34850 34692 34860
rect 34748 34468 34804 34860
rect 35308 34914 35364 34926
rect 35308 34862 35310 34914
rect 35362 34862 35364 34914
rect 35308 34804 35364 34862
rect 35420 34916 35476 34926
rect 35420 34822 35476 34860
rect 35308 34738 35364 34748
rect 34972 34692 35028 34702
rect 34972 34690 35252 34692
rect 34972 34638 34974 34690
rect 35026 34638 35252 34690
rect 34972 34636 35252 34638
rect 34972 34626 35028 34636
rect 34748 34412 35028 34468
rect 34524 34300 34916 34356
rect 33964 33842 34020 33852
rect 34188 33796 34244 33806
rect 34860 33796 34916 34300
rect 33846 33740 34110 33750
rect 33902 33684 33950 33740
rect 34006 33684 34054 33740
rect 33404 33628 33684 33684
rect 33846 33674 34110 33684
rect 32956 33618 33012 33628
rect 33404 33124 33460 33134
rect 33628 33124 33684 33628
rect 33404 32452 33460 33068
rect 33404 32386 33460 32396
rect 33516 33068 33684 33124
rect 32732 31836 33012 31892
rect 32620 30258 32676 30268
rect 32844 31750 32900 31762
rect 32844 31698 32846 31750
rect 32898 31698 32900 31750
rect 32396 30182 32452 30194
rect 32396 30130 32398 30182
rect 32450 30130 32452 30182
rect 32396 30100 32452 30130
rect 32396 30034 32452 30044
rect 32060 29922 32116 29932
rect 32508 29764 32564 29774
rect 32060 29652 32116 29662
rect 32060 29538 32116 29596
rect 32060 29486 32062 29538
rect 32114 29486 32116 29538
rect 32060 28980 32116 29486
rect 32060 28914 32116 28924
rect 32060 28644 32116 28654
rect 32060 28550 32116 28588
rect 32302 28532 32358 28542
rect 32302 28438 32358 28476
rect 32172 28420 32228 28430
rect 32172 27858 32228 28364
rect 32508 28084 32564 29708
rect 32844 29092 32900 31698
rect 32844 29026 32900 29036
rect 32844 28868 32900 28878
rect 32172 27806 32174 27858
rect 32226 27806 32228 27858
rect 32172 27794 32228 27806
rect 32396 28028 32564 28084
rect 32732 28756 32788 28766
rect 32396 27870 32452 28028
rect 32396 27858 32470 27870
rect 32396 27806 32416 27858
rect 32468 27806 32470 27858
rect 32396 27804 32470 27806
rect 32414 27794 32470 27804
rect 32732 27310 32788 28700
rect 32844 28642 32900 28812
rect 32844 28590 32846 28642
rect 32898 28590 32900 28642
rect 32844 28578 32900 28590
rect 32956 28420 33012 31836
rect 33162 31220 33218 31230
rect 33162 31106 33218 31164
rect 33162 31054 33164 31106
rect 33216 31054 33218 31106
rect 33162 31042 33218 31054
rect 33404 30996 33460 31006
rect 33404 30902 33460 30940
rect 33404 30772 33460 30782
rect 33236 30100 33292 30110
rect 33404 30100 33460 30716
rect 33516 30212 33572 33068
rect 34076 32452 34132 32462
rect 34076 32358 34132 32396
rect 33846 32172 34110 32182
rect 33902 32116 33950 32172
rect 34006 32116 34054 32172
rect 33846 32106 34110 32116
rect 34188 31890 34244 33740
rect 34636 33740 34916 33796
rect 34412 33236 34468 33246
rect 34412 32676 34468 33180
rect 34412 32610 34468 32620
rect 34188 31838 34190 31890
rect 34242 31838 34244 31890
rect 34188 31826 34244 31838
rect 34300 32564 34356 32574
rect 34300 32004 34356 32508
rect 34076 30996 34132 31006
rect 34076 30994 34244 30996
rect 33908 30938 33964 30950
rect 33908 30886 33910 30938
rect 33962 30886 33964 30938
rect 34076 30942 34078 30994
rect 34130 30942 34244 30994
rect 34076 30940 34244 30942
rect 34076 30930 34132 30940
rect 33908 30884 33964 30886
rect 33908 30818 33964 30828
rect 33846 30604 34110 30614
rect 33902 30548 33950 30604
rect 34006 30548 34054 30604
rect 33846 30538 34110 30548
rect 34188 30212 34244 30940
rect 33516 30156 33908 30212
rect 33404 30044 33572 30100
rect 33236 29650 33292 30044
rect 33236 29598 33238 29650
rect 33290 29598 33292 29650
rect 33236 29586 33292 29598
rect 33068 28644 33124 28654
rect 33068 28550 33124 28588
rect 33348 28532 33404 28542
rect 32396 27300 32452 27310
rect 31948 27074 32004 27086
rect 31948 27022 31950 27074
rect 32002 27022 32004 27074
rect 31948 26964 32004 27022
rect 32284 27074 32340 27086
rect 32284 27022 32286 27074
rect 32338 27022 32340 27074
rect 32060 26964 32116 26974
rect 31948 26908 32060 26964
rect 31836 25890 31892 25900
rect 31836 25732 31892 25742
rect 31500 25450 31556 25462
rect 31500 25398 31502 25450
rect 31554 25398 31556 25450
rect 31500 25396 31556 25398
rect 31500 25330 31556 25340
rect 31836 25338 31892 25676
rect 31948 25508 32004 25518
rect 32060 25508 32116 26908
rect 31948 25506 32116 25508
rect 31948 25454 31950 25506
rect 32002 25454 32116 25506
rect 31948 25452 32116 25454
rect 31948 25442 32004 25452
rect 31388 24882 31444 24892
rect 31724 25284 31780 25294
rect 31836 25286 31838 25338
rect 31890 25286 31892 25338
rect 31836 25274 31892 25286
rect 31724 24836 31780 25228
rect 31612 24780 31780 24836
rect 32060 24948 32116 25452
rect 32284 25284 32340 27022
rect 32396 27074 32452 27244
rect 32676 27298 32788 27310
rect 32676 27246 32678 27298
rect 32730 27246 32788 27298
rect 32676 27244 32788 27246
rect 32844 28364 33012 28420
rect 33236 28530 33404 28532
rect 33236 28478 33350 28530
rect 33402 28478 33404 28530
rect 33236 28476 33404 28478
rect 32676 27234 32732 27244
rect 32396 27022 32398 27074
rect 32450 27022 32452 27074
rect 32396 27010 32452 27022
rect 32508 27188 32564 27198
rect 32284 25218 32340 25228
rect 32396 26180 32452 26190
rect 32172 24948 32228 24958
rect 32060 24946 32228 24948
rect 32060 24894 32174 24946
rect 32226 24894 32228 24946
rect 32060 24892 32228 24894
rect 31612 24766 31668 24780
rect 31388 24724 31444 24734
rect 31612 24714 31614 24766
rect 31666 24714 31668 24766
rect 31612 24702 31668 24714
rect 32060 24724 32116 24892
rect 32172 24882 32228 24892
rect 31388 24630 31444 24668
rect 32060 24658 32116 24668
rect 31724 24612 31780 24622
rect 31724 24518 31780 24556
rect 31724 24388 31780 24398
rect 31500 23716 31556 23726
rect 31500 23714 31668 23716
rect 31500 23662 31502 23714
rect 31554 23662 31668 23714
rect 31500 23660 31668 23662
rect 31500 23650 31556 23660
rect 31388 23380 31444 23390
rect 31276 22986 31332 22998
rect 31276 22934 31278 22986
rect 31330 22934 31332 22986
rect 31276 22932 31332 22934
rect 31276 22866 31332 22876
rect 31388 22372 31444 23324
rect 31612 23156 31668 23660
rect 31612 23062 31668 23100
rect 31388 22278 31444 22316
rect 31500 22538 31556 22550
rect 31500 22486 31502 22538
rect 31554 22486 31556 22538
rect 31164 21410 31220 21420
rect 31332 21588 31388 21598
rect 31332 21474 31388 21532
rect 31332 21422 31334 21474
rect 31386 21422 31388 21474
rect 31164 21252 31220 21262
rect 31164 20804 31220 21196
rect 31332 21028 31388 21422
rect 31332 20962 31388 20972
rect 31388 20804 31444 20814
rect 31164 20802 31444 20804
rect 31164 20750 31390 20802
rect 31442 20750 31444 20802
rect 31164 20748 31444 20750
rect 31388 20738 31444 20748
rect 30940 20356 30996 20366
rect 30940 20018 30996 20300
rect 30940 19966 30942 20018
rect 30994 19966 30996 20018
rect 30940 19954 30996 19966
rect 31052 20244 31108 20254
rect 31052 19290 31108 20188
rect 31276 20020 31332 20030
rect 31052 19238 31054 19290
rect 31106 19238 31108 19290
rect 31052 19236 31108 19238
rect 31052 19160 31108 19180
rect 31164 19572 31220 19582
rect 31164 19196 31220 19516
rect 31164 19144 31166 19196
rect 31218 19144 31220 19196
rect 31164 19132 31220 19144
rect 30268 18722 30324 18732
rect 30604 19012 30884 19068
rect 31276 19012 31332 19964
rect 31388 20018 31444 20030
rect 31388 19966 31390 20018
rect 31442 19966 31444 20018
rect 31388 19908 31444 19966
rect 31388 19842 31444 19852
rect 31500 19460 31556 22486
rect 31612 21588 31668 21598
rect 31612 21494 31668 21532
rect 31724 20916 31780 24332
rect 32284 24164 32340 24174
rect 32396 24164 32452 26124
rect 32508 25508 32564 27132
rect 32508 25506 32676 25508
rect 32508 25454 32510 25506
rect 32562 25454 32676 25506
rect 32508 25452 32676 25454
rect 32508 25442 32564 25452
rect 32508 25060 32564 25070
rect 32508 24722 32564 25004
rect 32508 24670 32510 24722
rect 32562 24670 32564 24722
rect 32508 24658 32564 24670
rect 32620 24388 32676 25452
rect 32732 25450 32788 25462
rect 32732 25398 32734 25450
rect 32786 25398 32788 25450
rect 32732 24612 32788 25398
rect 32844 25060 32900 28364
rect 33236 27914 33292 28476
rect 33348 28466 33404 28476
rect 33516 28308 33572 30044
rect 33852 29426 33908 30156
rect 33852 29374 33854 29426
rect 33906 29374 33908 29426
rect 33852 29362 33908 29374
rect 34076 30156 34244 30212
rect 34300 30994 34356 31948
rect 34300 30942 34302 30994
rect 34354 30942 34356 30994
rect 34076 29204 34132 30156
rect 34188 29988 34244 29998
rect 34188 29894 34244 29932
rect 34076 29148 34244 29204
rect 33846 29036 34110 29046
rect 33902 28980 33950 29036
rect 34006 28980 34054 29036
rect 33846 28970 34110 28980
rect 33068 27860 33124 27870
rect 32956 27858 33124 27860
rect 32956 27806 33070 27858
rect 33122 27806 33124 27858
rect 33236 27862 33238 27914
rect 33290 27862 33292 27914
rect 33236 27850 33292 27862
rect 33404 28252 33572 28308
rect 33740 28532 33796 28542
rect 32956 27804 33124 27806
rect 32956 25618 33012 27804
rect 33068 27794 33124 27804
rect 33404 27046 33460 28252
rect 33740 27860 33796 28476
rect 34188 27972 34244 29148
rect 34188 27906 34244 27916
rect 34300 27860 34356 30942
rect 34412 30884 34468 30894
rect 34412 29988 34468 30828
rect 34412 29204 34468 29932
rect 34412 29138 34468 29148
rect 34636 28868 34692 33740
rect 34972 33460 35028 34412
rect 34748 33404 35028 33460
rect 35084 34244 35140 34254
rect 35084 33460 35140 34188
rect 34748 30100 34804 33404
rect 35084 33394 35140 33404
rect 35028 33290 35084 33302
rect 34748 30034 34804 30044
rect 34860 33234 34916 33246
rect 34860 33182 34862 33234
rect 34914 33182 34916 33234
rect 34860 29204 34916 33182
rect 35028 33238 35030 33290
rect 35082 33238 35084 33290
rect 35028 33236 35084 33238
rect 35028 33170 35084 33180
rect 35196 32788 35252 34636
rect 35644 34468 35700 39200
rect 36148 36372 36204 36382
rect 36148 36278 36204 36316
rect 35980 36260 36036 36270
rect 35756 35700 35812 35710
rect 35756 35698 35924 35700
rect 35756 35646 35758 35698
rect 35810 35646 35924 35698
rect 35756 35644 35924 35646
rect 35756 35634 35812 35644
rect 35644 34402 35700 34412
rect 35756 34690 35812 34702
rect 35756 34638 35758 34690
rect 35810 34638 35812 34690
rect 35644 34018 35700 34030
rect 35644 33966 35646 34018
rect 35698 33966 35700 34018
rect 35420 33908 35476 33918
rect 35420 33460 35476 33852
rect 35644 33908 35700 33966
rect 35644 33842 35700 33852
rect 35756 33460 35812 34638
rect 35420 33404 35588 33460
rect 35532 33402 35588 33404
rect 35532 33350 35534 33402
rect 35586 33350 35588 33402
rect 35532 33338 35588 33350
rect 35644 33404 35812 33460
rect 35868 33460 35924 35644
rect 35084 32732 35252 32788
rect 35420 32900 35476 32910
rect 35084 31668 35140 32732
rect 35196 32562 35252 32574
rect 35196 32510 35198 32562
rect 35250 32510 35252 32562
rect 35196 31892 35252 32510
rect 35308 32564 35364 32574
rect 35308 32470 35364 32508
rect 35196 31826 35252 31836
rect 35084 31612 35252 31668
rect 35084 30884 35140 30894
rect 35084 30790 35140 30828
rect 35196 30212 35252 31612
rect 35420 31220 35476 32844
rect 35644 32340 35700 33404
rect 35868 33394 35924 33404
rect 35774 33236 35830 33246
rect 35644 32274 35700 32284
rect 35756 33234 35830 33236
rect 35756 33182 35776 33234
rect 35828 33182 35830 33234
rect 35756 33170 35830 33182
rect 35308 31164 35476 31220
rect 35756 31220 35812 33170
rect 35868 33012 35924 33022
rect 35868 32116 35924 32956
rect 35980 32228 36036 36204
rect 36428 35700 36484 35710
rect 36204 35698 36484 35700
rect 36204 35646 36430 35698
rect 36482 35646 36484 35698
rect 36204 35644 36484 35646
rect 36764 35700 36820 39200
rect 38332 37492 38388 37502
rect 37604 37044 37660 37054
rect 37604 36594 37660 36988
rect 37604 36542 37606 36594
rect 37658 36542 37660 36594
rect 37604 36530 37660 36542
rect 38332 37044 38388 37436
rect 38332 36482 38388 36988
rect 38332 36430 38334 36482
rect 38386 36430 38388 36482
rect 38332 36418 38388 36430
rect 37996 36258 38052 36270
rect 37996 36206 37998 36258
rect 38050 36206 38052 36258
rect 36764 35644 36932 35700
rect 36092 35474 36148 35486
rect 36092 35422 36094 35474
rect 36146 35422 36148 35474
rect 36092 32614 36148 35422
rect 36204 34356 36260 35644
rect 36428 35634 36484 35644
rect 36764 35476 36820 35486
rect 36540 35474 36820 35476
rect 36540 35422 36766 35474
rect 36818 35422 36820 35474
rect 36540 35420 36820 35422
rect 36372 34804 36428 34814
rect 36372 34710 36428 34748
rect 36204 34290 36260 34300
rect 36260 34132 36316 34142
rect 36260 34038 36316 34076
rect 36372 33124 36428 33134
rect 36372 33030 36428 33068
rect 36540 32900 36596 35420
rect 36764 35410 36820 35420
rect 36708 34020 36764 34030
rect 36652 34018 36764 34020
rect 36652 33966 36710 34018
rect 36762 33966 36764 34018
rect 36652 33954 36764 33966
rect 36652 33124 36708 33954
rect 36652 33058 36708 33068
rect 36540 32834 36596 32844
rect 36876 32788 36932 35644
rect 37996 35476 38052 36206
rect 38508 36092 38772 36102
rect 38564 36036 38612 36092
rect 38668 36036 38716 36092
rect 38508 36026 38772 36036
rect 37996 35410 38052 35420
rect 37828 34692 37884 34702
rect 37660 34690 37884 34692
rect 37660 34638 37830 34690
rect 37882 34638 37884 34690
rect 37660 34636 37884 34638
rect 37660 34130 37716 34636
rect 37828 34626 37884 34636
rect 38276 34692 38332 34702
rect 38276 34690 38388 34692
rect 38276 34638 38278 34690
rect 38330 34638 38388 34690
rect 38276 34626 38388 34638
rect 37660 34078 37662 34130
rect 37714 34078 37716 34130
rect 37324 34020 37380 34030
rect 37660 34020 37716 34078
rect 37324 33926 37380 33964
rect 37436 33964 37716 34020
rect 38332 34130 38388 34626
rect 38508 34524 38772 34534
rect 38564 34468 38612 34524
rect 38668 34468 38716 34524
rect 38508 34458 38772 34468
rect 38332 34078 38334 34130
rect 38386 34078 38388 34130
rect 37156 33290 37212 33302
rect 36988 33236 37044 33246
rect 36988 33142 37044 33180
rect 37156 33238 37158 33290
rect 37210 33238 37212 33290
rect 37156 32788 37212 33238
rect 37156 32732 37380 32788
rect 36876 32722 36932 32732
rect 36092 32558 36372 32614
rect 36092 32452 36148 32462
rect 36092 32358 36148 32396
rect 35980 32172 36148 32228
rect 35868 32050 35924 32060
rect 35924 31892 35980 31902
rect 35924 31798 35980 31836
rect 36092 31220 36148 32172
rect 36204 32116 36260 32126
rect 36316 32116 36372 32558
rect 36652 32228 36708 32238
rect 36540 32116 36596 32126
rect 36316 32060 36484 32116
rect 36204 32004 36260 32060
rect 36204 31948 36372 32004
rect 36204 31778 36260 31790
rect 36204 31726 36206 31778
rect 36258 31726 36260 31778
rect 36204 31332 36260 31726
rect 36316 31778 36372 31948
rect 36316 31726 36318 31778
rect 36370 31726 36372 31778
rect 36316 31714 36372 31726
rect 36204 31276 36372 31332
rect 36092 31164 36260 31220
rect 35308 30660 35364 31164
rect 35756 31154 35812 31164
rect 35308 30604 35812 30660
rect 35196 30182 35364 30212
rect 35196 30156 35310 30182
rect 35308 30130 35310 30156
rect 35362 30130 35364 30182
rect 35308 30118 35364 30130
rect 34972 29204 35028 29214
rect 34860 29148 34972 29204
rect 34748 28868 34804 28878
rect 34636 28866 34804 28868
rect 34636 28814 34750 28866
rect 34802 28814 34804 28866
rect 34636 28812 34804 28814
rect 34748 28802 34804 28812
rect 34860 28084 34916 28094
rect 34748 27860 34804 27870
rect 33740 27858 34132 27860
rect 33740 27806 33742 27858
rect 33794 27806 34132 27858
rect 33740 27804 34132 27806
rect 34300 27858 34804 27860
rect 34300 27806 34750 27858
rect 34802 27806 34804 27858
rect 34300 27804 34804 27806
rect 33740 27794 33796 27804
rect 34076 27748 34132 27804
rect 34748 27794 34804 27804
rect 34076 27692 34244 27748
rect 33982 27636 34038 27646
rect 33404 26994 33406 27046
rect 33458 26994 33460 27046
rect 33236 26516 33292 26526
rect 33404 26516 33460 26994
rect 33236 26514 33460 26516
rect 33236 26462 33238 26514
rect 33290 26462 33460 26514
rect 33236 26460 33460 26462
rect 33628 27634 34038 27636
rect 33628 27582 33984 27634
rect 34036 27582 34038 27634
rect 33628 27580 34038 27582
rect 33236 26450 33292 26460
rect 33628 26290 33684 27580
rect 33982 27570 34038 27580
rect 33846 27468 34110 27478
rect 33902 27412 33950 27468
rect 34006 27412 34054 27468
rect 33846 27402 34110 27412
rect 34188 26908 34244 27692
rect 34412 27636 34468 27646
rect 34188 26852 34356 26908
rect 33628 26238 33630 26290
rect 33682 26238 33684 26290
rect 33628 26226 33684 26238
rect 32956 25566 32958 25618
rect 33010 25566 33012 25618
rect 32956 25554 33012 25566
rect 33628 26068 33684 26078
rect 33180 25508 33236 25518
rect 33516 25508 33572 25518
rect 33180 25506 33460 25508
rect 33180 25454 33182 25506
rect 33234 25454 33460 25506
rect 33180 25452 33460 25454
rect 33180 25442 33236 25452
rect 33404 25060 33460 25452
rect 33516 25414 33572 25452
rect 33628 25338 33684 26012
rect 33846 25900 34110 25910
rect 33902 25844 33950 25900
rect 34006 25844 34054 25900
rect 33846 25834 34110 25844
rect 34188 25506 34244 25518
rect 33628 25286 33630 25338
rect 33682 25286 33684 25338
rect 33852 25450 33908 25462
rect 33852 25398 33854 25450
rect 33906 25398 33908 25450
rect 33852 25396 33908 25398
rect 33852 25330 33908 25340
rect 34188 25454 34190 25506
rect 34242 25454 34244 25506
rect 33628 25274 33684 25286
rect 34188 25284 34244 25454
rect 34188 25218 34244 25228
rect 32844 25004 33012 25060
rect 33404 25004 33796 25060
rect 32788 24556 32900 24612
rect 32732 24546 32788 24556
rect 32620 24332 32788 24388
rect 32284 24162 32676 24164
rect 32284 24110 32286 24162
rect 32338 24110 32676 24162
rect 32284 24108 32676 24110
rect 32284 24098 32340 24108
rect 31836 23940 31892 23950
rect 31836 23846 31892 23884
rect 31948 23940 32004 23950
rect 31948 23938 32116 23940
rect 31948 23886 31950 23938
rect 32002 23886 32116 23938
rect 31948 23884 32116 23886
rect 31948 23874 32004 23884
rect 31948 23604 32004 23614
rect 31836 22370 31892 22382
rect 31836 22318 31838 22370
rect 31890 22318 31892 22370
rect 31836 22036 31892 22318
rect 31836 21970 31892 21980
rect 31948 21642 32004 23548
rect 31948 21590 31950 21642
rect 32002 21590 32004 21642
rect 31948 21578 32004 21590
rect 32060 22932 32116 23884
rect 31948 21474 32004 21486
rect 31948 21422 31950 21474
rect 32002 21422 32004 21474
rect 31724 20860 31892 20916
rect 31724 20690 31780 20702
rect 31724 20638 31726 20690
rect 31778 20638 31780 20690
rect 31612 20020 31668 20030
rect 31612 19926 31668 19964
rect 29484 18620 29652 18676
rect 29484 18564 29540 18620
rect 29484 18470 29540 18508
rect 30268 18564 30324 18574
rect 28028 18452 28084 18462
rect 28028 18358 28084 18396
rect 29372 18450 29428 18462
rect 29372 18398 29374 18450
rect 29426 18398 29428 18450
rect 29820 18452 29876 18462
rect 29092 18228 29148 18238
rect 27916 18172 28084 18228
rect 27692 18060 27860 18116
rect 27692 16660 27748 18060
rect 27804 17444 27860 17454
rect 27804 17442 27972 17444
rect 27804 17390 27806 17442
rect 27858 17390 27972 17442
rect 27804 17388 27972 17390
rect 27804 17378 27860 17388
rect 27804 17220 27860 17230
rect 27804 16996 27860 17164
rect 27804 16882 27860 16940
rect 27804 16830 27806 16882
rect 27858 16830 27860 16882
rect 27804 16818 27860 16830
rect 27692 16604 27860 16660
rect 27468 15596 27636 15652
rect 27468 15426 27524 15596
rect 27468 15374 27470 15426
rect 27522 15374 27524 15426
rect 27468 15362 27524 15374
rect 27636 15258 27692 15270
rect 27636 15206 27638 15258
rect 27690 15206 27692 15258
rect 27636 15204 27692 15206
rect 27132 15148 27692 15204
rect 26124 15092 26628 15148
rect 25340 14438 25396 14476
rect 25900 14644 25956 14654
rect 25900 14530 25956 14588
rect 25900 14478 25902 14530
rect 25954 14478 25956 14530
rect 25900 14466 25956 14478
rect 26404 14532 26460 14552
rect 26404 14474 26460 14476
rect 24836 14420 24892 14430
rect 24836 14326 24892 14364
rect 25658 14420 25714 14430
rect 25788 14420 25844 14430
rect 25658 14418 25732 14420
rect 25658 14366 25660 14418
rect 25712 14366 25732 14418
rect 25658 14354 25732 14366
rect 25676 13746 25732 14354
rect 25676 13694 25678 13746
rect 25730 13694 25732 13746
rect 25676 13682 25732 13694
rect 25788 13746 25844 14364
rect 26404 14422 26406 14474
rect 26458 14422 26460 14474
rect 26572 14530 26628 15092
rect 27132 14654 27188 15148
rect 27076 14644 27188 14654
rect 27132 14588 27188 14644
rect 27076 14550 27132 14588
rect 26572 14478 26574 14530
rect 26626 14478 26628 14530
rect 26572 14466 26628 14478
rect 26404 14308 26460 14422
rect 25788 13694 25790 13746
rect 25842 13694 25844 13746
rect 25788 13682 25844 13694
rect 26348 14252 26460 14308
rect 24500 13634 24556 13646
rect 24500 13582 24502 13634
rect 24554 13582 24556 13634
rect 24332 13524 24388 13534
rect 24500 13524 24556 13582
rect 25340 13524 25396 13534
rect 26124 13524 26180 13534
rect 24500 13468 24948 13524
rect 24332 13074 24388 13468
rect 24522 13356 24786 13366
rect 24578 13300 24626 13356
rect 24682 13300 24730 13356
rect 24522 13290 24786 13300
rect 24892 13300 24948 13468
rect 25340 13430 25396 13468
rect 25900 13522 26180 13524
rect 25900 13470 26126 13522
rect 26178 13470 26180 13522
rect 25900 13468 26180 13470
rect 24892 13234 24948 13244
rect 24332 13022 24334 13074
rect 24386 13022 24388 13074
rect 24332 13010 24388 13022
rect 24220 12684 24388 12740
rect 23324 12402 23436 12414
rect 23324 12350 23382 12402
rect 23434 12350 23436 12402
rect 23324 12348 23436 12350
rect 23380 12338 23436 12348
rect 23212 11778 23268 11788
rect 23044 11508 23100 11518
rect 22764 11506 23100 11508
rect 22764 11454 23046 11506
rect 23098 11454 23100 11506
rect 22764 11452 23100 11454
rect 22184 11330 22240 11340
rect 22428 9828 22484 9838
rect 22428 9734 22484 9772
rect 21980 9202 22036 9212
rect 22764 9268 22820 11452
rect 23044 11442 23100 11452
rect 23884 10610 23940 10622
rect 23884 10558 23886 10610
rect 23938 10558 23940 10610
rect 23548 10388 23604 10398
rect 23212 10386 23604 10388
rect 23212 10334 23550 10386
rect 23602 10334 23604 10386
rect 23212 10332 23604 10334
rect 23212 9938 23268 10332
rect 23548 10322 23604 10332
rect 23884 10164 23940 10558
rect 23884 10098 23940 10108
rect 23212 9886 23214 9938
rect 23266 9886 23268 9938
rect 23212 9874 23268 9886
rect 22764 9202 22820 9212
rect 24332 8428 24388 12684
rect 25116 12180 25172 12190
rect 25116 12086 25172 12124
rect 25900 12178 25956 13468
rect 26124 13458 26180 13468
rect 26236 13076 26292 13086
rect 26348 13076 26404 14252
rect 27244 14196 27300 14206
rect 27244 13746 27300 14140
rect 27244 13694 27246 13746
rect 27298 13694 27300 13746
rect 27244 13682 27300 13694
rect 26236 13074 26404 13076
rect 26236 13022 26238 13074
rect 26290 13022 26404 13074
rect 26236 13020 26404 13022
rect 27804 13076 27860 16604
rect 27916 16098 27972 17388
rect 27916 16046 27918 16098
rect 27970 16046 27972 16098
rect 27916 16034 27972 16046
rect 28028 15148 28084 18172
rect 28924 18226 29148 18228
rect 28924 18174 29094 18226
rect 29146 18174 29148 18226
rect 28924 18172 29148 18174
rect 28644 17780 28700 17790
rect 28644 17686 28700 17724
rect 28140 17556 28196 17566
rect 28140 17106 28196 17500
rect 28140 17054 28142 17106
rect 28194 17054 28196 17106
rect 28140 17042 28196 17054
rect 28588 16884 28644 16894
rect 28588 16790 28644 16828
rect 28924 16882 28980 18172
rect 29092 18162 29148 18172
rect 29372 18228 29428 18398
rect 29372 18162 29428 18172
rect 29652 18394 29708 18406
rect 29652 18342 29654 18394
rect 29706 18342 29708 18394
rect 29820 18358 29876 18396
rect 30268 18450 30324 18508
rect 30268 18398 30270 18450
rect 30322 18398 30324 18450
rect 30268 18386 30324 18398
rect 29652 17790 29708 18342
rect 30156 18282 30212 18294
rect 30156 18230 30158 18282
rect 30210 18230 30212 18282
rect 30156 17892 30212 18230
rect 29372 17780 29428 17790
rect 29372 17666 29428 17724
rect 29596 17780 29708 17790
rect 29652 17724 29708 17780
rect 29932 17836 30212 17892
rect 30268 18228 30324 18238
rect 29596 17714 29652 17724
rect 29372 17614 29374 17666
rect 29426 17614 29428 17666
rect 29372 17602 29428 17614
rect 29820 17668 29876 17678
rect 29820 17574 29876 17612
rect 29932 17666 29988 17836
rect 29932 17614 29934 17666
rect 29986 17614 29988 17666
rect 29204 17444 29260 17454
rect 29932 17444 29988 17614
rect 29036 17442 29260 17444
rect 29036 17390 29206 17442
rect 29258 17390 29260 17442
rect 29036 17388 29260 17390
rect 29036 17220 29092 17388
rect 29204 17378 29260 17388
rect 29552 17388 29988 17444
rect 30098 17610 30154 17622
rect 30098 17558 30100 17610
rect 30152 17558 30154 17610
rect 30098 17444 30154 17558
rect 29184 17276 29448 17286
rect 29240 17220 29288 17276
rect 29344 17220 29392 17276
rect 29184 17210 29448 17220
rect 29036 17154 29092 17164
rect 29552 16922 29608 17388
rect 30098 17378 30154 17388
rect 30268 17220 30324 18172
rect 30492 17780 30548 17790
rect 30156 17164 30324 17220
rect 30380 17778 30548 17780
rect 30380 17726 30494 17778
rect 30546 17726 30548 17778
rect 30380 17724 30548 17726
rect 28924 16830 28926 16882
rect 28978 16830 28980 16882
rect 28924 16818 28980 16830
rect 29372 16884 29428 16894
rect 29552 16870 29554 16922
rect 29606 16870 29608 16922
rect 29552 16858 29608 16870
rect 29708 16918 29764 16930
rect 29708 16866 29710 16918
rect 29762 16866 29764 16918
rect 29036 16714 29092 16726
rect 29036 16662 29038 16714
rect 29090 16662 29092 16714
rect 28588 16548 28644 16558
rect 28252 16436 28308 16446
rect 28252 16042 28308 16380
rect 28364 16212 28420 16222
rect 28364 16118 28420 16156
rect 28252 15990 28254 16042
rect 28306 15990 28308 16042
rect 28252 15978 28308 15990
rect 28588 16098 28644 16492
rect 28588 16046 28590 16098
rect 28642 16046 28644 16098
rect 28140 15316 28196 15326
rect 28140 15222 28196 15260
rect 28588 15316 28644 16046
rect 29036 16100 29092 16662
rect 29372 16548 29428 16828
rect 29036 16034 29092 16044
rect 29328 16492 29428 16548
rect 29484 16770 29540 16782
rect 29484 16718 29486 16770
rect 29538 16718 29540 16770
rect 29328 16065 29384 16492
rect 29328 16013 29330 16065
rect 29382 16013 29384 16065
rect 29328 16001 29384 16013
rect 29484 16061 29540 16718
rect 29484 16009 29486 16061
rect 29538 16009 29540 16061
rect 29148 15986 29204 15998
rect 29484 15997 29540 16009
rect 29148 15934 29150 15986
rect 29202 15934 29204 15986
rect 29148 15876 29204 15934
rect 29148 15820 29652 15876
rect 29184 15708 29448 15718
rect 29240 15652 29288 15708
rect 29344 15652 29392 15708
rect 29184 15642 29448 15652
rect 28588 15250 28644 15260
rect 28812 15314 28868 15326
rect 28812 15262 28814 15314
rect 28866 15262 28868 15314
rect 26236 13010 26292 13020
rect 27804 12290 27860 13020
rect 27804 12238 27806 12290
rect 27858 12238 27860 12290
rect 27804 12226 27860 12238
rect 27916 15092 28084 15148
rect 25900 12126 25902 12178
rect 25954 12126 25956 12178
rect 25900 12114 25956 12126
rect 24522 11788 24786 11798
rect 24578 11732 24626 11788
rect 24682 11732 24730 11788
rect 24522 11722 24786 11732
rect 25116 11732 25172 11742
rect 25116 10612 25172 11676
rect 26348 11394 26404 11406
rect 26348 11342 26350 11394
rect 26402 11342 26404 11394
rect 26068 11284 26124 11294
rect 26068 11282 26180 11284
rect 26068 11230 26070 11282
rect 26122 11230 26180 11282
rect 26068 11218 26180 11230
rect 25004 10610 25172 10612
rect 25004 10558 25118 10610
rect 25170 10558 25172 10610
rect 25004 10556 25172 10558
rect 24522 10220 24786 10230
rect 24578 10164 24626 10220
rect 24682 10164 24730 10220
rect 24522 10154 24786 10164
rect 24522 8652 24786 8662
rect 24578 8596 24626 8652
rect 24682 8596 24730 8652
rect 24522 8586 24786 8596
rect 19628 7980 20020 8036
rect 18956 7644 19236 7700
rect 17108 7410 17164 7420
rect 17276 7476 17332 7486
rect 17276 7382 17332 7420
rect 18060 7362 18116 7374
rect 18060 7310 18062 7362
rect 18114 7310 18116 7362
rect 17948 6916 18004 6926
rect 18060 6916 18116 7310
rect 17948 6914 18116 6916
rect 17948 6862 17950 6914
rect 18002 6862 18116 6914
rect 17948 6860 18116 6862
rect 17948 6850 18004 6860
rect 19012 6804 19068 6814
rect 19012 6746 19068 6748
rect 18844 6692 18900 6702
rect 18844 6598 18900 6636
rect 19012 6694 19014 6746
rect 19066 6694 19068 6746
rect 18060 6580 18116 6590
rect 16940 6402 16996 6412
rect 17948 6468 18004 6478
rect 16100 6066 16156 6076
rect 16492 6132 16548 6142
rect 16268 5236 16324 5246
rect 16268 5142 16324 5180
rect 15820 4398 15822 4450
rect 15874 4398 15876 4450
rect 15820 4386 15876 4398
rect 15260 4340 15316 4350
rect 15260 4246 15316 4284
rect 15988 4340 16044 4350
rect 15988 4246 16044 4284
rect 16492 4338 16548 6076
rect 17500 6132 17556 6142
rect 17500 5933 17556 6076
rect 17500 5881 17502 5933
rect 17554 5881 17556 5933
rect 17500 5869 17556 5881
rect 17388 5684 17444 5694
rect 17388 4676 17444 5628
rect 17276 4620 17444 4676
rect 16492 4286 16494 4338
rect 16546 4286 16548 4338
rect 16492 4274 16548 4286
rect 16734 4340 16790 4350
rect 16734 4246 16790 4284
rect 15198 3948 15462 3958
rect 15254 3892 15302 3948
rect 15358 3892 15406 3948
rect 15198 3882 15462 3892
rect 14588 3490 14644 3500
rect 13916 3462 13972 3474
rect 15596 3332 15652 3342
rect 15484 3330 15652 3332
rect 15484 3278 15598 3330
rect 15650 3278 15652 3330
rect 15484 3276 15652 3278
rect 15484 800 15540 3276
rect 15596 3266 15652 3276
rect 17276 800 17332 4620
rect 17444 4452 17500 4462
rect 17444 4358 17500 4396
rect 17724 4340 17780 4350
rect 17724 4246 17780 4284
rect 17948 4338 18004 6412
rect 17948 4286 17950 4338
rect 18002 4286 18004 4338
rect 17948 4274 18004 4286
rect 18060 3526 18116 6524
rect 19012 6580 19068 6694
rect 19012 6514 19068 6524
rect 19180 6692 19236 7644
rect 18172 6132 18228 6142
rect 18172 5234 18228 6076
rect 19180 6020 19236 6636
rect 19516 6690 19572 6702
rect 19516 6638 19518 6690
rect 19570 6638 19572 6690
rect 19516 6580 19572 6638
rect 19516 6514 19572 6524
rect 19180 5954 19236 5964
rect 18508 5684 18564 5694
rect 18508 5590 18564 5628
rect 18172 5182 18174 5234
rect 18226 5182 18228 5234
rect 18172 5170 18228 5182
rect 19628 5236 19684 7980
rect 19860 7868 20124 7878
rect 19916 7812 19964 7868
rect 20020 7812 20068 7868
rect 19860 7802 20124 7812
rect 20524 7476 20580 8372
rect 21756 8260 21812 8270
rect 20636 8146 20692 8158
rect 20636 8094 20638 8146
rect 20690 8094 20692 8146
rect 20636 7700 20692 8094
rect 20636 7644 21308 7700
rect 20748 7476 20804 7486
rect 20524 7420 20692 7476
rect 19964 7362 20020 7374
rect 19964 7310 19966 7362
rect 20018 7310 20020 7362
rect 19964 6804 20020 7310
rect 20506 7250 20562 7262
rect 20506 7198 20508 7250
rect 20560 7198 20562 7250
rect 20506 7140 20562 7198
rect 19964 6738 20020 6748
rect 20412 7084 20562 7140
rect 19758 6692 19814 6702
rect 19758 6598 19814 6636
rect 20076 6692 20132 6702
rect 20300 6692 20356 6702
rect 20076 6690 20244 6692
rect 20076 6638 20078 6690
rect 20130 6638 20244 6690
rect 20076 6636 20244 6638
rect 20076 6468 20132 6636
rect 20188 6468 20244 6636
rect 20300 6598 20356 6636
rect 20300 6468 20356 6478
rect 20188 6412 20300 6468
rect 20076 6402 20132 6412
rect 19860 6300 20124 6310
rect 19916 6244 19964 6300
rect 20020 6244 20068 6300
rect 19860 6234 20124 6244
rect 20300 5906 20356 6412
rect 20300 5854 20302 5906
rect 20354 5854 20356 5906
rect 20300 5842 20356 5854
rect 20412 5906 20468 7084
rect 20636 6702 20692 7420
rect 20748 7474 21028 7476
rect 20748 7422 20750 7474
rect 20802 7422 21028 7474
rect 20748 7420 21028 7422
rect 20748 7410 20804 7420
rect 20580 6690 20692 6702
rect 20580 6638 20582 6690
rect 20634 6638 20692 6690
rect 20580 6636 20692 6638
rect 20580 6626 20636 6636
rect 20412 5854 20414 5906
rect 20466 5854 20468 5906
rect 20412 5842 20468 5854
rect 20972 5794 21028 7420
rect 21252 7418 21308 7644
rect 21252 7366 21254 7418
rect 21306 7366 21308 7418
rect 21420 7476 21476 7486
rect 21420 7474 21588 7476
rect 21420 7422 21422 7474
rect 21474 7422 21588 7474
rect 21420 7420 21588 7422
rect 21420 7410 21476 7420
rect 21252 6804 21308 7366
rect 21196 6748 21308 6804
rect 20972 5742 20974 5794
rect 21026 5742 21028 5794
rect 20692 5684 20748 5694
rect 20692 5682 20916 5684
rect 20692 5630 20694 5682
rect 20746 5630 20916 5682
rect 20692 5628 20916 5630
rect 20692 5618 20748 5628
rect 19628 5170 19684 5180
rect 20860 5122 20916 5628
rect 20860 5070 20862 5122
rect 20914 5070 20916 5122
rect 20860 5058 20916 5070
rect 18788 5012 18844 5022
rect 18788 4898 18844 4956
rect 18788 4846 18790 4898
rect 18842 4846 18844 4898
rect 18340 4340 18396 4350
rect 18508 4340 18564 4350
rect 18788 4340 18844 4846
rect 19404 4898 19460 4910
rect 19404 4846 19406 4898
rect 19458 4846 19460 4898
rect 18340 4338 18844 4340
rect 18340 4286 18342 4338
rect 18394 4286 18510 4338
rect 18562 4286 18844 4338
rect 18340 4284 18844 4286
rect 19292 4340 19348 4350
rect 19404 4340 19460 4846
rect 19860 4732 20124 4742
rect 19916 4676 19964 4732
rect 20020 4676 20068 4732
rect 19860 4666 20124 4676
rect 19292 4338 19460 4340
rect 19292 4286 19294 4338
rect 19346 4286 19460 4338
rect 19292 4284 19460 4286
rect 18340 4274 18396 4284
rect 18508 4274 18564 4284
rect 19292 4274 19348 4284
rect 20972 3780 21028 5742
rect 20972 3714 21028 3724
rect 21084 6580 21140 6590
rect 21196 6580 21252 6748
rect 21140 6524 21252 6580
rect 18060 3474 18062 3526
rect 18114 3474 18116 3526
rect 18060 3462 18116 3474
rect 20860 3668 20916 3678
rect 19068 3330 19124 3342
rect 19068 3278 19070 3330
rect 19122 3278 19124 3330
rect 19068 800 19124 3278
rect 19860 3164 20124 3174
rect 19916 3108 19964 3164
rect 20020 3108 20068 3164
rect 19860 3098 20124 3108
rect 20860 800 20916 3612
rect 21084 3526 21140 6524
rect 21420 6468 21476 6478
rect 21420 6374 21476 6412
rect 21532 6244 21588 7420
rect 21756 6690 21812 8204
rect 21868 7474 21924 8428
rect 24220 8372 24388 8428
rect 24892 8484 24948 8494
rect 25004 8484 25060 10556
rect 25116 10546 25172 10556
rect 25900 11172 25956 11182
rect 25900 10610 25956 11116
rect 25900 10558 25902 10610
rect 25954 10558 25956 10610
rect 25900 10546 25956 10558
rect 26012 10836 26068 10846
rect 26012 10164 26068 10780
rect 26124 10276 26180 11218
rect 26348 10836 26404 11342
rect 26572 11394 26628 11406
rect 26572 11342 26574 11394
rect 26626 11342 26628 11394
rect 26572 10836 26628 11342
rect 27244 11396 27300 11406
rect 27244 11394 27524 11396
rect 27244 11342 27246 11394
rect 27298 11342 27524 11394
rect 27244 11340 27524 11342
rect 27244 11330 27300 11340
rect 26908 11172 26964 11182
rect 26908 11078 26964 11116
rect 26572 10780 27076 10836
rect 26348 10770 26404 10780
rect 26124 10220 26684 10276
rect 25676 10052 25732 10062
rect 26012 10052 26068 10108
rect 26012 9996 26516 10052
rect 25116 9828 25172 9838
rect 25116 9734 25172 9772
rect 24948 8428 25060 8484
rect 25676 8428 25732 9996
rect 26124 9828 26180 9838
rect 26180 9772 26292 9828
rect 26124 9734 26180 9772
rect 25882 9716 25938 9726
rect 25882 9714 26068 9716
rect 25882 9662 25884 9714
rect 25936 9662 26068 9714
rect 25882 9660 26068 9662
rect 25882 9650 25938 9660
rect 26012 9044 26068 9660
rect 26012 8988 26180 9044
rect 25994 8820 26050 8830
rect 26124 8820 26180 8988
rect 26236 9042 26292 9772
rect 26460 9716 26516 9996
rect 26628 9882 26684 10220
rect 27020 10052 27076 10780
rect 26628 9830 26630 9882
rect 26682 9830 26684 9882
rect 26628 9818 26684 9830
rect 26908 9996 27076 10052
rect 26796 9716 26852 9726
rect 26460 9660 26628 9716
rect 26572 9210 26628 9660
rect 26796 9622 26852 9660
rect 26236 8990 26238 9042
rect 26290 8990 26292 9042
rect 26236 8978 26292 8990
rect 26460 9156 26516 9166
rect 26572 9158 26574 9210
rect 26626 9158 26628 9210
rect 26572 9146 26628 9158
rect 26124 8764 26404 8820
rect 25994 8726 26050 8764
rect 22204 8260 22260 8270
rect 22204 8166 22260 8204
rect 23324 8258 23380 8270
rect 23324 8206 23326 8258
rect 23378 8206 23380 8258
rect 23044 8148 23100 8158
rect 22876 8146 23100 8148
rect 22876 8094 23046 8146
rect 23098 8094 23100 8146
rect 22876 8092 23100 8094
rect 22540 8034 22596 8046
rect 22540 7982 22542 8034
rect 22594 7982 22596 8034
rect 22540 7588 22596 7982
rect 22540 7532 22820 7588
rect 21868 7422 21870 7474
rect 21922 7422 21924 7474
rect 21868 7410 21924 7422
rect 22652 7362 22708 7374
rect 22652 7310 22654 7362
rect 22706 7310 22708 7362
rect 22540 6916 22596 6926
rect 22652 6916 22708 7310
rect 22540 6914 22708 6916
rect 22540 6862 22542 6914
rect 22594 6862 22708 6914
rect 22540 6860 22708 6862
rect 22540 6850 22596 6860
rect 21756 6638 21758 6690
rect 21810 6638 21812 6690
rect 21756 6626 21812 6638
rect 21420 6188 21588 6244
rect 21420 6020 21476 6188
rect 21420 5926 21476 5964
rect 21756 6020 21812 6030
rect 21588 5906 21644 5918
rect 21588 5854 21590 5906
rect 21642 5854 21644 5906
rect 21196 5796 21252 5806
rect 21588 5796 21644 5854
rect 21196 5794 21644 5796
rect 21196 5742 21198 5794
rect 21250 5742 21644 5794
rect 21196 5740 21644 5742
rect 21196 5730 21252 5740
rect 21756 4450 21812 5964
rect 22092 6020 22148 6030
rect 22092 5906 22148 5964
rect 22092 5854 22094 5906
rect 22146 5854 22148 5906
rect 22092 5842 22148 5854
rect 22764 5908 22820 7532
rect 22876 6692 22932 8092
rect 23044 8082 23100 8092
rect 23324 7700 23380 8206
rect 23548 8260 23604 8270
rect 23548 8258 23828 8260
rect 23548 8206 23550 8258
rect 23602 8206 23828 8258
rect 23548 8204 23828 8206
rect 23548 8194 23604 8204
rect 23324 7634 23380 7644
rect 22876 6626 22932 6636
rect 22764 5814 22820 5852
rect 22876 5906 22932 5918
rect 22876 5854 22878 5906
rect 22930 5854 22932 5906
rect 22334 5684 22390 5694
rect 22876 5684 22932 5854
rect 23772 5796 23828 8204
rect 23996 6692 24052 6702
rect 23996 6598 24052 6636
rect 23772 5730 23828 5740
rect 24108 5906 24164 5918
rect 24108 5854 24110 5906
rect 24162 5854 24164 5906
rect 24108 5796 24164 5854
rect 24108 5730 24164 5740
rect 22334 5682 22932 5684
rect 22334 5630 22336 5682
rect 22388 5630 22932 5682
rect 22334 5628 22932 5630
rect 23156 5682 23212 5694
rect 23156 5630 23158 5682
rect 23210 5630 23212 5682
rect 22334 5618 22390 5628
rect 23156 5124 23212 5630
rect 23156 5058 23212 5068
rect 23660 5124 23716 5134
rect 23660 5030 23716 5068
rect 21756 4398 21758 4450
rect 21810 4398 21812 4450
rect 21756 4386 21812 4398
rect 22540 4898 22596 4910
rect 22540 4846 22542 4898
rect 22594 4846 22596 4898
rect 22540 4340 22596 4846
rect 22540 4274 22596 4284
rect 23660 4340 23716 4350
rect 23660 4246 23716 4284
rect 21196 4226 21252 4238
rect 21196 4174 21198 4226
rect 21250 4174 21252 4226
rect 21196 3780 21252 4174
rect 21196 3714 21252 3724
rect 22092 3668 22148 3678
rect 22092 3574 22148 3612
rect 22652 3668 22708 3678
rect 21084 3474 21086 3526
rect 21138 3474 21140 3526
rect 21084 3462 21140 3474
rect 22652 800 22708 3612
rect 24220 2548 24276 8372
rect 24556 7476 24612 7486
rect 24556 7382 24612 7420
rect 24522 7084 24786 7094
rect 24578 7028 24626 7084
rect 24682 7028 24730 7084
rect 24522 7018 24786 7028
rect 24668 6690 24724 6702
rect 24668 6638 24670 6690
rect 24722 6638 24724 6690
rect 24668 6030 24724 6638
rect 24612 6018 24724 6030
rect 24612 5966 24614 6018
rect 24666 5966 24724 6018
rect 24612 5964 24724 5966
rect 24612 5954 24668 5964
rect 24332 5908 24388 5918
rect 24332 5814 24388 5852
rect 24332 5684 24388 5694
rect 24332 2884 24388 5628
rect 24522 5516 24786 5526
rect 24578 5460 24626 5516
rect 24682 5460 24730 5516
rect 24522 5450 24786 5460
rect 24780 5124 24836 5134
rect 24892 5124 24948 8428
rect 25676 8372 26124 8428
rect 26068 8370 26124 8372
rect 26068 8318 26070 8370
rect 26122 8318 26124 8370
rect 26068 8306 26124 8318
rect 26348 8258 26404 8764
rect 26348 8206 26350 8258
rect 26402 8206 26404 8258
rect 26348 8194 26404 8206
rect 26460 8258 26516 9100
rect 26740 8986 26796 8998
rect 26740 8934 26742 8986
rect 26794 8934 26796 8986
rect 26740 8708 26796 8934
rect 26740 8652 26852 8708
rect 26796 8372 26852 8652
rect 26908 8596 26964 9996
rect 27300 9884 27356 9894
rect 27020 9882 27356 9884
rect 27020 9830 27302 9882
rect 27354 9830 27356 9882
rect 27020 9828 27356 9830
rect 27020 8820 27076 9828
rect 27300 9818 27356 9828
rect 27132 9714 27188 9726
rect 27132 9662 27134 9714
rect 27186 9662 27188 9714
rect 27132 9604 27188 9662
rect 27468 9604 27524 11340
rect 27804 10498 27860 10510
rect 27804 10446 27806 10498
rect 27858 10446 27860 10498
rect 27804 9884 27860 10446
rect 27916 10052 27972 15092
rect 28382 15090 28438 15102
rect 28382 15038 28384 15090
rect 28436 15038 28438 15090
rect 28382 14532 28438 15038
rect 28588 14532 28644 14542
rect 28382 14530 28644 14532
rect 28382 14478 28590 14530
rect 28642 14478 28644 14530
rect 28382 14476 28644 14478
rect 28588 14466 28644 14476
rect 28252 14306 28308 14318
rect 28252 14254 28254 14306
rect 28306 14254 28308 14306
rect 28028 13748 28084 13758
rect 28252 13748 28308 14254
rect 28812 14196 28868 15262
rect 29596 15314 29652 15820
rect 29596 15262 29598 15314
rect 29650 15262 29652 15314
rect 29596 15250 29652 15262
rect 29316 14644 29372 14654
rect 29316 14550 29372 14588
rect 28812 14130 28868 14140
rect 29184 14140 29448 14150
rect 29240 14084 29288 14140
rect 29344 14084 29392 14140
rect 29184 14074 29448 14084
rect 29708 13972 29764 16866
rect 30156 16918 30212 17164
rect 30156 16866 30158 16918
rect 30210 16866 30212 16918
rect 30156 16660 30212 16866
rect 30380 16884 30436 17724
rect 30492 17714 30548 17724
rect 30492 16996 30548 17006
rect 30492 16938 30548 16940
rect 30492 16886 30494 16938
rect 30546 16886 30548 16938
rect 30492 16874 30548 16886
rect 30380 16818 30436 16828
rect 30156 16594 30212 16604
rect 29708 13906 29764 13916
rect 29820 16548 29876 16558
rect 29820 13860 29876 16492
rect 29932 16212 29988 16222
rect 29932 16061 29988 16156
rect 29932 16009 29934 16061
rect 29986 16009 29988 16061
rect 29932 15997 29988 16009
rect 30380 16212 30436 16222
rect 30380 16065 30436 16156
rect 30380 16013 30382 16065
rect 30434 16013 30436 16065
rect 30380 16001 30436 16013
rect 30604 15876 30660 19012
rect 31008 18956 31332 19012
rect 31388 19404 31556 19460
rect 31008 18488 31064 18956
rect 31164 18788 31220 18798
rect 31220 18732 31332 18788
rect 31164 18722 31220 18732
rect 31008 18436 31010 18488
rect 31062 18436 31064 18488
rect 31008 18424 31064 18436
rect 31164 18450 31220 18462
rect 31164 18398 31166 18450
rect 31218 18398 31220 18450
rect 31164 18228 31220 18398
rect 31276 18340 31332 18732
rect 31388 18452 31444 19404
rect 31724 19348 31780 20638
rect 31836 19918 31892 20860
rect 31948 20132 32004 21422
rect 32060 20802 32116 22876
rect 32284 23154 32340 23166
rect 32284 23102 32286 23154
rect 32338 23102 32340 23154
rect 32284 22932 32340 23102
rect 32172 22484 32228 22522
rect 32172 22418 32228 22428
rect 32172 22314 32228 22326
rect 32172 22262 32174 22314
rect 32226 22262 32228 22314
rect 32172 22148 32228 22262
rect 32172 22082 32228 22092
rect 32284 22036 32340 22876
rect 32396 22986 32452 22998
rect 32396 22934 32398 22986
rect 32450 22934 32452 22986
rect 32396 22820 32452 22934
rect 32396 22754 32452 22764
rect 32508 22596 32564 22606
rect 32284 21970 32340 21980
rect 32396 22372 32452 22382
rect 32284 21588 32340 21598
rect 32284 21494 32340 21532
rect 32060 20750 32062 20802
rect 32114 20750 32116 20802
rect 32060 20738 32116 20750
rect 32284 20804 32340 20814
rect 32396 20804 32452 22316
rect 32508 22370 32564 22540
rect 32508 22318 32510 22370
rect 32562 22318 32564 22370
rect 32508 22306 32564 22318
rect 32620 21588 32676 24108
rect 32732 22820 32788 24332
rect 32732 21812 32788 22764
rect 32844 23604 32900 24556
rect 32844 22370 32900 23548
rect 32956 23492 33012 25004
rect 33404 24836 33460 24846
rect 33404 24722 33460 24780
rect 33404 24670 33406 24722
rect 33458 24670 33460 24722
rect 33404 24658 33460 24670
rect 32956 23426 33012 23436
rect 33516 22596 33572 25004
rect 33740 24946 33796 25004
rect 33740 24894 33742 24946
rect 33794 24894 33796 24946
rect 33740 24882 33796 24894
rect 33846 24332 34110 24342
rect 33902 24276 33950 24332
rect 34006 24276 34054 24332
rect 33846 24266 34110 24276
rect 33846 22764 34110 22774
rect 33902 22708 33950 22764
rect 34006 22708 34054 22764
rect 33846 22698 34110 22708
rect 34300 22596 34356 26852
rect 34412 25732 34468 27580
rect 34748 27300 34804 27310
rect 34860 27300 34916 28028
rect 34748 27298 34916 27300
rect 34748 27246 34750 27298
rect 34802 27246 34916 27298
rect 34748 27244 34916 27246
rect 34748 27234 34804 27244
rect 34412 25666 34468 25676
rect 34692 25396 34748 25406
rect 34692 24834 34748 25340
rect 34692 24782 34694 24834
rect 34746 24782 34748 24834
rect 34692 24770 34748 24782
rect 34972 24724 35028 29148
rect 35532 27746 35588 27758
rect 35532 27694 35534 27746
rect 35586 27694 35588 27746
rect 35532 26908 35588 27694
rect 35084 26852 35588 26908
rect 35084 26514 35140 26852
rect 35084 26462 35086 26514
rect 35138 26462 35140 26514
rect 35084 26450 35140 26462
rect 35756 26317 35812 30604
rect 36036 30324 36092 30334
rect 36036 30230 36092 30268
rect 36204 29764 36260 31164
rect 36092 29708 36260 29764
rect 36316 29764 36372 31276
rect 36092 29453 36148 29708
rect 36316 29698 36372 29708
rect 36092 29401 36094 29453
rect 36146 29401 36148 29453
rect 36092 29389 36148 29401
rect 36428 28614 36484 32060
rect 36540 30324 36596 32060
rect 36540 30258 36596 30268
rect 36428 28562 36430 28614
rect 36482 28562 36484 28614
rect 36428 28550 36484 28562
rect 36484 27076 36540 27086
rect 36484 26982 36540 27020
rect 36652 26908 36708 32172
rect 37156 31778 37212 31790
rect 37156 31726 37158 31778
rect 37210 31726 37212 31778
rect 36988 31666 37044 31678
rect 36988 31614 36990 31666
rect 37042 31614 37044 31666
rect 36988 31220 37044 31614
rect 37156 31444 37212 31726
rect 37156 31378 37212 31388
rect 37324 31332 37380 32732
rect 37436 31668 37492 33964
rect 37996 33908 38052 33918
rect 37996 33814 38052 33852
rect 37660 33348 37716 33358
rect 37660 33254 37716 33292
rect 38220 33348 38276 33358
rect 37902 33236 37958 33246
rect 37772 33234 37958 33236
rect 37772 33182 37904 33234
rect 37956 33182 37958 33234
rect 37772 33180 37958 33182
rect 37772 32614 37828 33180
rect 37902 33170 37958 33180
rect 38108 33236 38164 33246
rect 37436 31602 37492 31612
rect 37548 32558 37828 32614
rect 37324 31276 37492 31332
rect 37212 31220 37268 31230
rect 36988 31164 37156 31220
rect 36988 30996 37044 31006
rect 36988 30902 37044 30940
rect 37100 30436 37156 31164
rect 36988 30380 37156 30436
rect 37212 30436 37268 31164
rect 37324 31108 37380 31118
rect 37324 30994 37380 31052
rect 37324 30942 37326 30994
rect 37378 30942 37380 30994
rect 37324 30930 37380 30942
rect 37212 30380 37380 30436
rect 36988 30324 37044 30380
rect 36764 30268 37044 30324
rect 36764 29204 36820 30268
rect 37156 30212 37212 30222
rect 37156 30118 37212 30156
rect 36764 29110 36820 29148
rect 36988 30098 37044 30110
rect 36988 30046 36990 30098
rect 37042 30046 37044 30098
rect 36988 28756 37044 30046
rect 37324 29204 37380 30380
rect 36988 28690 37044 28700
rect 37156 29148 37380 29204
rect 37156 28698 37212 29148
rect 37156 28646 37158 28698
rect 37210 28646 37212 28698
rect 37156 28634 37212 28646
rect 37436 28644 37492 31276
rect 36988 28530 37044 28542
rect 36988 28478 36990 28530
rect 37042 28478 37044 28530
rect 36988 27076 37044 28478
rect 37436 27970 37492 28588
rect 37436 27918 37438 27970
rect 37490 27918 37492 27970
rect 37436 27906 37492 27918
rect 37548 27748 37604 32558
rect 37660 32452 37716 32462
rect 37660 31778 37716 32396
rect 37996 32452 38052 32462
rect 37996 32358 38052 32396
rect 37660 31726 37662 31778
rect 37714 31726 37716 31778
rect 37660 31108 37716 31726
rect 37902 31666 37958 31678
rect 37902 31614 37904 31666
rect 37956 31614 37958 31666
rect 37902 31108 37958 31614
rect 37660 31042 37716 31052
rect 37772 31052 37958 31108
rect 37660 30884 37716 30894
rect 37660 30790 37716 30828
rect 37660 30210 37716 30222
rect 37660 30158 37662 30210
rect 37714 30158 37716 30210
rect 37660 29988 37716 30158
rect 37660 29922 37716 29932
rect 37660 28644 37716 28654
rect 37772 28644 37828 31052
rect 37902 30100 37958 30110
rect 37902 30006 37958 30044
rect 38108 29428 38164 33180
rect 38220 30996 38276 33292
rect 38220 30930 38276 30940
rect 38220 29428 38276 29438
rect 38108 29426 38276 29428
rect 38108 29374 38222 29426
rect 38274 29374 38276 29426
rect 38108 29372 38276 29374
rect 38220 29204 38276 29372
rect 38332 29428 38388 34078
rect 39004 33908 39060 33918
rect 38508 32956 38772 32966
rect 38564 32900 38612 32956
rect 38668 32900 38716 32956
rect 38508 32890 38772 32900
rect 38508 31388 38772 31398
rect 38564 31332 38612 31388
rect 38668 31332 38716 31388
rect 38508 31322 38772 31332
rect 38508 29820 38772 29830
rect 38564 29764 38612 29820
rect 38668 29764 38716 29820
rect 38508 29754 38772 29764
rect 38332 29362 38388 29372
rect 38220 29148 38948 29204
rect 37660 28642 37828 28644
rect 37660 28590 37662 28642
rect 37714 28590 37828 28642
rect 37660 28588 37828 28590
rect 37660 28578 37716 28588
rect 37902 28532 37958 28542
rect 37772 28530 37958 28532
rect 37772 28478 37904 28530
rect 37956 28478 37958 28530
rect 37772 28476 37958 28478
rect 37772 27748 37828 28476
rect 37902 28466 37958 28476
rect 38508 28252 38772 28262
rect 38564 28196 38612 28252
rect 38668 28196 38716 28252
rect 38508 28186 38772 28196
rect 36876 27020 37044 27076
rect 37324 27692 37604 27748
rect 37660 27692 37828 27748
rect 38332 27858 38388 27870
rect 38332 27806 38334 27858
rect 38386 27806 38388 27858
rect 37324 27074 37380 27692
rect 37324 27022 37326 27074
rect 37378 27022 37380 27074
rect 36876 26964 36932 27020
rect 37324 27010 37380 27022
rect 36652 26852 36820 26908
rect 35756 26265 35758 26317
rect 35810 26265 35812 26317
rect 35756 26253 35812 26265
rect 36764 26178 36820 26852
rect 36876 26852 36932 26908
rect 37082 26964 37138 26974
rect 37082 26962 37268 26964
rect 37082 26910 37084 26962
rect 37136 26910 37268 26962
rect 37082 26908 37268 26910
rect 37082 26898 37138 26908
rect 37212 26852 37380 26908
rect 36876 26796 37044 26852
rect 36764 26126 36766 26178
rect 36818 26126 36820 26178
rect 36764 26114 36820 26126
rect 35756 25508 35812 25518
rect 36988 25508 37044 26796
rect 35364 25450 35420 25462
rect 35364 25398 35366 25450
rect 35418 25398 35420 25450
rect 35756 25414 35812 25452
rect 35980 25450 36036 25462
rect 35364 25396 35420 25398
rect 35364 25330 35420 25340
rect 35532 25396 35588 25406
rect 35532 25302 35588 25340
rect 35980 25398 35982 25450
rect 36034 25398 36036 25450
rect 35980 25060 36036 25398
rect 36876 25452 37044 25508
rect 37324 25506 37380 26852
rect 37660 26180 37716 27692
rect 37996 27636 38052 27646
rect 37996 27634 38276 27636
rect 37996 27582 37998 27634
rect 38050 27582 38276 27634
rect 37996 27580 38276 27582
rect 37996 27570 38052 27580
rect 37828 27132 38164 27188
rect 37828 27130 37884 27132
rect 37828 27078 37830 27130
rect 37882 27078 37884 27130
rect 37828 27066 37884 27078
rect 37996 26964 38052 27002
rect 37996 26898 38052 26908
rect 37660 26124 37884 26180
rect 37324 25454 37326 25506
rect 37378 25454 37380 25506
rect 37828 25562 37884 26124
rect 37828 25510 37830 25562
rect 37882 25510 37884 25562
rect 37828 25498 37884 25510
rect 36036 25004 36260 25060
rect 35980 24994 36036 25004
rect 34972 24630 35028 24668
rect 35196 24836 35252 24846
rect 35196 24722 35252 24780
rect 35196 24670 35198 24722
rect 35250 24670 35252 24722
rect 34580 24164 34636 24174
rect 34580 24050 34636 24108
rect 34580 23998 34582 24050
rect 34634 23998 34636 24050
rect 34580 23986 34636 23998
rect 34860 24050 34916 24062
rect 34860 23998 34862 24050
rect 34914 23998 34916 24050
rect 34860 23380 34916 23998
rect 34972 23894 35028 23906
rect 34972 23842 34974 23894
rect 35026 23842 35028 23894
rect 34972 23828 35028 23842
rect 34972 23762 35028 23772
rect 35196 23604 35252 24670
rect 36204 24612 36260 25004
rect 36876 24836 36932 25452
rect 37324 25442 37380 25454
rect 37082 25396 37138 25406
rect 37082 25394 37268 25396
rect 37082 25342 37084 25394
rect 37136 25342 37268 25394
rect 37082 25340 37268 25342
rect 37082 25330 37138 25340
rect 37212 24948 37268 25340
rect 37996 25394 38052 25406
rect 37996 25342 37998 25394
rect 38050 25342 38052 25394
rect 37212 24892 37828 24948
rect 36876 24770 36932 24780
rect 37212 24724 37268 24734
rect 37212 24630 37268 24668
rect 37436 24724 37492 24734
rect 36204 24546 36260 24556
rect 36092 24500 36148 24510
rect 35980 24498 36148 24500
rect 35980 24446 36094 24498
rect 36146 24446 36148 24498
rect 35980 24444 36148 24446
rect 35308 24164 35364 24174
rect 35308 23938 35364 24108
rect 35308 23886 35310 23938
rect 35362 23886 35364 23938
rect 35308 23874 35364 23886
rect 35420 24052 35476 24062
rect 35196 23538 35252 23548
rect 35420 23380 35476 23996
rect 35644 24052 35700 24062
rect 35644 23938 35700 23996
rect 35644 23886 35646 23938
rect 35698 23886 35700 23938
rect 35644 23874 35700 23886
rect 35756 23994 35868 24052
rect 35756 23942 35814 23994
rect 35866 23942 35868 23994
rect 35756 23930 35868 23942
rect 35980 23940 36036 24444
rect 36092 24434 36148 24444
rect 35756 23716 35812 23930
rect 35980 23846 36036 23884
rect 36092 23940 36148 23950
rect 36372 23940 36428 23950
rect 36092 23938 36260 23940
rect 36092 23886 36094 23938
rect 36146 23886 36260 23938
rect 36092 23884 36260 23886
rect 36092 23874 36148 23884
rect 35644 23660 35812 23716
rect 35420 23324 35588 23380
rect 34860 23314 34916 23324
rect 34524 23156 34580 23166
rect 34524 23062 34580 23100
rect 35420 23156 35476 23166
rect 35420 23062 35476 23100
rect 34860 22932 34916 22942
rect 34860 22838 34916 22876
rect 33572 22540 33796 22596
rect 33516 22530 33572 22540
rect 32844 22318 32846 22370
rect 32898 22318 32900 22370
rect 32844 22306 32900 22318
rect 33404 22484 33460 22494
rect 33404 22370 33460 22428
rect 33404 22318 33406 22370
rect 33458 22318 33460 22370
rect 33740 22372 33796 22540
rect 33404 22306 33460 22318
rect 33572 22314 33628 22326
rect 33572 22262 33574 22314
rect 33626 22262 33628 22314
rect 33572 21812 33628 22262
rect 32732 21746 32788 21756
rect 33348 21756 33628 21812
rect 33348 21698 33404 21756
rect 33348 21646 33350 21698
rect 33402 21646 33404 21698
rect 33348 21634 33404 21646
rect 32620 21522 32676 21532
rect 33628 21586 33684 21598
rect 33628 21534 33630 21586
rect 33682 21534 33684 21586
rect 32284 20802 32452 20804
rect 32284 20750 32286 20802
rect 32338 20750 32452 20802
rect 32284 20748 32452 20750
rect 33516 21364 33572 21374
rect 32284 20738 32340 20748
rect 32564 20690 32620 20702
rect 32564 20638 32566 20690
rect 32618 20638 32620 20690
rect 32564 20356 32620 20638
rect 33516 20580 33572 21308
rect 33628 20804 33684 21534
rect 33740 21586 33796 22316
rect 34076 22540 34356 22596
rect 34076 22370 34132 22540
rect 34076 22318 34078 22370
rect 34130 22318 34132 22370
rect 33740 21534 33742 21586
rect 33794 21534 33796 21586
rect 33740 21522 33796 21534
rect 33964 22260 34020 22270
rect 33964 21586 34020 22204
rect 33964 21534 33966 21586
rect 34018 21534 34020 21586
rect 33964 21522 34020 21534
rect 34076 21364 34132 22318
rect 34636 22372 34692 22382
rect 34636 22278 34692 22316
rect 34860 22370 34916 22382
rect 34860 22318 34862 22370
rect 34914 22318 34916 22370
rect 34318 22260 34374 22270
rect 34318 22166 34374 22204
rect 34076 21308 34244 21364
rect 33846 21196 34110 21206
rect 33902 21140 33950 21196
rect 34006 21140 34054 21196
rect 33846 21130 34110 21140
rect 34188 21028 34244 21308
rect 34860 21140 34916 22318
rect 35140 22260 35196 22270
rect 34972 22258 35196 22260
rect 34972 22206 35142 22258
rect 35194 22206 35196 22258
rect 34972 22204 35196 22206
rect 34972 21364 35028 22204
rect 35140 22194 35196 22204
rect 35532 21476 35588 23324
rect 35644 22932 35700 23660
rect 35868 23604 35924 23614
rect 35756 23548 35868 23604
rect 35756 23154 35812 23548
rect 35868 23538 35924 23548
rect 36204 23268 36260 23884
rect 36372 23846 36428 23884
rect 37324 23940 37380 23950
rect 37324 23846 37380 23884
rect 37082 23826 37138 23838
rect 37082 23774 37084 23826
rect 37136 23774 37138 23826
rect 37082 23716 37138 23774
rect 36988 23660 37138 23716
rect 37436 23828 37492 24668
rect 37548 24612 37604 24622
rect 37548 24518 37604 24556
rect 37772 24500 37828 24892
rect 37884 24836 37940 24846
rect 37884 24722 37940 24780
rect 37884 24670 37886 24722
rect 37938 24670 37940 24722
rect 37884 24658 37940 24670
rect 37996 24612 38052 25342
rect 37996 24546 38052 24556
rect 37772 24444 37884 24500
rect 37828 23994 37884 24444
rect 37828 23942 37830 23994
rect 37882 23942 37884 23994
rect 37828 23930 37884 23942
rect 37996 24164 38052 24174
rect 37996 23938 38052 24108
rect 37996 23886 37998 23938
rect 38050 23886 38052 23938
rect 37996 23874 38052 23886
rect 36410 23268 36466 23278
rect 36204 23266 36466 23268
rect 36204 23214 36412 23266
rect 36464 23214 36466 23266
rect 36204 23212 36466 23214
rect 36410 23202 36466 23212
rect 36652 23156 36708 23166
rect 35756 23102 35758 23154
rect 35810 23102 35812 23154
rect 35756 23090 35812 23102
rect 36540 23154 36708 23156
rect 36540 23102 36654 23154
rect 36706 23102 36708 23154
rect 36540 23100 36708 23102
rect 35644 22866 35700 22876
rect 35980 21586 36036 21598
rect 35980 21534 35982 21586
rect 36034 21534 36036 21586
rect 35532 21420 35924 21476
rect 34972 21298 35028 21308
rect 35420 21364 35476 21374
rect 35420 21362 35812 21364
rect 35420 21310 35422 21362
rect 35474 21310 35812 21362
rect 35420 21308 35812 21310
rect 35420 21298 35476 21308
rect 34860 21074 34916 21084
rect 35644 21140 35700 21150
rect 33964 20972 34244 21028
rect 33852 20804 33908 20814
rect 33628 20748 33852 20804
rect 33852 20710 33908 20748
rect 32564 20290 32620 20300
rect 33460 20524 33572 20580
rect 33292 20132 33348 20142
rect 31948 20130 33348 20132
rect 31948 20078 33294 20130
rect 33346 20078 33348 20130
rect 31948 20076 33348 20078
rect 33292 20066 33348 20076
rect 33460 20074 33516 20524
rect 33460 20022 33462 20074
rect 33514 20022 33516 20074
rect 33460 20010 33516 20022
rect 33964 20018 34020 20972
rect 34206 20356 34262 20366
rect 34206 20130 34262 20300
rect 34206 20078 34208 20130
rect 34260 20078 34262 20130
rect 34206 20066 34262 20078
rect 35644 20130 35700 21084
rect 35756 20914 35812 21308
rect 35756 20862 35758 20914
rect 35810 20862 35812 20914
rect 35756 20850 35812 20862
rect 35644 20078 35646 20130
rect 35698 20078 35700 20130
rect 35644 20066 35700 20078
rect 33964 19966 33966 20018
rect 34018 19966 34020 20018
rect 33964 19954 34020 19966
rect 31836 19906 31948 19918
rect 31836 19854 31894 19906
rect 31946 19854 31948 19906
rect 31836 19852 31948 19854
rect 31892 19842 31948 19852
rect 32060 19908 32116 19918
rect 31612 19292 31780 19348
rect 31892 19684 31948 19694
rect 31388 18396 31556 18452
rect 31276 18284 31388 18340
rect 31332 18282 31388 18284
rect 31332 18230 31334 18282
rect 31386 18230 31388 18282
rect 31332 18218 31388 18230
rect 31164 18162 31220 18172
rect 31108 17780 31164 17790
rect 31108 17106 31164 17724
rect 31108 17054 31110 17106
rect 31162 17054 31164 17106
rect 31108 16996 31164 17054
rect 31108 16930 31164 16940
rect 30716 16548 30772 16558
rect 30716 16098 30772 16492
rect 30716 16046 30718 16098
rect 30770 16046 30772 16098
rect 30716 16034 30772 16046
rect 30828 16436 30884 16446
rect 30828 16098 30884 16380
rect 31388 16212 31444 16222
rect 31388 16118 31444 16156
rect 30828 16046 30830 16098
rect 30882 16046 30884 16098
rect 30828 16034 30884 16046
rect 30994 16100 31050 16110
rect 30994 16006 31050 16044
rect 30604 15820 30772 15876
rect 29932 13860 29988 13870
rect 30716 13860 30772 15820
rect 31500 15764 31556 18396
rect 29820 13858 29988 13860
rect 29820 13806 29934 13858
rect 29986 13806 29988 13858
rect 29820 13804 29988 13806
rect 29932 13794 29988 13804
rect 30492 13804 30772 13860
rect 30828 15708 31556 15764
rect 28028 13746 28308 13748
rect 28028 13694 28030 13746
rect 28082 13694 28308 13746
rect 28028 13692 28308 13694
rect 28028 13682 28084 13692
rect 29932 13524 29988 13534
rect 28700 12962 28756 12974
rect 28700 12910 28702 12962
rect 28754 12910 28756 12962
rect 28588 12292 28644 12302
rect 28588 12205 28644 12236
rect 28588 12153 28590 12205
rect 28642 12153 28644 12205
rect 28084 11508 28140 11518
rect 28084 11414 28140 11452
rect 28588 11508 28644 12153
rect 28700 11732 28756 12910
rect 29596 12964 29652 12974
rect 29596 12870 29652 12908
rect 29932 12962 29988 13468
rect 30156 13412 30212 13422
rect 29932 12910 29934 12962
rect 29986 12910 29988 12962
rect 29932 12898 29988 12910
rect 30044 12962 30100 12974
rect 30044 12910 30046 12962
rect 30098 12910 30100 12962
rect 29184 12572 29448 12582
rect 29240 12516 29288 12572
rect 29344 12516 29392 12572
rect 29184 12506 29448 12516
rect 28700 11666 28756 11676
rect 29372 11956 29428 11966
rect 30044 11956 30100 12910
rect 29372 11954 30100 11956
rect 29372 11902 29374 11954
rect 29426 11902 30100 11954
rect 29372 11900 30100 11902
rect 29372 11732 29428 11900
rect 30156 11844 30212 13356
rect 30492 12404 30548 13804
rect 30660 13636 30716 13646
rect 30660 13542 30716 13580
rect 30828 13188 30884 15708
rect 31388 15540 31444 15550
rect 31388 15148 31444 15484
rect 31500 15428 31556 15438
rect 31500 15334 31556 15372
rect 31388 15092 31556 15148
rect 31500 14530 31556 15092
rect 31500 14478 31502 14530
rect 31554 14478 31556 14530
rect 31276 13746 31332 13758
rect 31276 13694 31278 13746
rect 31330 13694 31332 13746
rect 30996 13524 31052 13534
rect 30996 13430 31052 13468
rect 31164 13524 31220 13534
rect 31164 13300 31220 13468
rect 30492 12338 30548 12348
rect 30716 13132 30884 13188
rect 31052 13244 31220 13300
rect 31276 13300 31332 13694
rect 31388 13746 31444 13758
rect 31388 13694 31390 13746
rect 31442 13694 31444 13746
rect 31388 13636 31444 13694
rect 31388 13570 31444 13580
rect 31500 13412 31556 14478
rect 31612 13748 31668 19292
rect 31892 19290 31948 19628
rect 31892 19238 31894 19290
rect 31946 19238 31948 19290
rect 31892 19226 31948 19238
rect 31724 19122 31780 19134
rect 31724 19070 31726 19122
rect 31778 19070 31780 19122
rect 31724 16884 31780 19070
rect 31724 16818 31780 16828
rect 31836 19124 31892 19134
rect 31724 16660 31780 16670
rect 31724 15428 31780 16604
rect 31836 15540 31892 19068
rect 32060 17780 32116 19852
rect 34636 19908 34692 19918
rect 32340 19684 32396 19694
rect 32340 19346 32396 19628
rect 33846 19628 34110 19638
rect 33902 19572 33950 19628
rect 34006 19572 34054 19628
rect 33846 19562 34110 19572
rect 32340 19294 32342 19346
rect 32394 19294 32396 19346
rect 32340 19282 32396 19294
rect 33964 18450 34020 18462
rect 33964 18398 33966 18450
rect 34018 18398 34020 18450
rect 33796 18340 33852 18350
rect 33964 18340 34020 18398
rect 33796 18338 34020 18340
rect 33796 18286 33798 18338
rect 33850 18286 34020 18338
rect 33796 18284 34020 18286
rect 34188 18450 34244 18462
rect 34188 18398 34190 18450
rect 34242 18398 34244 18450
rect 33796 18228 33852 18284
rect 32060 17714 32116 17724
rect 33516 18172 33852 18228
rect 32172 16884 32228 16894
rect 32004 16660 32060 16670
rect 32004 16436 32060 16604
rect 32004 16210 32060 16380
rect 32004 16158 32006 16210
rect 32058 16158 32060 16210
rect 32004 16146 32060 16158
rect 31836 15474 31892 15484
rect 31724 15362 31780 15372
rect 31836 14306 31892 14318
rect 31836 14254 31838 14306
rect 31890 14254 31892 14306
rect 31836 13748 31892 14254
rect 31836 13692 32004 13748
rect 31612 13682 31668 13692
rect 31612 13524 31668 13534
rect 31836 13524 31892 13534
rect 31668 13522 31892 13524
rect 31668 13470 31838 13522
rect 31890 13470 31892 13522
rect 31668 13468 31892 13470
rect 31612 13458 31668 13468
rect 31836 13458 31892 13468
rect 31500 13346 31556 13356
rect 29372 11666 29428 11676
rect 30044 11788 30212 11844
rect 28588 11442 28644 11452
rect 29596 11340 29876 11396
rect 29184 11004 29448 11014
rect 29240 10948 29288 11004
rect 29344 10948 29392 11004
rect 29184 10938 29448 10948
rect 29596 10734 29652 11340
rect 29708 11170 29764 11182
rect 29708 11118 29710 11170
rect 29762 11118 29764 11170
rect 29708 10836 29764 11118
rect 29820 11172 29876 11340
rect 30044 11394 30100 11788
rect 30044 11342 30046 11394
rect 30098 11342 30100 11394
rect 30044 11330 30100 11342
rect 30156 11394 30212 11406
rect 30156 11342 30158 11394
rect 30210 11342 30212 11394
rect 30156 11172 30212 11342
rect 29820 11116 30212 11172
rect 30492 11172 30548 11182
rect 30492 11078 30548 11116
rect 29708 10780 29988 10836
rect 29540 10722 29652 10734
rect 29540 10670 29542 10722
rect 29594 10670 29652 10722
rect 29540 10668 29652 10670
rect 29540 10658 29596 10668
rect 28700 10612 28756 10622
rect 28588 10610 28756 10612
rect 28588 10558 28702 10610
rect 28754 10558 28756 10610
rect 28588 10556 28756 10558
rect 27916 9986 27972 9996
rect 28364 10386 28420 10398
rect 28364 10334 28366 10386
rect 28418 10334 28420 10386
rect 27804 9828 28308 9884
rect 27804 9826 27860 9828
rect 27804 9774 27806 9826
rect 27858 9774 27860 9826
rect 27804 9762 27860 9774
rect 28046 9716 28102 9726
rect 27132 9538 27188 9548
rect 27300 9548 27524 9604
rect 27916 9714 28102 9716
rect 27916 9662 28048 9714
rect 28100 9662 28102 9714
rect 27916 9660 28102 9662
rect 27300 9154 27356 9548
rect 27916 9380 27972 9660
rect 28046 9650 28102 9660
rect 27300 9102 27302 9154
rect 27354 9102 27356 9154
rect 27300 9090 27356 9102
rect 27580 9324 27972 9380
rect 27580 9042 27636 9324
rect 27580 8990 27582 9042
rect 27634 8990 27636 9042
rect 27580 8978 27636 8990
rect 27804 9156 27860 9166
rect 27804 9042 27860 9100
rect 27804 8990 27806 9042
rect 27858 8990 27860 9042
rect 27804 8978 27860 8990
rect 28122 9044 28178 9054
rect 28252 9044 28308 9828
rect 28364 9828 28420 10334
rect 28364 9268 28420 9772
rect 28364 9202 28420 9212
rect 28364 9044 28420 9054
rect 28252 9042 28420 9044
rect 28252 8990 28366 9042
rect 28418 8990 28420 9042
rect 28252 8988 28420 8990
rect 28122 8950 28178 8988
rect 28364 8978 28420 8988
rect 27020 8754 27076 8764
rect 26908 8540 27300 8596
rect 26908 8372 26964 8382
rect 26796 8316 26908 8372
rect 26908 8306 26964 8316
rect 27132 8260 27188 8270
rect 26460 8206 26462 8258
rect 26514 8206 26516 8258
rect 26460 8194 26516 8206
rect 27020 8258 27188 8260
rect 27020 8206 27134 8258
rect 27186 8206 27188 8258
rect 27020 8204 27188 8206
rect 26852 8148 26908 8158
rect 26572 8146 26908 8148
rect 26572 8094 26854 8146
rect 26906 8094 26908 8146
rect 26572 8092 26908 8094
rect 26572 7812 26628 8092
rect 26852 8082 26908 8092
rect 26180 7756 26628 7812
rect 25434 7700 25490 7710
rect 25434 7586 25490 7644
rect 25434 7534 25436 7586
rect 25488 7534 25490 7586
rect 25434 7522 25490 7534
rect 26180 7530 26236 7756
rect 27020 7642 27076 8204
rect 27132 8194 27188 8204
rect 27244 8258 27300 8540
rect 27244 8206 27246 8258
rect 27298 8206 27300 8258
rect 25676 7476 25732 7486
rect 26180 7478 26182 7530
rect 26234 7478 26236 7530
rect 26348 7588 26404 7598
rect 26348 7494 26404 7532
rect 27020 7590 27022 7642
rect 27074 7590 27076 7642
rect 26180 7466 26236 7478
rect 25676 7382 25732 7420
rect 26852 7418 26908 7430
rect 26852 7366 26854 7418
rect 26906 7366 26908 7418
rect 26852 7364 26908 7366
rect 26852 7298 26908 7308
rect 27020 6916 27076 7590
rect 27020 6850 27076 6860
rect 26684 6690 26740 6702
rect 26684 6638 26686 6690
rect 26738 6638 26740 6690
rect 25788 6468 25844 6478
rect 25564 6466 25844 6468
rect 25564 6414 25790 6466
rect 25842 6414 25844 6466
rect 25564 6412 25844 6414
rect 25228 6020 25284 6030
rect 25228 5933 25284 5964
rect 25228 5881 25230 5933
rect 25282 5881 25284 5933
rect 25228 5869 25284 5881
rect 25564 5234 25620 6412
rect 25788 6402 25844 6412
rect 25564 5182 25566 5234
rect 25618 5182 25620 5234
rect 25564 5170 25620 5182
rect 25788 5796 25844 5806
rect 24444 5122 24948 5124
rect 24444 5070 24782 5122
rect 24834 5070 24948 5122
rect 24444 5068 24948 5070
rect 24444 4340 24500 5068
rect 24780 5058 24836 5068
rect 25788 4340 25844 5740
rect 26236 5684 26292 5694
rect 26236 5590 26292 5628
rect 26236 4900 26292 4910
rect 26012 4340 26068 4350
rect 25788 4338 26068 4340
rect 25788 4286 26014 4338
rect 26066 4286 26068 4338
rect 25788 4284 26068 4286
rect 24444 4246 24500 4284
rect 26012 4274 26068 4284
rect 26236 4338 26292 4844
rect 26516 4452 26572 4462
rect 26684 4452 26740 6638
rect 26516 4450 26740 4452
rect 26516 4398 26518 4450
rect 26570 4398 26740 4450
rect 26516 4396 26740 4398
rect 26516 4386 26572 4396
rect 26236 4286 26238 4338
rect 26290 4286 26292 4338
rect 26236 4274 26292 4286
rect 26908 4340 26964 4350
rect 26908 4246 26964 4284
rect 24522 3948 24786 3958
rect 24578 3892 24626 3948
rect 24682 3892 24730 3948
rect 24522 3882 24786 3892
rect 24556 3780 24612 3790
rect 27244 3780 27300 8206
rect 27468 8372 27524 8382
rect 27356 7476 27412 7486
rect 27356 7382 27412 7420
rect 27468 7364 27524 8316
rect 28588 8260 28644 10556
rect 28700 10546 28756 10556
rect 29148 10610 29204 10622
rect 29148 10558 29150 10610
rect 29202 10558 29204 10610
rect 29036 10164 29092 10174
rect 29036 9154 29092 10108
rect 29148 9828 29204 10558
rect 29260 10612 29316 10622
rect 29260 10610 29428 10612
rect 29260 10558 29262 10610
rect 29314 10558 29428 10610
rect 29260 10556 29428 10558
rect 29260 10546 29316 10556
rect 29260 10388 29316 10398
rect 29260 9938 29316 10332
rect 29260 9886 29262 9938
rect 29314 9886 29316 9938
rect 29260 9874 29316 9886
rect 29148 9762 29204 9772
rect 29372 9604 29428 10556
rect 29932 10610 29988 10780
rect 29932 10558 29934 10610
rect 29986 10558 29988 10610
rect 30604 10610 30660 10622
rect 29708 10388 29764 10398
rect 29372 9548 29652 9604
rect 29184 9436 29448 9446
rect 29240 9380 29288 9436
rect 29344 9380 29392 9436
rect 29184 9370 29448 9380
rect 29036 9102 29038 9154
rect 29090 9102 29092 9154
rect 29036 9090 29092 9102
rect 29466 9156 29522 9166
rect 29596 9156 29652 9548
rect 29466 9154 29652 9156
rect 29466 9102 29468 9154
rect 29520 9102 29652 9154
rect 29466 9100 29652 9102
rect 29466 9090 29522 9100
rect 29708 9042 29764 10332
rect 29932 10164 29988 10558
rect 30100 10554 30156 10566
rect 30100 10502 30102 10554
rect 30154 10502 30156 10554
rect 30100 10164 30156 10502
rect 30604 10558 30606 10610
rect 30658 10558 30660 10610
rect 30604 10388 30660 10558
rect 30604 10322 30660 10332
rect 30716 10276 30772 13132
rect 30828 12964 30884 12974
rect 30828 12870 30884 12908
rect 31052 12292 31108 13244
rect 31276 13234 31332 13244
rect 31948 13076 32004 13692
rect 32172 13746 32228 16828
rect 32844 16884 32900 16894
rect 32844 16098 32900 16828
rect 33516 16324 33572 18172
rect 33846 18060 34110 18070
rect 33902 18004 33950 18060
rect 34006 18004 34054 18060
rect 33846 17994 34110 18004
rect 33684 17640 33740 17652
rect 33684 17588 33686 17640
rect 33738 17588 33740 17640
rect 33684 17108 33740 17588
rect 34188 17332 34244 18398
rect 34468 18452 34524 18462
rect 34468 18358 34524 18396
rect 34412 18228 34468 18238
rect 34412 17778 34468 18172
rect 34412 17726 34414 17778
rect 34466 17726 34468 17778
rect 34412 17714 34468 17726
rect 34188 17266 34244 17276
rect 33684 17106 34580 17108
rect 33684 17054 33686 17106
rect 33738 17054 34580 17106
rect 33684 17052 34580 17054
rect 33684 16324 33740 17052
rect 34412 16882 34468 16894
rect 34412 16830 34414 16882
rect 34466 16830 34468 16882
rect 34076 16772 34132 16782
rect 34076 16678 34132 16716
rect 33846 16492 34110 16502
rect 33902 16436 33950 16492
rect 34006 16436 34054 16492
rect 33846 16426 34110 16436
rect 34412 16324 34468 16830
rect 34524 16884 34580 17052
rect 34636 16884 34692 19852
rect 35252 19908 35308 19918
rect 35252 19814 35308 19852
rect 35868 19348 35924 21420
rect 35980 20356 36036 21534
rect 36540 21028 36596 23100
rect 36652 23090 36708 23100
rect 36988 21140 37044 23660
rect 37156 23492 37212 23502
rect 37156 23210 37212 23436
rect 37156 23158 37158 23210
rect 37210 23158 37212 23210
rect 37324 23268 37380 23278
rect 37436 23268 37492 23772
rect 37996 23604 38052 23614
rect 37996 23378 38052 23548
rect 37996 23326 37998 23378
rect 38050 23326 38052 23378
rect 37996 23314 38052 23326
rect 37324 23266 37492 23268
rect 37324 23214 37326 23266
rect 37378 23214 37492 23266
rect 37324 23212 37492 23214
rect 37324 23202 37380 23212
rect 37156 23146 37212 23158
rect 37436 21362 37492 21374
rect 37436 21310 37438 21362
rect 37490 21310 37492 21362
rect 36988 21084 37380 21140
rect 35980 20290 36036 20300
rect 36316 20972 36596 21028
rect 35868 19292 35980 19348
rect 34748 18452 34804 18462
rect 34748 18358 34804 18396
rect 35756 18450 35812 18462
rect 35756 18398 35758 18450
rect 35810 18398 35812 18450
rect 35084 18228 35140 18238
rect 35084 18134 35140 18172
rect 34524 16882 34692 16884
rect 34524 16830 34526 16882
rect 34578 16830 34692 16882
rect 34524 16828 34692 16830
rect 35084 17332 35140 17342
rect 35756 17332 35812 18398
rect 35924 18282 35980 19292
rect 35924 18230 35926 18282
rect 35978 18230 35980 18282
rect 35924 18218 35980 18230
rect 36316 17780 36372 20972
rect 36988 20916 37044 20926
rect 36540 20804 36596 20814
rect 36428 20802 36596 20804
rect 36428 20750 36542 20802
rect 36594 20750 36596 20802
rect 36428 20748 36596 20750
rect 36428 19908 36484 20748
rect 36540 20738 36596 20748
rect 36988 20802 37044 20860
rect 36988 20750 36990 20802
rect 37042 20750 37044 20802
rect 36988 20738 37044 20750
rect 37156 20804 37212 20814
rect 37156 20710 37212 20748
rect 36428 19460 36484 19852
rect 36428 19394 36484 19404
rect 37156 19460 37212 19470
rect 37156 19346 37212 19404
rect 37156 19294 37158 19346
rect 37210 19294 37212 19346
rect 37156 17780 37212 19294
rect 36316 17724 36708 17780
rect 36316 17554 36372 17566
rect 36316 17502 36318 17554
rect 36370 17502 36372 17554
rect 36316 17332 36372 17502
rect 34524 16818 34580 16828
rect 35084 16334 35140 17276
rect 35532 17276 36372 17332
rect 35308 16772 35364 16782
rect 35308 16678 35364 16716
rect 33516 16258 33572 16268
rect 33628 16268 33852 16324
rect 32844 16046 32846 16098
rect 32898 16046 32900 16098
rect 32844 16034 32900 16046
rect 33180 15876 33236 15886
rect 33180 15782 33236 15820
rect 32956 15314 33012 15326
rect 32956 15262 32958 15314
rect 33010 15262 33012 15314
rect 32340 15202 32396 15214
rect 32340 15150 32342 15202
rect 32394 15150 32396 15202
rect 32340 15148 32396 15150
rect 32340 15092 32676 15148
rect 32172 13694 32174 13746
rect 32226 13694 32228 13746
rect 32172 13682 32228 13694
rect 32620 14502 32676 15092
rect 32956 15092 33012 15262
rect 32956 15026 33012 15036
rect 33628 15092 33684 16268
rect 33796 16210 33852 16268
rect 34412 16258 34468 16268
rect 35066 16322 35140 16334
rect 35066 16270 35068 16322
rect 35120 16270 35140 16322
rect 35066 16268 35140 16270
rect 35066 16258 35122 16268
rect 33796 16158 33798 16210
rect 33850 16158 33852 16210
rect 33796 16146 33852 16158
rect 34524 16100 34580 16110
rect 34412 16098 34580 16100
rect 34412 16046 34526 16098
rect 34578 16046 34580 16098
rect 34412 16044 34580 16046
rect 33852 15876 33908 15886
rect 33852 15426 33908 15820
rect 34188 15876 34244 15886
rect 34188 15874 34356 15876
rect 34188 15822 34190 15874
rect 34242 15822 34356 15874
rect 34188 15820 34356 15822
rect 34188 15810 34244 15820
rect 33852 15374 33854 15426
rect 33906 15374 33908 15426
rect 33852 15204 33908 15374
rect 33852 15138 33908 15148
rect 34020 15258 34076 15270
rect 34020 15206 34022 15258
rect 34074 15206 34076 15258
rect 32620 14450 32622 14502
rect 32674 14450 32676 14502
rect 31948 13010 32004 13020
rect 32060 13300 32116 13310
rect 31612 12740 31668 12750
rect 31164 12292 31220 12302
rect 31052 12290 31556 12292
rect 31052 12238 31166 12290
rect 31218 12238 31556 12290
rect 31052 12236 31556 12238
rect 31164 12226 31220 12236
rect 31332 12122 31388 12134
rect 31332 12070 31334 12122
rect 31386 12070 31388 12122
rect 31332 11508 31388 12070
rect 30940 11452 31388 11508
rect 30940 11284 30996 11452
rect 30846 11228 30996 11284
rect 30846 10722 30902 11228
rect 30846 10670 30848 10722
rect 30900 10670 30902 10722
rect 30846 10658 30902 10670
rect 31164 11172 31220 11182
rect 30716 10220 30996 10276
rect 29932 10098 29988 10108
rect 30044 10108 30156 10164
rect 30044 9940 30100 10108
rect 28868 8988 28924 8998
rect 28588 8194 28644 8204
rect 28700 8986 28924 8988
rect 28700 8934 28870 8986
rect 28922 8934 28924 8986
rect 29708 8990 29710 9042
rect 29762 8990 29764 9042
rect 29708 8978 29764 8990
rect 29932 9884 30100 9940
rect 28700 8932 28924 8934
rect 28588 7588 28644 7598
rect 27468 5796 27524 7308
rect 28364 7474 28420 7486
rect 28364 7422 28366 7474
rect 28418 7422 28420 7474
rect 27598 7252 27654 7262
rect 28122 7252 28178 7262
rect 27580 7250 27654 7252
rect 27580 7198 27600 7250
rect 27652 7198 27654 7250
rect 27580 7186 27654 7198
rect 27916 7250 28178 7252
rect 27916 7198 28124 7250
rect 28176 7198 28178 7250
rect 27916 7196 28178 7198
rect 27580 6020 27636 7186
rect 27580 5954 27636 5964
rect 27804 6466 27860 6478
rect 27804 6414 27806 6466
rect 27858 6414 27860 6466
rect 27468 5740 27636 5796
rect 27468 5236 27524 5246
rect 27468 5142 27524 5180
rect 27468 3780 27524 3790
rect 27244 3778 27524 3780
rect 27244 3726 27470 3778
rect 27522 3726 27524 3778
rect 27244 3724 27524 3726
rect 27580 3780 27636 5740
rect 27692 4340 27748 4350
rect 27804 4340 27860 6414
rect 27916 5124 27972 7196
rect 28122 7186 28178 7196
rect 28364 6692 28420 7422
rect 28364 6626 28420 6636
rect 28122 5908 28178 5918
rect 28122 5814 28178 5852
rect 28364 5908 28420 5918
rect 28588 5908 28644 7532
rect 28700 6132 28756 8932
rect 28868 8922 28924 8932
rect 29036 8260 29092 8270
rect 29036 8166 29092 8204
rect 29372 8036 29428 8046
rect 29372 8034 29876 8036
rect 29372 7982 29374 8034
rect 29426 7982 29876 8034
rect 29372 7980 29876 7982
rect 29372 7970 29428 7980
rect 29184 7868 29448 7878
rect 29240 7812 29288 7868
rect 29344 7812 29392 7868
rect 29184 7802 29448 7812
rect 29036 7588 29092 7598
rect 29036 7494 29092 7532
rect 28868 7418 28924 7430
rect 28868 7366 28870 7418
rect 28922 7366 28924 7418
rect 28868 6804 28924 7366
rect 29484 6916 29540 6926
rect 28868 6748 29092 6804
rect 29036 6132 29092 6748
rect 29484 6690 29540 6860
rect 29484 6638 29486 6690
rect 29538 6638 29540 6690
rect 29484 6626 29540 6638
rect 29652 6692 29708 6702
rect 29652 6690 29764 6692
rect 29652 6638 29654 6690
rect 29706 6638 29764 6690
rect 29652 6626 29764 6638
rect 29596 6468 29652 6478
rect 29184 6300 29448 6310
rect 29240 6244 29288 6300
rect 29344 6244 29392 6300
rect 29184 6234 29448 6244
rect 29036 6076 29522 6132
rect 28700 6066 28756 6076
rect 28868 6020 28924 6030
rect 28868 5962 28924 5964
rect 28868 5910 28870 5962
rect 28922 5910 28924 5962
rect 29466 6018 29522 6076
rect 29466 5966 29468 6018
rect 29520 5966 29522 6018
rect 29466 5954 29522 5966
rect 28588 5852 28756 5908
rect 28868 5898 28924 5910
rect 29036 5906 29092 5918
rect 28364 5236 28420 5852
rect 28700 5796 28756 5852
rect 29036 5854 29038 5906
rect 29090 5854 29092 5906
rect 29036 5796 29092 5854
rect 28700 5740 29092 5796
rect 28364 5170 28420 5180
rect 27916 5058 27972 5068
rect 29184 4732 29448 4742
rect 29240 4676 29288 4732
rect 29344 4676 29392 4732
rect 29184 4666 29448 4676
rect 29596 4450 29652 6412
rect 29708 6356 29764 6626
rect 29820 6580 29876 7980
rect 29820 6514 29876 6524
rect 29708 6290 29764 6300
rect 29932 6356 29988 9884
rect 30380 9604 30436 9614
rect 30380 9156 30436 9548
rect 30380 9062 30436 9100
rect 30212 9044 30268 9054
rect 30212 8950 30268 8988
rect 30716 9044 30772 9054
rect 30716 8950 30772 8988
rect 30940 8260 30996 10220
rect 31164 9938 31220 11116
rect 31164 9886 31166 9938
rect 31218 9886 31220 9938
rect 31164 9874 31220 9886
rect 31500 9156 31556 12236
rect 31500 9090 31556 9100
rect 31612 9044 31668 12684
rect 32060 12302 32116 13244
rect 32060 12290 32134 12302
rect 32060 12238 32080 12290
rect 32132 12238 32134 12290
rect 32060 12236 32134 12238
rect 32078 12226 32134 12236
rect 32620 12292 32676 14450
rect 33628 14642 33684 15036
rect 34020 15092 34076 15206
rect 34020 15026 34076 15036
rect 33846 14924 34110 14934
rect 33902 14868 33950 14924
rect 34006 14868 34054 14924
rect 33846 14858 34110 14868
rect 33628 14590 33630 14642
rect 33682 14590 33684 14642
rect 33068 13748 33124 13758
rect 33068 13654 33124 13692
rect 33628 13748 33684 14590
rect 33180 13076 33236 13086
rect 32620 12226 32676 12236
rect 32732 12964 32788 12974
rect 32732 12850 32788 12908
rect 33180 12962 33236 13020
rect 33180 12910 33182 12962
rect 33234 12910 33236 12962
rect 33180 12898 33236 12910
rect 33348 12906 33404 12918
rect 32732 12798 32734 12850
rect 32786 12798 32788 12850
rect 31836 12180 31892 12190
rect 31836 12086 31892 12124
rect 32732 12180 32788 12798
rect 33348 12854 33350 12906
rect 33402 12854 33404 12906
rect 33348 12404 33404 12854
rect 33348 12348 33572 12404
rect 32732 12114 32788 12124
rect 31948 9826 32004 9838
rect 31948 9774 31950 9826
rect 32002 9774 32004 9826
rect 31948 9604 32004 9774
rect 32620 9828 32676 9838
rect 32620 9734 32676 9772
rect 32844 9828 32900 9838
rect 32844 9734 32900 9772
rect 33124 9828 33180 9838
rect 33404 9828 33460 9838
rect 33124 9826 33460 9828
rect 33124 9774 33126 9826
rect 33178 9774 33406 9826
rect 33458 9774 33460 9826
rect 33124 9772 33460 9774
rect 33124 9762 33180 9772
rect 33404 9762 33460 9772
rect 31948 9538 32004 9548
rect 32340 9604 32396 9614
rect 32340 9510 32396 9548
rect 32956 9604 33012 9614
rect 31612 8978 31668 8988
rect 32060 9044 32116 9054
rect 30604 8034 30660 8046
rect 30604 7982 30606 8034
rect 30658 7982 30660 8034
rect 30268 7588 30324 7598
rect 29932 6290 29988 6300
rect 30044 6916 30100 6926
rect 30044 6074 30100 6860
rect 30156 6692 30212 6702
rect 30156 6598 30212 6636
rect 30268 6356 30324 7532
rect 30604 7588 30660 7982
rect 30604 7522 30660 7532
rect 30940 7474 30996 8204
rect 32060 8258 32116 8988
rect 32172 8820 32228 8830
rect 32172 8726 32228 8764
rect 32060 8206 32062 8258
rect 32114 8206 32116 8258
rect 32060 8194 32116 8206
rect 32172 8260 32228 8270
rect 32172 8166 32228 8204
rect 30940 7422 30942 7474
rect 30994 7422 30996 7474
rect 30940 7410 30996 7422
rect 32508 8034 32564 8046
rect 32508 7982 32510 8034
rect 32562 7982 32564 8034
rect 32508 7476 32564 7982
rect 32508 7410 32564 7420
rect 30604 7250 30660 7262
rect 30604 7198 30606 7250
rect 30658 7198 30660 7250
rect 30604 6916 30660 7198
rect 30604 6850 30660 6860
rect 30716 6690 30772 6702
rect 30716 6638 30718 6690
rect 30770 6638 30772 6690
rect 30398 6580 30454 6590
rect 30716 6580 30772 6638
rect 30940 6692 30996 6702
rect 30940 6690 31108 6692
rect 30940 6638 30942 6690
rect 30994 6638 31108 6690
rect 30940 6636 31108 6638
rect 30940 6626 30996 6636
rect 30398 6578 30660 6580
rect 30398 6526 30400 6578
rect 30452 6526 30660 6578
rect 30398 6524 30660 6526
rect 30398 6514 30454 6524
rect 30268 6300 30548 6356
rect 30044 6022 30046 6074
rect 30098 6022 30100 6074
rect 30044 6010 30100 6022
rect 30212 6132 30268 6142
rect 30212 5962 30268 6076
rect 30492 6020 30548 6300
rect 30604 6244 30660 6524
rect 30716 6514 30772 6524
rect 30604 6188 30940 6244
rect 30716 6020 30772 6030
rect 30492 6018 30772 6020
rect 30492 5966 30718 6018
rect 30770 5966 30772 6018
rect 30492 5964 30772 5966
rect 29708 5908 29764 5918
rect 30212 5910 30214 5962
rect 30266 5910 30268 5962
rect 30716 5954 30772 5964
rect 30884 5962 30940 6188
rect 31052 6132 31108 6636
rect 31220 6580 31276 6590
rect 31948 6580 32004 6590
rect 31220 6578 31892 6580
rect 31220 6526 31222 6578
rect 31274 6526 31892 6578
rect 31220 6524 31892 6526
rect 31220 6514 31276 6524
rect 31052 6076 31686 6132
rect 30212 5908 30268 5910
rect 29708 5814 29764 5852
rect 30156 5852 30268 5908
rect 30884 5910 30886 5962
rect 30938 5910 30940 5962
rect 31630 6018 31686 6076
rect 31630 5966 31632 6018
rect 31684 5966 31686 6018
rect 31630 5954 31686 5966
rect 30884 5898 30940 5910
rect 31388 5906 31444 5918
rect 31388 5854 31390 5906
rect 31442 5854 31444 5906
rect 29596 4398 29598 4450
rect 29650 4398 29652 4450
rect 29596 4386 29652 4398
rect 29932 5122 29988 5134
rect 29932 5070 29934 5122
rect 29986 5070 29988 5122
rect 27692 4338 27860 4340
rect 27692 4286 27694 4338
rect 27746 4286 27860 4338
rect 27692 4284 27860 4286
rect 29932 4340 29988 5070
rect 27692 4274 27748 4284
rect 29932 4274 29988 4284
rect 28476 3780 28532 3790
rect 27580 3778 28532 3780
rect 27580 3726 28478 3778
rect 28530 3726 28532 3778
rect 27580 3724 28532 3726
rect 24556 3526 24612 3724
rect 27468 3714 27524 3724
rect 28476 3714 28532 3724
rect 30156 3778 30212 5852
rect 31388 5460 31444 5854
rect 31388 5394 31444 5404
rect 30716 5122 30772 5134
rect 30716 5070 30718 5122
rect 30770 5070 30772 5122
rect 30716 4562 30772 5070
rect 30716 4510 30718 4562
rect 30770 4510 30772 4562
rect 30716 4498 30772 4510
rect 31836 4338 31892 6524
rect 31948 5906 32004 6524
rect 31948 5854 31950 5906
rect 32002 5854 32004 5906
rect 31948 5842 32004 5854
rect 32172 6580 32228 6590
rect 32172 5906 32228 6524
rect 32172 5854 32174 5906
rect 32226 5854 32228 5906
rect 32172 5842 32228 5854
rect 32284 6356 32340 6366
rect 31836 4286 31838 4338
rect 31890 4286 31892 4338
rect 31836 4274 31892 4286
rect 30156 3726 30158 3778
rect 30210 3726 30212 3778
rect 30156 3714 30212 3726
rect 32284 3780 32340 6300
rect 32452 5684 32508 5694
rect 32452 5682 32900 5684
rect 32452 5630 32454 5682
rect 32506 5630 32900 5682
rect 32452 5628 32900 5630
rect 32452 5618 32508 5628
rect 32620 5460 32676 5470
rect 32620 5234 32676 5404
rect 32620 5182 32622 5234
rect 32674 5182 32676 5234
rect 32620 5170 32676 5182
rect 32844 4340 32900 5628
rect 32956 5122 33012 9548
rect 33516 9380 33572 12348
rect 33628 10612 33684 13692
rect 33852 14420 33908 14430
rect 33852 13746 33908 14364
rect 34300 14420 34356 15820
rect 34300 14354 34356 14364
rect 34412 13972 34468 16044
rect 34524 16034 34580 16044
rect 35308 16100 35364 16110
rect 35532 16100 35588 17276
rect 35308 16098 35588 16100
rect 35308 16046 35310 16098
rect 35362 16046 35588 16098
rect 36204 16268 36540 16324
rect 35308 16044 35588 16046
rect 35308 16034 35364 16044
rect 35812 16042 35868 16054
rect 35812 15990 35814 16042
rect 35866 15990 35868 16042
rect 35812 15764 35868 15990
rect 35980 15986 36036 15998
rect 35980 15934 35982 15986
rect 36034 15934 36036 15986
rect 35980 15876 36036 15934
rect 35980 15810 36036 15820
rect 35290 15708 35868 15764
rect 35290 15426 35346 15708
rect 36204 15652 36260 16268
rect 36484 16212 36540 16268
rect 36484 16118 36540 16156
rect 35290 15374 35292 15426
rect 35344 15374 35346 15426
rect 35290 15362 35346 15374
rect 35868 15596 36260 15652
rect 36316 16100 36372 16110
rect 34524 15314 34580 15326
rect 34524 15262 34526 15314
rect 34578 15262 34580 15314
rect 34524 14084 34580 15262
rect 35532 15316 35588 15326
rect 35532 15222 35588 15260
rect 35308 15204 35364 15214
rect 34766 15092 34822 15102
rect 35308 15092 35476 15148
rect 34766 15090 35028 15092
rect 34766 15038 34768 15090
rect 34820 15038 35028 15090
rect 34766 15036 35028 15038
rect 34766 15026 34822 15036
rect 34524 14018 34580 14028
rect 34412 13906 34468 13916
rect 33852 13694 33854 13746
rect 33906 13694 33908 13746
rect 33852 13682 33908 13694
rect 34300 13412 34356 13422
rect 34972 13412 35028 15036
rect 35420 14418 35476 15092
rect 35420 14366 35422 14418
rect 35474 14366 35476 14418
rect 33846 13356 34110 13366
rect 33902 13300 33950 13356
rect 34006 13300 34054 13356
rect 33846 13290 34110 13300
rect 33852 12964 33908 12974
rect 33852 12870 33908 12908
rect 34094 12852 34150 12862
rect 34094 12758 34150 12796
rect 33908 12740 33964 12750
rect 33908 12402 33964 12684
rect 33908 12350 33910 12402
rect 33962 12350 33964 12402
rect 33908 12338 33964 12350
rect 34300 12302 34356 13356
rect 34244 12290 34356 12302
rect 34244 12238 34246 12290
rect 34298 12238 34356 12290
rect 34244 12236 34356 12238
rect 34524 13356 35028 13412
rect 35308 14084 35364 14094
rect 34244 12226 34300 12236
rect 34524 12178 34580 13356
rect 34636 13188 34692 13198
rect 34636 12964 34692 13132
rect 35308 12962 35364 14028
rect 35420 13412 35476 14366
rect 35588 14474 35644 14486
rect 35588 14422 35590 14474
rect 35642 14422 35644 14474
rect 35588 14196 35644 14422
rect 35588 14130 35644 14140
rect 35756 13748 35812 13758
rect 35756 13654 35812 13692
rect 35420 13346 35476 13356
rect 34636 12870 34692 12908
rect 34804 12906 34860 12918
rect 34804 12854 34806 12906
rect 34858 12854 34860 12906
rect 35308 12910 35310 12962
rect 35362 12910 35364 12962
rect 35308 12898 35364 12910
rect 35550 12964 35606 12974
rect 35550 12870 35606 12908
rect 35868 12962 35924 15596
rect 36204 15428 36260 15438
rect 36204 15334 36260 15372
rect 36036 15258 36092 15270
rect 36036 15206 36038 15258
rect 36090 15206 36092 15258
rect 36036 15148 36092 15206
rect 35980 15092 36092 15148
rect 36204 15092 36260 15102
rect 35980 14308 36036 15092
rect 36092 14532 36148 14542
rect 36204 14532 36260 15036
rect 36316 14766 36372 16044
rect 36316 14754 36390 14766
rect 36316 14702 36336 14754
rect 36388 14702 36390 14754
rect 36316 14700 36390 14702
rect 36334 14690 36390 14700
rect 36092 14530 36260 14532
rect 36092 14478 36094 14530
rect 36146 14478 36260 14530
rect 36092 14476 36260 14478
rect 36092 14466 36148 14476
rect 35980 14252 36148 14308
rect 36092 13748 36148 14252
rect 36298 14196 36354 14206
rect 36298 13858 36354 14140
rect 36298 13806 36300 13858
rect 36352 13806 36354 13858
rect 36298 13794 36354 13806
rect 36092 13692 36260 13748
rect 35868 12910 35870 12962
rect 35922 12910 35924 12962
rect 34524 12126 34526 12178
rect 34578 12126 34580 12178
rect 34524 12114 34580 12126
rect 34636 12740 34692 12750
rect 34636 12178 34692 12684
rect 34804 12404 34860 12854
rect 35868 12852 35924 12910
rect 35868 12786 35924 12796
rect 36092 12962 36148 12974
rect 36092 12910 36094 12962
rect 36146 12910 36148 12962
rect 36092 12852 36148 12910
rect 36092 12786 36148 12796
rect 34636 12126 34638 12178
rect 34690 12126 34692 12178
rect 34636 12114 34692 12126
rect 34748 12348 34860 12404
rect 35252 12740 35308 12750
rect 35252 12402 35308 12684
rect 35252 12350 35254 12402
rect 35306 12350 35308 12402
rect 33846 11788 34110 11798
rect 33902 11732 33950 11788
rect 34006 11732 34054 11788
rect 33846 11722 34110 11732
rect 34748 10724 34804 12348
rect 35252 12338 35308 12350
rect 35644 12740 35700 12750
rect 35644 12290 35700 12684
rect 35644 12238 35646 12290
rect 35698 12238 35700 12290
rect 35644 12226 35700 12238
rect 35252 11172 35308 11182
rect 34524 10668 34804 10724
rect 34972 11170 35308 11172
rect 34972 11118 35254 11170
rect 35306 11118 35308 11170
rect 34972 11116 35308 11118
rect 33964 10612 34020 10622
rect 33628 10610 34020 10612
rect 33628 10558 33966 10610
rect 34018 10558 34020 10610
rect 33628 10556 34020 10558
rect 33628 9604 33684 10556
rect 33964 10546 34020 10556
rect 33846 10220 34110 10230
rect 33902 10164 33950 10220
rect 34006 10164 34054 10220
rect 33846 10154 34110 10164
rect 33628 9538 33684 9548
rect 33516 9324 33684 9380
rect 33292 8820 33348 8830
rect 33292 6690 33348 8764
rect 33292 6638 33294 6690
rect 33346 6638 33348 6690
rect 33292 6626 33348 6638
rect 33460 6634 33516 6646
rect 33460 6582 33462 6634
rect 33514 6582 33516 6634
rect 33460 6132 33516 6582
rect 33162 6076 33516 6132
rect 33628 6468 33684 9324
rect 33846 8652 34110 8662
rect 33902 8596 33950 8652
rect 34006 8596 34054 8652
rect 33846 8586 34110 8596
rect 34412 8372 34468 8382
rect 34188 8258 34244 8270
rect 34188 8206 34190 8258
rect 34242 8206 34244 8258
rect 33846 7084 34110 7094
rect 33902 7028 33950 7084
rect 34006 7028 34054 7084
rect 33846 7018 34110 7028
rect 34188 6916 34244 8206
rect 34412 8258 34468 8316
rect 34412 8206 34414 8258
rect 34466 8206 34468 8258
rect 34412 8194 34468 8206
rect 34524 7700 34580 10668
rect 34748 10498 34804 10510
rect 34748 10446 34750 10498
rect 34802 10446 34804 10498
rect 34748 10052 34804 10446
rect 34860 10052 34916 10062
rect 34748 10050 34916 10052
rect 34748 9998 34862 10050
rect 34914 9998 34916 10050
rect 34748 9996 34916 9998
rect 34860 9986 34916 9996
rect 34972 9604 35028 11116
rect 35252 11106 35308 11116
rect 34972 9538 35028 9548
rect 35252 9604 35308 9614
rect 35252 9266 35308 9548
rect 35252 9214 35254 9266
rect 35306 9214 35308 9266
rect 35252 9202 35308 9214
rect 35980 9268 36036 9278
rect 35644 8932 35700 8942
rect 35644 8930 35812 8932
rect 35644 8878 35646 8930
rect 35698 8878 35812 8930
rect 35644 8876 35812 8878
rect 35644 8866 35700 8876
rect 35756 8260 35812 8876
rect 35980 8382 36036 9212
rect 35980 8370 36054 8382
rect 35980 8318 36000 8370
rect 36052 8318 36054 8370
rect 35980 8316 36054 8318
rect 35998 8306 36054 8316
rect 35252 8202 35308 8214
rect 34692 8148 34748 8158
rect 34692 8054 34748 8092
rect 35084 8146 35140 8158
rect 35084 8094 35086 8146
rect 35138 8094 35140 8146
rect 34524 7644 34692 7700
rect 34076 6860 34244 6916
rect 34300 7476 34356 7486
rect 33964 6692 34020 6702
rect 33964 6598 34020 6636
rect 34076 6468 34132 6860
rect 34300 6804 34356 7420
rect 34468 7418 34524 7430
rect 34468 7366 34470 7418
rect 34522 7366 34524 7418
rect 34468 7364 34524 7366
rect 34468 7298 34524 7308
rect 34636 6916 34692 7644
rect 34524 6860 34692 6916
rect 34972 7474 35028 7486
rect 34972 7422 34974 7474
rect 35026 7422 35028 7474
rect 34300 6748 34468 6804
rect 34206 6580 34262 6590
rect 34206 6486 34262 6524
rect 33628 6412 33964 6468
rect 33162 6018 33218 6076
rect 33162 5966 33164 6018
rect 33216 5966 33218 6018
rect 33162 5954 33218 5966
rect 33404 5906 33460 5918
rect 33404 5854 33406 5906
rect 33458 5854 33460 5906
rect 33404 5460 33460 5854
rect 33404 5394 33460 5404
rect 32956 5070 32958 5122
rect 33010 5070 33012 5122
rect 32956 5058 33012 5070
rect 32956 4340 33012 4350
rect 32844 4338 33012 4340
rect 32844 4286 32958 4338
rect 33010 4286 33012 4338
rect 32844 4284 33012 4286
rect 32956 4274 33012 4284
rect 32396 3780 32452 3790
rect 32284 3778 32452 3780
rect 32284 3726 32398 3778
rect 32450 3726 32452 3778
rect 32284 3724 32452 3726
rect 33628 3780 33684 6412
rect 33908 5962 33964 6412
rect 34076 6132 34132 6412
rect 34076 6076 34244 6132
rect 33908 5910 33910 5962
rect 33962 5910 33964 5962
rect 33908 5898 33964 5910
rect 34076 5906 34132 5918
rect 34076 5854 34078 5906
rect 34130 5854 34132 5906
rect 34076 5684 34132 5854
rect 34188 5908 34244 6076
rect 34188 5842 34244 5852
rect 34412 5684 34468 6748
rect 34524 6244 34580 6860
rect 34972 6804 35028 7422
rect 35084 7476 35140 8094
rect 35252 8150 35254 8202
rect 35306 8150 35308 8202
rect 35756 8166 35812 8204
rect 35252 8036 35308 8150
rect 35252 7970 35308 7980
rect 35532 8148 35588 8158
rect 35214 7700 35270 7710
rect 35214 7586 35270 7644
rect 35214 7534 35216 7586
rect 35268 7534 35270 7586
rect 35214 7522 35270 7534
rect 35084 7410 35140 7420
rect 35532 7474 35588 8092
rect 36204 8036 36260 13692
rect 36540 13746 36596 13758
rect 36540 13694 36542 13746
rect 36594 13694 36596 13746
rect 36372 13524 36428 13534
rect 36372 13186 36428 13468
rect 36372 13134 36374 13186
rect 36426 13134 36428 13186
rect 36372 13122 36428 13134
rect 36540 12740 36596 13694
rect 36540 12674 36596 12684
rect 36652 12404 36708 17724
rect 37100 17778 37212 17780
rect 37100 17726 37158 17778
rect 37210 17726 37212 17778
rect 37100 17714 37212 17726
rect 36988 16772 37044 16782
rect 36876 16212 36932 16222
rect 36876 16098 36932 16156
rect 36876 16046 36878 16098
rect 36930 16046 36932 16098
rect 36876 16034 36932 16046
rect 36876 15428 36932 15438
rect 36876 13300 36932 15372
rect 36988 15316 37044 16716
rect 37100 16548 37156 17714
rect 37212 16772 37268 16782
rect 37212 16678 37268 16716
rect 37324 16660 37380 21084
rect 37436 20020 37492 21310
rect 37660 21140 37716 21150
rect 37660 20802 37716 21084
rect 37902 21028 37958 21038
rect 38108 21028 38164 27132
rect 38220 24836 38276 27580
rect 38332 27076 38388 27806
rect 38332 25844 38388 27020
rect 38508 26684 38772 26694
rect 38564 26628 38612 26684
rect 38668 26628 38716 26684
rect 38508 26618 38772 26628
rect 38332 25778 38388 25788
rect 38508 25116 38772 25126
rect 38564 25060 38612 25116
rect 38668 25060 38716 25116
rect 38508 25050 38772 25060
rect 38220 24770 38276 24780
rect 38276 24612 38332 24622
rect 38276 24164 38332 24556
rect 38276 24098 38332 24108
rect 38508 23548 38772 23558
rect 38564 23492 38612 23548
rect 38668 23492 38716 23548
rect 38508 23482 38772 23492
rect 38332 23154 38388 23166
rect 38332 23102 38334 23154
rect 38386 23102 38388 23154
rect 38332 22932 38388 23102
rect 38332 22494 38388 22876
rect 38276 22482 38388 22494
rect 38276 22430 38278 22482
rect 38330 22430 38388 22482
rect 38276 22428 38388 22430
rect 38276 22418 38332 22428
rect 38508 21980 38772 21990
rect 38564 21924 38612 21980
rect 38668 21924 38716 21980
rect 38508 21914 38772 21924
rect 37902 21026 38164 21028
rect 37902 20974 37904 21026
rect 37956 20974 38164 21026
rect 37902 20972 38164 20974
rect 37902 20962 37958 20972
rect 38892 20916 38948 29148
rect 39004 24612 39060 33852
rect 39004 24546 39060 24556
rect 38892 20850 38948 20860
rect 37660 20750 37662 20802
rect 37714 20750 37716 20802
rect 37660 20738 37716 20750
rect 37996 20804 38052 20814
rect 37548 20020 37604 20030
rect 37436 20018 37604 20020
rect 37436 19966 37550 20018
rect 37602 19966 37604 20018
rect 37436 19964 37604 19966
rect 37548 19954 37604 19964
rect 37996 19458 38052 20748
rect 38508 20412 38772 20422
rect 38564 20356 38612 20412
rect 38668 20356 38716 20412
rect 38508 20346 38772 20356
rect 37996 19406 37998 19458
rect 38050 19406 38052 19458
rect 37996 19394 38052 19406
rect 38332 20018 38388 20030
rect 38332 19966 38334 20018
rect 38386 19966 38388 20018
rect 38332 19460 38388 19966
rect 38332 19394 38388 19404
rect 38444 20020 38500 20030
rect 37604 19236 37660 19246
rect 37604 19142 37660 19180
rect 38332 19236 38388 19246
rect 38444 19236 38500 19964
rect 38388 19180 38500 19236
rect 38332 19142 38388 19180
rect 38508 18844 38772 18854
rect 38564 18788 38612 18844
rect 38668 18788 38716 18844
rect 38508 18778 38772 18788
rect 38332 17666 38388 17678
rect 38332 17614 38334 17666
rect 38386 17614 38388 17666
rect 37604 17442 37660 17454
rect 37604 17390 37606 17442
rect 37658 17390 37660 17442
rect 37604 17108 37660 17390
rect 37996 17442 38052 17454
rect 37996 17390 37998 17442
rect 38050 17390 38052 17442
rect 37996 17220 38052 17390
rect 37996 17154 38052 17164
rect 37604 17042 37660 17052
rect 38332 17108 38388 17614
rect 38508 17276 38772 17286
rect 38564 17220 38612 17276
rect 38668 17220 38716 17276
rect 38508 17210 38772 17220
rect 38332 17042 38388 17052
rect 37324 16594 37380 16604
rect 37100 16492 37268 16548
rect 37100 16100 37156 16110
rect 37100 16006 37156 16044
rect 36988 15250 37044 15260
rect 37212 14654 37268 16492
rect 37380 16324 37436 16334
rect 37380 16230 37436 16268
rect 38508 15708 38772 15718
rect 38564 15652 38612 15708
rect 38668 15652 38716 15708
rect 38508 15642 38772 15652
rect 37156 14644 37268 14654
rect 37156 14642 38276 14644
rect 37156 14590 37158 14642
rect 37210 14590 38276 14642
rect 37156 14588 38276 14590
rect 37156 14578 37212 14588
rect 37996 14420 38052 14430
rect 37996 14326 38052 14364
rect 37604 14308 37660 14318
rect 37604 14214 37660 14252
rect 37044 13916 37380 13972
rect 37044 13802 37100 13916
rect 37044 13750 37046 13802
rect 37098 13750 37100 13802
rect 37044 13738 37100 13750
rect 37212 13746 37268 13758
rect 37212 13694 37214 13746
rect 37266 13694 37268 13746
rect 36876 13234 36932 13244
rect 36988 13412 37044 13422
rect 36988 12962 37044 13356
rect 37212 13412 37268 13694
rect 37212 13346 37268 13356
rect 37324 13300 37380 13916
rect 37436 13746 37492 13758
rect 37436 13694 37438 13746
rect 37490 13694 37492 13746
rect 37436 13524 37492 13694
rect 37772 13524 37828 13534
rect 37436 13458 37492 13468
rect 37548 13522 37828 13524
rect 37548 13470 37774 13522
rect 37826 13470 37828 13522
rect 37548 13468 37828 13470
rect 37324 13244 37492 13300
rect 36988 12910 36990 12962
rect 37042 12910 37044 12962
rect 36988 12898 37044 12910
rect 37156 12964 37212 12974
rect 37156 12870 37212 12908
rect 36428 12348 36708 12404
rect 36428 11620 36484 12348
rect 36428 11564 36708 11620
rect 36652 10724 36708 11564
rect 37268 10836 37324 10846
rect 37268 10742 37324 10780
rect 36652 10630 36708 10668
rect 37156 9770 37212 9782
rect 37156 9718 37158 9770
rect 37210 9718 37212 9770
rect 37156 9268 37212 9718
rect 37156 9202 37212 9212
rect 37324 9658 37380 9670
rect 37324 9606 37326 9658
rect 37378 9606 37380 9658
rect 37324 8820 37380 9606
rect 37324 8754 37380 8764
rect 36988 8708 37044 8718
rect 36204 7970 36260 7980
rect 36652 8484 36708 8494
rect 36652 7698 36708 8428
rect 36652 7646 36654 7698
rect 36706 7646 36708 7698
rect 36652 7634 36708 7646
rect 36988 8146 37044 8652
rect 36988 8094 36990 8146
rect 37042 8094 37044 8146
rect 35532 7422 35534 7474
rect 35586 7422 35588 7474
rect 35532 7410 35588 7422
rect 34972 6748 35252 6804
rect 34636 6692 34692 6702
rect 34636 6690 35140 6692
rect 34636 6638 34638 6690
rect 34690 6638 35140 6690
rect 34636 6636 35140 6638
rect 34636 6626 34692 6636
rect 34524 6188 35028 6244
rect 34860 6020 34916 6030
rect 34636 5908 34692 5918
rect 34636 5814 34692 5852
rect 34860 5906 34916 5964
rect 34860 5854 34862 5906
rect 34914 5854 34916 5906
rect 34860 5842 34916 5854
rect 34972 5796 35028 6188
rect 35084 6030 35140 6636
rect 35196 6580 35252 6748
rect 35196 6514 35252 6524
rect 35644 6692 35700 6702
rect 35084 6018 35196 6030
rect 35084 5966 35142 6018
rect 35194 5966 35196 6018
rect 35084 5964 35196 5966
rect 35140 5954 35196 5964
rect 35420 5906 35476 5918
rect 35420 5854 35422 5906
rect 35474 5854 35476 5906
rect 34972 5740 35252 5796
rect 34076 5628 35140 5684
rect 33846 5516 34110 5526
rect 33902 5460 33950 5516
rect 34006 5460 34054 5516
rect 33846 5450 34110 5460
rect 33740 5122 33796 5134
rect 33740 5070 33742 5122
rect 33794 5070 33796 5122
rect 33740 4564 33796 5070
rect 34076 4564 34132 4574
rect 33740 4562 34132 4564
rect 33740 4510 34078 4562
rect 34130 4510 34132 4562
rect 33740 4508 34132 4510
rect 34076 4498 34132 4508
rect 35084 4450 35140 5628
rect 35196 4900 35252 5740
rect 35420 5236 35476 5854
rect 35420 5170 35476 5180
rect 35644 5234 35700 6636
rect 36988 6690 37044 8094
rect 37156 8202 37212 8214
rect 37156 8150 37158 8202
rect 37210 8150 37212 8202
rect 37156 7700 37212 8150
rect 37156 7634 37212 7644
rect 37324 8036 37380 8046
rect 36988 6638 36990 6690
rect 37042 6638 37044 6690
rect 36988 6626 37044 6638
rect 37156 6634 37212 6646
rect 37156 6582 37158 6634
rect 37210 6582 37212 6634
rect 36092 6466 36148 6478
rect 36092 6414 36094 6466
rect 36146 6414 36148 6466
rect 35644 5182 35646 5234
rect 35698 5182 35700 5234
rect 35196 4844 35308 4900
rect 35084 4398 35086 4450
rect 35138 4398 35140 4450
rect 35084 4386 35140 4398
rect 35252 4394 35308 4844
rect 35252 4342 35254 4394
rect 35306 4342 35308 4394
rect 33846 3948 34110 3958
rect 33902 3892 33950 3948
rect 34006 3892 34054 3948
rect 33846 3882 34110 3892
rect 33852 3780 33908 3790
rect 33628 3778 33908 3780
rect 33628 3726 33854 3778
rect 33906 3726 33908 3778
rect 33628 3724 33908 3726
rect 32396 3714 32452 3724
rect 33852 3714 33908 3724
rect 35252 3780 35308 4342
rect 35644 4340 35700 5182
rect 35980 6132 36036 6142
rect 35980 4462 36036 6076
rect 36092 5908 36148 6414
rect 37156 6132 37212 6582
rect 37156 6066 37212 6076
rect 36204 5908 36260 5918
rect 36092 5906 36260 5908
rect 36092 5854 36206 5906
rect 36258 5854 36260 5906
rect 36092 5852 36260 5854
rect 36204 5842 36260 5852
rect 36260 5236 36316 5246
rect 36260 5142 36316 5180
rect 37156 5236 37212 5246
rect 37156 5142 37212 5180
rect 35980 4450 36054 4462
rect 35980 4398 36000 4450
rect 36052 4398 36054 4450
rect 35980 4396 36054 4398
rect 35998 4386 36054 4396
rect 35756 4340 35812 4350
rect 35644 4338 35812 4340
rect 35644 4286 35758 4338
rect 35810 4286 35812 4338
rect 35644 4284 35812 4286
rect 35756 4274 35812 4284
rect 35252 3714 35308 3724
rect 36204 3780 36260 3790
rect 36204 3686 36260 3724
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 24556 3474 24558 3526
rect 24610 3474 24612 3526
rect 24556 3462 24612 3474
rect 26236 3556 26292 3566
rect 24332 2828 24500 2884
rect 24220 2482 24276 2492
rect 24444 800 24500 2828
rect 26236 800 26292 3500
rect 27804 3556 27860 3566
rect 27804 3462 27860 3500
rect 28028 3556 28084 3566
rect 28028 800 28084 3500
rect 28812 3556 28868 3566
rect 28812 3462 28868 3500
rect 29652 3556 29708 3566
rect 29204 3444 29260 3482
rect 29652 3462 29708 3500
rect 29820 3556 29876 3566
rect 29204 3378 29260 3388
rect 29184 3164 29448 3174
rect 29240 3108 29288 3164
rect 29344 3108 29392 3164
rect 29184 3098 29448 3108
rect 29820 800 29876 3500
rect 30492 3556 30548 3566
rect 30492 3462 30548 3500
rect 30884 3556 30940 3566
rect 31668 3556 31724 3566
rect 30884 3462 30940 3500
rect 31612 3554 31724 3556
rect 31612 3502 31670 3554
rect 31722 3502 31724 3554
rect 31612 3490 31724 3502
rect 32060 3554 32116 3566
rect 33516 3556 33572 3566
rect 32060 3502 32062 3554
rect 32114 3502 32116 3554
rect 31612 3388 31668 3490
rect 32060 3388 32116 3502
rect 33404 3554 33572 3556
rect 33404 3502 33518 3554
rect 33570 3502 33572 3554
rect 33404 3500 33572 3502
rect 33404 3454 33460 3500
rect 33516 3490 33572 3500
rect 35868 3554 35924 3566
rect 35868 3502 35870 3554
rect 35922 3502 35924 3554
rect 31612 3332 32116 3388
rect 33348 3442 33460 3454
rect 33348 3390 33350 3442
rect 33402 3390 33460 3442
rect 33348 3332 33460 3390
rect 35476 3444 35532 3454
rect 35868 3444 35924 3502
rect 37100 3554 37156 3566
rect 37100 3502 37102 3554
rect 37154 3502 37156 3554
rect 35476 3442 35924 3444
rect 35476 3390 35478 3442
rect 35530 3390 35924 3442
rect 35476 3388 35924 3390
rect 36932 3442 36988 3454
rect 36932 3390 36934 3442
rect 36986 3390 36988 3442
rect 36932 3388 36988 3390
rect 37100 3388 37156 3502
rect 37324 3556 37380 7980
rect 37436 7364 37492 13244
rect 37548 12178 37604 13468
rect 37772 13458 37828 13468
rect 38108 13076 38164 13086
rect 37660 12962 37716 12974
rect 37660 12910 37662 12962
rect 37714 12910 37716 12962
rect 37660 12740 37716 12910
rect 37902 12852 37958 12862
rect 37902 12758 37958 12796
rect 37660 12674 37716 12684
rect 37548 12126 37550 12178
rect 37602 12126 37604 12178
rect 37548 12114 37604 12126
rect 37996 11620 38052 11630
rect 38108 11620 38164 13020
rect 37996 11618 38164 11620
rect 37996 11566 37998 11618
rect 38050 11566 38164 11618
rect 37996 11564 38164 11566
rect 38220 12180 38276 14588
rect 38332 14530 38388 14542
rect 38332 14478 38334 14530
rect 38386 14478 38388 14530
rect 38332 14308 38388 14478
rect 38332 14242 38388 14252
rect 38508 14140 38772 14150
rect 38564 14084 38612 14140
rect 38668 14084 38716 14140
rect 38508 14074 38772 14084
rect 38508 12572 38772 12582
rect 38564 12516 38612 12572
rect 38668 12516 38716 12572
rect 38508 12506 38772 12516
rect 38332 12180 38388 12190
rect 38220 12178 38388 12180
rect 38220 12126 38334 12178
rect 38386 12126 38388 12178
rect 38220 12124 38388 12126
rect 37996 11554 38052 11564
rect 37604 11284 37660 11294
rect 37604 11190 37660 11228
rect 38220 10836 38276 12124
rect 38332 12114 38388 12124
rect 38332 11394 38388 11406
rect 38332 11342 38334 11394
rect 38386 11342 38388 11394
rect 38332 11284 38388 11342
rect 38332 11218 38388 11228
rect 38508 11004 38772 11014
rect 38564 10948 38612 11004
rect 38668 10948 38716 11004
rect 38508 10938 38772 10948
rect 37660 10724 37716 10734
rect 37660 9826 37716 10668
rect 37660 9774 37662 9826
rect 37714 9774 37716 9826
rect 37660 9762 37716 9774
rect 37902 9828 37958 9838
rect 37902 9734 37958 9772
rect 38108 9156 38164 9166
rect 37548 8930 37604 8942
rect 37548 8878 37550 8930
rect 37602 8878 37604 8930
rect 37548 8484 37604 8878
rect 37548 8418 37604 8428
rect 37902 8372 37958 8382
rect 37902 8278 37958 8316
rect 37660 8260 37716 8270
rect 37660 8166 37716 8204
rect 37996 7700 38052 7710
rect 38108 7700 38164 9100
rect 37996 7698 38164 7700
rect 37996 7646 37998 7698
rect 38050 7646 38164 7698
rect 37996 7644 38164 7646
rect 38220 9044 38276 10780
rect 38508 9436 38772 9446
rect 38564 9380 38612 9436
rect 38668 9380 38716 9436
rect 38508 9370 38772 9380
rect 38332 9044 38388 9054
rect 38220 9042 38388 9044
rect 38220 8990 38334 9042
rect 38386 8990 38388 9042
rect 38220 8988 38388 8990
rect 37996 7634 38052 7644
rect 37436 3778 37492 7308
rect 37772 7476 37828 7486
rect 37660 6690 37716 6702
rect 37660 6638 37662 6690
rect 37714 6638 37716 6690
rect 37660 6580 37716 6638
rect 37660 6514 37716 6524
rect 37772 5124 37828 7420
rect 37902 6578 37958 6590
rect 37902 6526 37904 6578
rect 37956 6526 37958 6578
rect 37902 6020 37958 6526
rect 37902 5954 37958 5964
rect 38108 6580 38164 6590
rect 38108 6018 38164 6524
rect 38108 5966 38110 6018
rect 38162 5966 38164 6018
rect 38108 5954 38164 5966
rect 37996 5348 38052 5358
rect 37996 5254 38052 5292
rect 38220 5236 38276 8988
rect 38332 8978 38388 8988
rect 38332 8372 38388 8382
rect 38332 7476 38388 8316
rect 38508 7868 38772 7878
rect 38564 7812 38612 7868
rect 38668 7812 38716 7868
rect 38508 7802 38772 7812
rect 38332 7382 38388 7420
rect 38508 6300 38772 6310
rect 38564 6244 38612 6300
rect 38668 6244 38716 6300
rect 38508 6234 38772 6244
rect 38220 5170 38276 5180
rect 38332 5460 38388 5470
rect 37660 5068 37828 5124
rect 38332 5122 38388 5404
rect 38332 5070 38334 5122
rect 38386 5070 38388 5122
rect 37660 4910 37716 5068
rect 37604 4898 37716 4910
rect 37604 4846 37606 4898
rect 37658 4846 37716 4898
rect 37604 4844 37716 4846
rect 37604 4834 37660 4844
rect 38332 4574 38388 5070
rect 38508 4732 38772 4742
rect 38564 4676 38612 4732
rect 38668 4676 38716 4732
rect 38508 4666 38772 4676
rect 38276 4562 38388 4574
rect 38276 4510 38278 4562
rect 38330 4510 38388 4562
rect 38276 4508 38388 4510
rect 38276 4498 38332 4508
rect 37828 4228 37884 4238
rect 37828 4226 38388 4228
rect 37828 4174 37830 4226
rect 37882 4174 38388 4226
rect 37828 4172 38388 4174
rect 37828 4162 37884 4172
rect 37436 3726 37438 3778
rect 37490 3726 37492 3778
rect 37436 3714 37492 3726
rect 37996 3556 38052 3566
rect 37324 3554 38052 3556
rect 37324 3502 37998 3554
rect 38050 3502 38052 3554
rect 37324 3500 38052 3502
rect 37996 3490 38052 3500
rect 38332 3554 38388 4172
rect 38332 3502 38334 3554
rect 38386 3502 38388 3554
rect 31612 3276 31780 3332
rect 31612 800 31668 3276
rect 33404 800 33460 3332
rect 35196 3332 35532 3388
rect 36932 3332 37156 3388
rect 35196 800 35252 3332
rect 36988 800 37044 3332
rect 38332 2660 38388 3502
rect 38508 3164 38772 3174
rect 38564 3108 38612 3164
rect 38668 3108 38716 3164
rect 38508 3098 38772 3108
rect 38332 2604 38836 2660
rect 38780 800 38836 2604
rect 1120 0 1232 800
rect 2912 0 3024 800
rect 4704 0 4816 800
rect 6496 0 6608 800
rect 8288 0 8400 800
rect 10080 0 10192 800
rect 11872 0 11984 800
rect 13664 0 13776 800
rect 15456 0 15568 800
rect 17248 0 17360 800
rect 19040 0 19152 800
rect 20832 0 20944 800
rect 22624 0 22736 800
rect 24416 0 24528 800
rect 26208 0 26320 800
rect 28000 0 28112 800
rect 29792 0 29904 800
rect 31584 0 31696 800
rect 33376 0 33488 800
rect 35168 0 35280 800
rect 36960 0 37072 800
rect 38752 0 38864 800
<< via2 >>
rect 5874 36874 5930 36876
rect 5874 36822 5876 36874
rect 5876 36822 5928 36874
rect 5928 36822 5930 36874
rect 5874 36820 5930 36822
rect 5978 36874 6034 36876
rect 5978 36822 5980 36874
rect 5980 36822 6032 36874
rect 6032 36822 6034 36874
rect 5978 36820 6034 36822
rect 6082 36874 6138 36876
rect 6082 36822 6084 36874
rect 6084 36822 6136 36874
rect 6136 36822 6138 36874
rect 6082 36820 6138 36822
rect 8876 36204 8932 36260
rect 5516 35644 5572 35700
rect 5180 35420 5236 35476
rect 2492 31836 2548 31892
rect 1988 31052 2044 31108
rect 5796 35698 5852 35700
rect 5796 35646 5798 35698
rect 5798 35646 5850 35698
rect 5850 35646 5852 35698
rect 5796 35644 5852 35646
rect 6188 35698 6244 35700
rect 6188 35646 6190 35698
rect 6190 35646 6242 35698
rect 6242 35646 6244 35698
rect 6188 35644 6244 35646
rect 6972 35586 7028 35588
rect 6972 35534 6974 35586
rect 6974 35534 7026 35586
rect 7026 35534 7028 35586
rect 6972 35532 7028 35534
rect 8764 35532 8820 35588
rect 5874 35306 5930 35308
rect 5874 35254 5876 35306
rect 5876 35254 5928 35306
rect 5928 35254 5930 35306
rect 5874 35252 5930 35254
rect 5978 35306 6034 35308
rect 5978 35254 5980 35306
rect 5980 35254 6032 35306
rect 6032 35254 6034 35306
rect 5978 35252 6034 35254
rect 6082 35306 6138 35308
rect 6082 35254 6084 35306
rect 6084 35254 6136 35306
rect 6136 35254 6138 35306
rect 6082 35252 6138 35254
rect 7532 35308 7588 35364
rect 5874 33738 5930 33740
rect 5874 33686 5876 33738
rect 5876 33686 5928 33738
rect 5928 33686 5930 33738
rect 5874 33684 5930 33686
rect 5978 33738 6034 33740
rect 5978 33686 5980 33738
rect 5980 33686 6032 33738
rect 6032 33686 6034 33738
rect 5978 33684 6034 33686
rect 6082 33738 6138 33740
rect 6082 33686 6084 33738
rect 6084 33686 6136 33738
rect 6136 33686 6138 33738
rect 6082 33684 6138 33686
rect 9548 35644 9604 35700
rect 10108 35196 10164 35252
rect 8204 34802 8260 34804
rect 8204 34750 8206 34802
rect 8206 34750 8258 34802
rect 8258 34750 8260 34802
rect 8204 34748 8260 34750
rect 8596 34130 8652 34132
rect 8596 34078 8598 34130
rect 8598 34078 8650 34130
rect 8650 34078 8652 34130
rect 8596 34076 8652 34078
rect 7532 33180 7588 33236
rect 4284 31948 4340 32004
rect 5180 31836 5236 31892
rect 5404 31836 5460 31892
rect 4284 31388 4340 31444
rect 4620 31778 4676 31780
rect 4620 31726 4622 31778
rect 4622 31726 4674 31778
rect 4674 31726 4676 31778
rect 4620 31724 4676 31726
rect 5068 31724 5124 31780
rect 3052 30994 3108 30996
rect 3052 30942 3054 30994
rect 3054 30942 3106 30994
rect 3106 30942 3108 30994
rect 3052 30940 3108 30942
rect 2734 30882 2790 30884
rect 2734 30830 2736 30882
rect 2736 30830 2788 30882
rect 2788 30830 2790 30882
rect 2734 30828 2790 30830
rect 2044 30268 2100 30324
rect 1876 30210 1932 30212
rect 1876 30158 1878 30210
rect 1878 30158 1930 30210
rect 1930 30158 1932 30210
rect 1876 30156 1932 30158
rect 1708 26236 1764 26292
rect 2380 30268 2436 30324
rect 2622 30268 2678 30324
rect 4060 30268 4116 30324
rect 5068 31164 5124 31220
rect 2044 25228 2100 25284
rect 3052 29148 3108 29204
rect 3612 29202 3668 29204
rect 3612 29150 3614 29202
rect 3614 29150 3666 29202
rect 3666 29150 3668 29202
rect 3612 29148 3668 29150
rect 3276 27858 3332 27860
rect 3276 27806 3278 27858
rect 3278 27806 3330 27858
rect 3330 27806 3332 27858
rect 3276 27804 3332 27806
rect 3612 27580 3668 27636
rect 3108 26348 3164 26404
rect 2940 26290 2996 26292
rect 2940 26238 2942 26290
rect 2942 26238 2994 26290
rect 2994 26238 2996 26290
rect 4228 27580 4284 27636
rect 7196 32396 7252 32452
rect 7364 32508 7420 32564
rect 5874 32170 5930 32172
rect 5874 32118 5876 32170
rect 5876 32118 5928 32170
rect 5928 32118 5930 32170
rect 5874 32116 5930 32118
rect 5978 32170 6034 32172
rect 5978 32118 5980 32170
rect 5980 32118 6032 32170
rect 6032 32118 6034 32170
rect 5978 32116 6034 32118
rect 6082 32170 6138 32172
rect 6082 32118 6084 32170
rect 6084 32118 6136 32170
rect 6136 32118 6138 32170
rect 6082 32116 6138 32118
rect 7084 31666 7140 31668
rect 7084 31614 7086 31666
rect 7086 31614 7138 31666
rect 7138 31614 7140 31666
rect 7084 31612 7140 31614
rect 6580 31388 6636 31444
rect 6300 31164 6356 31220
rect 5740 31106 5796 31108
rect 5740 31054 5742 31106
rect 5742 31054 5794 31106
rect 5794 31054 5796 31106
rect 5740 31052 5796 31054
rect 5628 30940 5684 30996
rect 6076 30828 6132 30884
rect 5874 30602 5930 30604
rect 5874 30550 5876 30602
rect 5876 30550 5928 30602
rect 5928 30550 5930 30602
rect 5874 30548 5930 30550
rect 5978 30602 6034 30604
rect 5978 30550 5980 30602
rect 5980 30550 6032 30602
rect 6032 30550 6034 30602
rect 5978 30548 6034 30550
rect 6082 30602 6138 30604
rect 6082 30550 6084 30602
rect 6084 30550 6136 30602
rect 6136 30550 6138 30602
rect 6082 30548 6138 30550
rect 4844 27804 4900 27860
rect 2940 26236 2996 26238
rect 2268 25228 2324 25284
rect 4060 26236 4116 26292
rect 3612 25004 3668 25060
rect 3836 24892 3892 24948
rect 3948 24780 4004 24836
rect 4956 29426 5012 29428
rect 4956 29374 4958 29426
rect 4958 29374 5010 29426
rect 5010 29374 5012 29426
rect 4956 29372 5012 29374
rect 4956 26348 5012 26404
rect 6748 30156 6804 30212
rect 5874 29034 5930 29036
rect 5874 28982 5876 29034
rect 5876 28982 5928 29034
rect 5928 28982 5930 29034
rect 5874 28980 5930 28982
rect 5978 29034 6034 29036
rect 5978 28982 5980 29034
rect 5980 28982 6032 29034
rect 6032 28982 6034 29034
rect 5978 28980 6034 28982
rect 6082 29034 6138 29036
rect 6082 28982 6084 29034
rect 6084 28982 6136 29034
rect 6136 28982 6138 29034
rect 6082 28980 6138 28982
rect 6580 29036 6636 29092
rect 7308 30957 7310 30996
rect 7310 30957 7362 30996
rect 7362 30957 7364 30996
rect 7308 30940 7364 30957
rect 7756 32732 7812 32788
rect 7644 32396 7700 32452
rect 7756 31052 7812 31108
rect 7532 30210 7588 30212
rect 7532 30158 7534 30210
rect 7534 30158 7586 30210
rect 7586 30158 7588 30210
rect 7532 30156 7588 30158
rect 8428 32732 8484 32788
rect 8764 33068 8820 33124
rect 8428 32562 8484 32564
rect 8428 32510 8430 32562
rect 8430 32510 8482 32562
rect 8482 32510 8484 32562
rect 8428 32508 8484 32510
rect 8988 33740 9044 33796
rect 10536 36090 10592 36092
rect 10536 36038 10538 36090
rect 10538 36038 10590 36090
rect 10590 36038 10592 36090
rect 10536 36036 10592 36038
rect 10640 36090 10696 36092
rect 10640 36038 10642 36090
rect 10642 36038 10694 36090
rect 10694 36038 10696 36090
rect 10640 36036 10696 36038
rect 10744 36090 10800 36092
rect 10744 36038 10746 36090
rect 10746 36038 10798 36090
rect 10798 36038 10800 36090
rect 10744 36036 10800 36038
rect 12348 36482 12404 36484
rect 12348 36430 12350 36482
rect 12350 36430 12402 36482
rect 12402 36430 12404 36482
rect 12348 36428 12404 36430
rect 10948 35196 11004 35252
rect 10220 34748 10276 34804
rect 9436 34130 9492 34132
rect 9436 34078 9438 34130
rect 9438 34078 9490 34130
rect 9490 34078 9492 34130
rect 9436 34076 9492 34078
rect 9436 33740 9492 33796
rect 9436 33404 9492 33460
rect 10052 33346 10108 33348
rect 10052 33294 10054 33346
rect 10054 33294 10106 33346
rect 10106 33294 10108 33346
rect 10052 33292 10108 33294
rect 9884 32620 9940 32676
rect 8092 32284 8148 32340
rect 8204 31948 8260 32004
rect 7998 31778 8054 31780
rect 7998 31726 8000 31778
rect 8000 31726 8052 31778
rect 8052 31726 8054 31778
rect 7998 31724 8054 31726
rect 8428 31666 8484 31668
rect 8428 31614 8430 31666
rect 8430 31614 8482 31666
rect 8482 31614 8484 31666
rect 8428 31612 8484 31614
rect 9996 32508 10052 32564
rect 8932 32338 8988 32340
rect 8932 32286 8934 32338
rect 8934 32286 8986 32338
rect 8986 32286 8988 32338
rect 8932 32284 8988 32286
rect 9342 32172 9398 32228
rect 9100 31836 9156 31892
rect 10108 32060 10164 32116
rect 10052 31500 10108 31556
rect 7774 30210 7830 30212
rect 7774 30158 7776 30210
rect 7776 30158 7828 30210
rect 7828 30158 7830 30210
rect 7774 30156 7830 30158
rect 7644 30044 7700 30100
rect 7980 29596 8036 29652
rect 7308 29260 7364 29316
rect 8540 30044 8596 30100
rect 8764 30940 8820 30996
rect 9660 31276 9716 31332
rect 10536 34522 10592 34524
rect 10536 34470 10538 34522
rect 10538 34470 10590 34522
rect 10590 34470 10592 34522
rect 10536 34468 10592 34470
rect 10640 34522 10696 34524
rect 10640 34470 10642 34522
rect 10642 34470 10694 34522
rect 10694 34470 10696 34522
rect 10640 34468 10696 34470
rect 10744 34522 10800 34524
rect 10744 34470 10746 34522
rect 10746 34470 10798 34522
rect 10798 34470 10800 34522
rect 10744 34468 10800 34470
rect 11228 33516 11284 33572
rect 10444 33458 10500 33460
rect 10444 33406 10446 33458
rect 10446 33406 10498 33458
rect 10498 33406 10500 33458
rect 10444 33404 10500 33406
rect 10780 33346 10836 33348
rect 10780 33294 10782 33346
rect 10782 33294 10834 33346
rect 10834 33294 10836 33346
rect 10780 33292 10836 33294
rect 11116 33122 11172 33124
rect 11116 33070 11118 33122
rect 11118 33070 11170 33122
rect 11170 33070 11172 33122
rect 11116 33068 11172 33070
rect 10536 32954 10592 32956
rect 10536 32902 10538 32954
rect 10538 32902 10590 32954
rect 10590 32902 10592 32954
rect 10536 32900 10592 32902
rect 10640 32954 10696 32956
rect 10640 32902 10642 32954
rect 10642 32902 10694 32954
rect 10694 32902 10696 32954
rect 10640 32900 10696 32902
rect 10744 32954 10800 32956
rect 10744 32902 10746 32954
rect 10746 32902 10798 32954
rect 10798 32902 10800 32954
rect 10744 32900 10800 32902
rect 10892 32844 10948 32900
rect 10892 32620 10948 32676
rect 10332 32172 10388 32228
rect 11340 33292 11396 33348
rect 11116 32562 11172 32564
rect 11116 32510 11118 32562
rect 11118 32510 11170 32562
rect 11170 32510 11172 32562
rect 11116 32508 11172 32510
rect 11228 32396 11284 32452
rect 10668 32172 10724 32228
rect 10444 32060 10500 32116
rect 10556 31750 10612 31780
rect 10556 31724 10558 31750
rect 10558 31724 10610 31750
rect 10610 31724 10612 31750
rect 10332 31276 10388 31332
rect 10536 31386 10592 31388
rect 10536 31334 10538 31386
rect 10538 31334 10590 31386
rect 10590 31334 10592 31386
rect 10536 31332 10592 31334
rect 10640 31386 10696 31388
rect 10640 31334 10642 31386
rect 10642 31334 10694 31386
rect 10694 31334 10696 31386
rect 10640 31332 10696 31334
rect 10744 31386 10800 31388
rect 10744 31334 10746 31386
rect 10746 31334 10798 31386
rect 10798 31334 10800 31386
rect 10744 31332 10800 31334
rect 10220 30828 10276 30884
rect 8988 30182 9044 30212
rect 8988 30156 8990 30182
rect 8990 30156 9042 30182
rect 9042 30156 9044 30182
rect 8764 30044 8820 30100
rect 5874 27466 5930 27468
rect 5874 27414 5876 27466
rect 5876 27414 5928 27466
rect 5928 27414 5930 27466
rect 5874 27412 5930 27414
rect 5978 27466 6034 27468
rect 5978 27414 5980 27466
rect 5980 27414 6032 27466
rect 6032 27414 6034 27466
rect 5978 27412 6034 27414
rect 6082 27466 6138 27468
rect 6082 27414 6084 27466
rect 6084 27414 6136 27466
rect 6136 27414 6138 27466
rect 6082 27412 6138 27414
rect 7980 28812 8036 28868
rect 7644 28700 7700 28756
rect 8540 29148 8596 29204
rect 8764 28924 8820 28980
rect 8204 28588 8260 28644
rect 8652 28812 8708 28868
rect 9548 30044 9604 30100
rect 9772 30268 9828 30324
rect 9548 29596 9604 29652
rect 9772 29372 9828 29428
rect 9884 29484 9940 29540
rect 9660 29260 9716 29316
rect 10220 30044 10276 30100
rect 10536 29818 10592 29820
rect 10536 29766 10538 29818
rect 10538 29766 10590 29818
rect 10590 29766 10592 29818
rect 10536 29764 10592 29766
rect 10640 29818 10696 29820
rect 10640 29766 10642 29818
rect 10642 29766 10694 29818
rect 10694 29766 10696 29818
rect 10640 29764 10696 29766
rect 10744 29818 10800 29820
rect 10744 29766 10746 29818
rect 10746 29766 10798 29818
rect 10798 29766 10800 29818
rect 11004 29820 11060 29876
rect 10744 29764 10800 29766
rect 10780 29426 10836 29428
rect 10780 29374 10782 29426
rect 10782 29374 10834 29426
rect 10834 29374 10836 29426
rect 10780 29372 10836 29374
rect 10108 29260 10164 29316
rect 9996 29148 10052 29204
rect 10444 29202 10500 29204
rect 10444 29150 10446 29202
rect 10446 29150 10498 29202
rect 10498 29150 10500 29202
rect 10444 29148 10500 29150
rect 10892 29036 10948 29092
rect 9436 28924 9492 28980
rect 9212 28812 9268 28868
rect 5516 26236 5572 26292
rect 5874 25898 5930 25900
rect 5874 25846 5876 25898
rect 5876 25846 5928 25898
rect 5928 25846 5930 25898
rect 5874 25844 5930 25846
rect 5978 25898 6034 25900
rect 5978 25846 5980 25898
rect 5980 25846 6032 25898
rect 6032 25846 6034 25898
rect 5978 25844 6034 25846
rect 6082 25898 6138 25900
rect 6082 25846 6084 25898
rect 6084 25846 6136 25898
rect 6136 25846 6138 25898
rect 6082 25844 6138 25846
rect 6188 25564 6244 25620
rect 4340 25282 4396 25284
rect 4340 25230 4342 25282
rect 4342 25230 4394 25282
rect 4394 25230 4396 25282
rect 4340 25228 4396 25230
rect 6972 25564 7028 25620
rect 6692 25506 6748 25508
rect 6692 25454 6694 25506
rect 6694 25454 6746 25506
rect 6746 25454 6748 25506
rect 6692 25452 6748 25454
rect 7196 25452 7252 25508
rect 4956 25228 5012 25284
rect 5740 25228 5796 25284
rect 4732 25004 4788 25060
rect 5068 24892 5124 24948
rect 4956 24668 5012 24724
rect 5572 24834 5628 24836
rect 5572 24782 5574 24834
rect 5574 24782 5626 24834
rect 5626 24782 5628 24834
rect 5572 24780 5628 24782
rect 4732 23660 4788 23716
rect 2940 23324 2996 23380
rect 4284 23378 4340 23380
rect 4284 23326 4286 23378
rect 4286 23326 4338 23378
rect 4338 23326 4340 23378
rect 4284 23324 4340 23326
rect 4844 23324 4900 23380
rect 4620 22988 4676 23044
rect 2044 22092 2100 22148
rect 2044 20802 2100 20804
rect 2044 20750 2046 20802
rect 2046 20750 2098 20802
rect 2098 20750 2100 20802
rect 2044 20748 2100 20750
rect 3164 21756 3220 21812
rect 4060 21644 4116 21700
rect 4732 21474 4788 21476
rect 4732 21422 4734 21474
rect 4734 21422 4786 21474
rect 4786 21422 4788 21474
rect 4732 21420 4788 21422
rect 5012 23042 5068 23044
rect 5012 22990 5014 23042
rect 5014 22990 5066 23042
rect 5066 22990 5068 23042
rect 5012 22988 5068 22990
rect 6636 24610 6692 24612
rect 6636 24558 6638 24610
rect 6638 24558 6690 24610
rect 6690 24558 6692 24610
rect 6636 24556 6692 24558
rect 7084 24444 7140 24500
rect 5874 24330 5930 24332
rect 5874 24278 5876 24330
rect 5876 24278 5928 24330
rect 5928 24278 5930 24330
rect 5874 24276 5930 24278
rect 5978 24330 6034 24332
rect 5978 24278 5980 24330
rect 5980 24278 6032 24330
rect 6032 24278 6034 24330
rect 5978 24276 6034 24278
rect 6082 24330 6138 24332
rect 6082 24278 6084 24330
rect 6084 24278 6136 24330
rect 6136 24278 6138 24330
rect 6082 24276 6138 24278
rect 5292 23324 5348 23380
rect 5740 23660 5796 23716
rect 6244 23266 6300 23268
rect 6244 23214 6246 23266
rect 6246 23214 6298 23266
rect 6298 23214 6300 23266
rect 6244 23212 6300 23214
rect 6860 23212 6916 23268
rect 6580 23154 6636 23156
rect 6580 23102 6582 23154
rect 6582 23102 6634 23154
rect 6634 23102 6636 23154
rect 6580 23100 6636 23102
rect 8876 28614 8932 28644
rect 8876 28588 8878 28614
rect 8878 28588 8930 28614
rect 8930 28588 8932 28614
rect 9100 27132 9156 27188
rect 8876 27074 8932 27076
rect 8876 27022 8878 27074
rect 8878 27022 8930 27074
rect 8930 27022 8932 27074
rect 8876 27020 8932 27022
rect 8764 26908 8820 26964
rect 8316 25452 8372 25508
rect 7196 23154 7252 23156
rect 7196 23102 7198 23154
rect 7198 23102 7250 23154
rect 7250 23102 7252 23154
rect 7196 23100 7252 23102
rect 6076 22988 6132 23044
rect 5874 22762 5930 22764
rect 5874 22710 5876 22762
rect 5876 22710 5928 22762
rect 5928 22710 5930 22762
rect 5874 22708 5930 22710
rect 5978 22762 6034 22764
rect 5978 22710 5980 22762
rect 5980 22710 6032 22762
rect 6032 22710 6034 22762
rect 5978 22708 6034 22710
rect 6082 22762 6138 22764
rect 6082 22710 6084 22762
rect 6084 22710 6136 22762
rect 6136 22710 6138 22762
rect 6082 22708 6138 22710
rect 5796 22146 5852 22148
rect 5796 22094 5798 22146
rect 5798 22094 5850 22146
rect 5850 22094 5852 22146
rect 5796 22092 5852 22094
rect 7756 24722 7812 24724
rect 7756 24670 7758 24722
rect 7758 24670 7810 24722
rect 7810 24670 7812 24722
rect 7756 24668 7812 24670
rect 8074 24498 8130 24500
rect 8074 24446 8076 24498
rect 8076 24446 8128 24498
rect 8128 24446 8130 24498
rect 8074 24444 8130 24446
rect 8988 24556 9044 24612
rect 7980 23212 8036 23268
rect 9324 23772 9380 23828
rect 11676 32620 11732 32676
rect 11676 32284 11732 32340
rect 12236 35420 12292 35476
rect 12348 35196 12404 35252
rect 12348 34860 12404 34916
rect 13244 36428 13300 36484
rect 13916 36204 13972 36260
rect 13356 35644 13412 35700
rect 12796 35420 12852 35476
rect 12012 33516 12068 33572
rect 12460 33516 12516 33572
rect 12236 32956 12292 33012
rect 12460 33180 12516 33236
rect 12348 32620 12404 32676
rect 12908 32956 12964 33012
rect 11900 32396 11956 32452
rect 11508 31500 11564 31556
rect 11658 31164 11714 31220
rect 11228 29932 11284 29988
rect 11452 29036 11508 29092
rect 10892 28812 10948 28868
rect 9716 28588 9772 28644
rect 10444 28642 10500 28644
rect 10444 28590 10446 28642
rect 10446 28590 10498 28642
rect 10498 28590 10500 28642
rect 10444 28588 10500 28590
rect 10780 28364 10836 28420
rect 10536 28250 10592 28252
rect 10536 28198 10538 28250
rect 10538 28198 10590 28250
rect 10590 28198 10592 28250
rect 10536 28196 10592 28198
rect 10640 28250 10696 28252
rect 10640 28198 10642 28250
rect 10642 28198 10694 28250
rect 10694 28198 10696 28250
rect 10640 28196 10696 28198
rect 10744 28250 10800 28252
rect 10744 28198 10746 28250
rect 10746 28198 10798 28250
rect 10798 28198 10800 28250
rect 10744 28196 10800 28198
rect 11900 30268 11956 30324
rect 11676 29932 11732 29988
rect 11844 29708 11900 29764
rect 11676 28812 11732 28868
rect 12124 31778 12180 31780
rect 12124 31726 12126 31778
rect 12126 31726 12178 31778
rect 12178 31726 12180 31778
rect 12124 31724 12180 31726
rect 12684 31836 12740 31892
rect 12796 31612 12852 31668
rect 12684 31500 12740 31556
rect 12236 30492 12292 30548
rect 12236 30210 12292 30212
rect 12236 30158 12238 30210
rect 12238 30158 12290 30210
rect 12290 30158 12292 30210
rect 12236 30156 12292 30158
rect 12124 29932 12180 29988
rect 12404 29708 12460 29764
rect 12572 30044 12628 30100
rect 12124 29650 12180 29652
rect 12124 29598 12126 29650
rect 12126 29598 12178 29650
rect 12178 29598 12180 29650
rect 12124 29596 12180 29598
rect 12236 29484 12292 29540
rect 14252 35196 14308 35252
rect 15198 36874 15254 36876
rect 15198 36822 15200 36874
rect 15200 36822 15252 36874
rect 15252 36822 15254 36874
rect 15198 36820 15254 36822
rect 15302 36874 15358 36876
rect 15302 36822 15304 36874
rect 15304 36822 15356 36874
rect 15356 36822 15358 36874
rect 15302 36820 15358 36822
rect 15406 36874 15462 36876
rect 15406 36822 15408 36874
rect 15408 36822 15460 36874
rect 15460 36822 15462 36874
rect 15406 36820 15462 36822
rect 14364 35084 14420 35140
rect 15596 35532 15652 35588
rect 15036 35196 15092 35252
rect 15198 35306 15254 35308
rect 15198 35254 15200 35306
rect 15200 35254 15252 35306
rect 15252 35254 15254 35306
rect 15198 35252 15254 35254
rect 15302 35306 15358 35308
rect 15302 35254 15304 35306
rect 15304 35254 15356 35306
rect 15356 35254 15358 35306
rect 15302 35252 15358 35254
rect 15406 35306 15462 35308
rect 15406 35254 15408 35306
rect 15408 35254 15460 35306
rect 15460 35254 15462 35306
rect 15406 35252 15462 35254
rect 13748 34914 13804 34916
rect 13748 34862 13750 34914
rect 13750 34862 13802 34914
rect 13802 34862 13804 34914
rect 13748 34860 13804 34862
rect 15820 35420 15876 35476
rect 15708 35084 15764 35140
rect 15036 33852 15092 33908
rect 14364 33740 14420 33796
rect 15198 33738 15254 33740
rect 15198 33686 15200 33738
rect 15200 33686 15252 33738
rect 15252 33686 15254 33738
rect 15198 33684 15254 33686
rect 15302 33738 15358 33740
rect 15302 33686 15304 33738
rect 15304 33686 15356 33738
rect 15356 33686 15358 33738
rect 15302 33684 15358 33686
rect 15406 33738 15462 33740
rect 15406 33686 15408 33738
rect 15408 33686 15460 33738
rect 15460 33686 15462 33738
rect 15406 33684 15462 33686
rect 15932 34914 15988 34916
rect 15932 34862 15934 34914
rect 15934 34862 15986 34914
rect 15986 34862 15988 34914
rect 15932 34860 15988 34862
rect 15932 34636 15988 34692
rect 15932 34300 15988 34356
rect 13356 32508 13412 32564
rect 13916 33346 13972 33348
rect 13916 33294 13918 33346
rect 13918 33294 13970 33346
rect 13970 33294 13972 33346
rect 13916 33292 13972 33294
rect 14252 33346 14308 33348
rect 14252 33294 14254 33346
rect 14254 33294 14306 33346
rect 14306 33294 14308 33346
rect 14252 33292 14308 33294
rect 14028 32284 14084 32340
rect 14364 32562 14420 32564
rect 14364 32510 14366 32562
rect 14366 32510 14418 32562
rect 14418 32510 14420 32562
rect 14364 32508 14420 32510
rect 14028 31836 14084 31892
rect 13468 31500 13524 31556
rect 13580 31164 13636 31220
rect 13692 31724 13748 31780
rect 13020 31052 13076 31108
rect 12908 29820 12964 29876
rect 12684 29596 12740 29652
rect 13524 30604 13580 30660
rect 13356 30492 13412 30548
rect 13524 30156 13580 30212
rect 13804 31612 13860 31668
rect 14364 31500 14420 31556
rect 13804 31164 13860 31220
rect 13244 29820 13300 29876
rect 14476 31388 14532 31444
rect 14812 32284 14868 32340
rect 16268 35685 16270 35700
rect 16270 35685 16322 35700
rect 16322 35685 16324 35700
rect 16268 35644 16324 35685
rect 16044 32844 16100 32900
rect 15198 32170 15254 32172
rect 15198 32118 15200 32170
rect 15200 32118 15252 32170
rect 15252 32118 15254 32170
rect 15198 32116 15254 32118
rect 15302 32170 15358 32172
rect 15302 32118 15304 32170
rect 15304 32118 15356 32170
rect 15356 32118 15358 32170
rect 15302 32116 15358 32118
rect 15406 32170 15462 32172
rect 15406 32118 15408 32170
rect 15408 32118 15460 32170
rect 15460 32118 15462 32170
rect 15406 32116 15462 32118
rect 18060 35586 18116 35588
rect 18060 35534 18062 35586
rect 18062 35534 18114 35586
rect 18114 35534 18116 35586
rect 18060 35532 18116 35534
rect 16604 34748 16660 34804
rect 16940 34636 16996 34692
rect 17276 34636 17332 34692
rect 16604 34300 16660 34356
rect 16828 33516 16884 33572
rect 16044 32450 16100 32452
rect 16044 32398 16046 32450
rect 16046 32398 16098 32450
rect 16098 32398 16100 32450
rect 16044 32396 16100 32398
rect 15036 31836 15092 31892
rect 15820 31836 15876 31892
rect 14924 31724 14980 31780
rect 14700 31500 14756 31556
rect 14588 31276 14644 31332
rect 14476 31164 14532 31220
rect 14924 30970 14926 30996
rect 14926 30970 14978 30996
rect 14978 30970 14980 30996
rect 14924 30940 14980 30970
rect 14364 30604 14420 30660
rect 14196 30492 14252 30548
rect 14028 30098 14084 30100
rect 14028 30046 14030 30098
rect 14030 30046 14082 30098
rect 14082 30046 14084 30098
rect 14028 30044 14084 30046
rect 15204 31388 15260 31444
rect 15540 31052 15596 31108
rect 15708 31500 15764 31556
rect 15036 30492 15092 30548
rect 15198 30602 15254 30604
rect 15198 30550 15200 30602
rect 15200 30550 15252 30602
rect 15252 30550 15254 30602
rect 15198 30548 15254 30550
rect 15302 30602 15358 30604
rect 15302 30550 15304 30602
rect 15304 30550 15356 30602
rect 15356 30550 15358 30602
rect 15302 30548 15358 30550
rect 15406 30602 15462 30604
rect 15406 30550 15408 30602
rect 15408 30550 15460 30602
rect 15460 30550 15462 30602
rect 15406 30548 15462 30550
rect 14942 30322 14998 30324
rect 14942 30270 14944 30322
rect 14944 30270 14996 30322
rect 14996 30270 14998 30322
rect 14942 30268 14998 30270
rect 14364 29708 14420 29764
rect 12460 28812 12516 28868
rect 9828 27858 9884 27860
rect 9828 27806 9830 27858
rect 9830 27806 9882 27858
rect 9882 27806 9884 27858
rect 9828 27804 9884 27806
rect 10724 27858 10780 27860
rect 10724 27806 10726 27858
rect 10726 27806 10778 27858
rect 10778 27806 10780 27858
rect 10724 27804 10780 27806
rect 10892 27356 10948 27412
rect 9996 27132 10052 27188
rect 9716 27020 9772 27076
rect 9660 26012 9716 26068
rect 10536 26682 10592 26684
rect 10536 26630 10538 26682
rect 10538 26630 10590 26682
rect 10590 26630 10592 26682
rect 10536 26628 10592 26630
rect 10640 26682 10696 26684
rect 10640 26630 10642 26682
rect 10642 26630 10694 26682
rect 10694 26630 10696 26682
rect 10640 26628 10696 26630
rect 10744 26682 10800 26684
rect 10744 26630 10746 26682
rect 10746 26630 10798 26682
rect 10798 26630 10800 26682
rect 10744 26628 10800 26630
rect 11508 27858 11564 27860
rect 11508 27806 11510 27858
rect 11510 27806 11562 27858
rect 11562 27806 11564 27858
rect 11508 27804 11564 27806
rect 11564 27356 11620 27412
rect 10444 26348 10500 26404
rect 10164 26012 10220 26068
rect 11284 26514 11340 26516
rect 11284 26462 11286 26514
rect 11286 26462 11338 26514
rect 11338 26462 11340 26514
rect 11284 26460 11340 26462
rect 11564 26460 11620 26516
rect 11452 26348 11508 26404
rect 11004 25506 11060 25508
rect 11004 25454 11006 25506
rect 11006 25454 11058 25506
rect 11058 25454 11060 25506
rect 11004 25452 11060 25454
rect 10536 25114 10592 25116
rect 10536 25062 10538 25114
rect 10538 25062 10590 25114
rect 10590 25062 10592 25114
rect 10536 25060 10592 25062
rect 10640 25114 10696 25116
rect 10640 25062 10642 25114
rect 10642 25062 10694 25114
rect 10694 25062 10696 25114
rect 10640 25060 10696 25062
rect 10744 25114 10800 25116
rect 10744 25062 10746 25114
rect 10746 25062 10798 25114
rect 10798 25062 10800 25114
rect 10744 25060 10800 25062
rect 9436 23324 9492 23380
rect 9212 23100 9268 23156
rect 9884 23154 9940 23156
rect 9884 23102 9886 23154
rect 9886 23102 9938 23154
rect 9938 23102 9940 23154
rect 9884 23100 9940 23102
rect 8652 22988 8708 23044
rect 7980 22652 8036 22708
rect 8204 22876 8260 22932
rect 7364 22146 7420 22148
rect 7364 22094 7366 22146
rect 7366 22094 7418 22146
rect 7418 22094 7420 22146
rect 7364 22092 7420 22094
rect 5274 21756 5330 21812
rect 6188 21698 6244 21700
rect 6188 21646 6190 21698
rect 6190 21646 6242 21698
rect 6242 21646 6244 21698
rect 6188 21644 6244 21646
rect 6524 21644 6580 21700
rect 5516 21420 5572 21476
rect 8316 22092 8372 22148
rect 8372 21474 8428 21476
rect 8372 21422 8374 21474
rect 8374 21422 8426 21474
rect 8426 21422 8428 21474
rect 8372 21420 8428 21422
rect 5874 21194 5930 21196
rect 5874 21142 5876 21194
rect 5876 21142 5928 21194
rect 5928 21142 5930 21194
rect 5874 21140 5930 21142
rect 5978 21194 6034 21196
rect 5978 21142 5980 21194
rect 5980 21142 6032 21194
rect 6032 21142 6034 21194
rect 5978 21140 6034 21142
rect 6082 21194 6138 21196
rect 6082 21142 6084 21194
rect 6084 21142 6136 21194
rect 6136 21142 6138 21194
rect 6082 21140 6138 21142
rect 5516 20972 5572 21028
rect 6468 20972 6524 21028
rect 2492 20748 2548 20804
rect 2156 19964 2212 20020
rect 5964 20802 6020 20804
rect 5964 20750 5966 20802
rect 5966 20750 6018 20802
rect 6018 20750 6020 20802
rect 5964 20748 6020 20750
rect 4060 20636 4116 20692
rect 6636 20524 6692 20580
rect 6860 20972 6916 21028
rect 4172 20018 4228 20020
rect 4172 19966 4174 20018
rect 4174 19966 4226 20018
rect 4226 19966 4228 20018
rect 4172 19964 4228 19966
rect 7308 20972 7364 21028
rect 7420 20748 7476 20804
rect 7066 20690 7122 20692
rect 7066 20638 7068 20690
rect 7068 20638 7120 20690
rect 7120 20638 7122 20690
rect 7066 20636 7122 20638
rect 7196 20524 7252 20580
rect 7812 20802 7868 20804
rect 7812 20750 7814 20802
rect 7814 20750 7866 20802
rect 7866 20750 7868 20802
rect 7812 20748 7868 20750
rect 7980 20524 8036 20580
rect 7420 20300 7476 20356
rect 8428 20188 8484 20244
rect 9642 22930 9698 22932
rect 9642 22878 9644 22930
rect 9644 22878 9696 22930
rect 9696 22878 9698 22930
rect 9642 22876 9698 22878
rect 5874 19626 5930 19628
rect 5874 19574 5876 19626
rect 5876 19574 5928 19626
rect 5928 19574 5930 19626
rect 5874 19572 5930 19574
rect 5978 19626 6034 19628
rect 5978 19574 5980 19626
rect 5980 19574 6032 19626
rect 6032 19574 6034 19626
rect 5978 19572 6034 19574
rect 6082 19626 6138 19628
rect 6082 19574 6084 19626
rect 6084 19574 6136 19626
rect 6136 19574 6138 19626
rect 6082 19572 6138 19574
rect 7980 19404 8036 19460
rect 4620 19180 4676 19236
rect 5516 19234 5572 19236
rect 5516 19182 5518 19234
rect 5518 19182 5570 19234
rect 5570 19182 5572 19234
rect 5516 19180 5572 19182
rect 7980 19234 8036 19236
rect 7980 19182 7982 19234
rect 7982 19182 8034 19234
rect 8034 19182 8036 19234
rect 7980 19180 8036 19182
rect 4172 18844 4228 18900
rect 5740 18844 5796 18900
rect 7812 18844 7868 18900
rect 8876 21420 8932 21476
rect 8204 18396 8260 18452
rect 10332 23772 10388 23828
rect 10536 23546 10592 23548
rect 10536 23494 10538 23546
rect 10538 23494 10590 23546
rect 10590 23494 10592 23546
rect 10536 23492 10592 23494
rect 10640 23546 10696 23548
rect 10640 23494 10642 23546
rect 10642 23494 10694 23546
rect 10694 23494 10696 23546
rect 10640 23492 10696 23494
rect 10744 23546 10800 23548
rect 10744 23494 10746 23546
rect 10746 23494 10798 23546
rect 10798 23494 10800 23546
rect 10744 23492 10800 23494
rect 10892 23548 10948 23604
rect 10780 23212 10836 23268
rect 10388 22988 10444 23044
rect 10892 22988 10948 23044
rect 9436 20188 9492 20244
rect 9604 20076 9660 20132
rect 5874 18058 5930 18060
rect 5874 18006 5876 18058
rect 5876 18006 5928 18058
rect 5928 18006 5930 18058
rect 5874 18004 5930 18006
rect 5978 18058 6034 18060
rect 5978 18006 5980 18058
rect 5980 18006 6032 18058
rect 6032 18006 6034 18058
rect 5978 18004 6034 18006
rect 6082 18058 6138 18060
rect 6082 18006 6084 18058
rect 6084 18006 6136 18058
rect 6136 18006 6138 18058
rect 8540 18060 8596 18116
rect 6082 18004 6138 18006
rect 8540 17890 8596 17892
rect 8540 17838 8542 17890
rect 8542 17838 8594 17890
rect 8594 17838 8596 17890
rect 8540 17836 8596 17838
rect 9044 18956 9100 19012
rect 9436 18450 9492 18452
rect 9436 18398 9438 18450
rect 9438 18398 9490 18450
rect 9490 18398 9492 18450
rect 9436 18396 9492 18398
rect 9660 18450 9716 18452
rect 9660 18398 9662 18450
rect 9662 18398 9714 18450
rect 9714 18398 9716 18450
rect 9660 18396 9716 18398
rect 10220 21756 10276 21812
rect 8764 17836 8820 17892
rect 8988 18060 9044 18116
rect 5874 16490 5930 16492
rect 5874 16438 5876 16490
rect 5876 16438 5928 16490
rect 5928 16438 5930 16490
rect 5874 16436 5930 16438
rect 5978 16490 6034 16492
rect 5978 16438 5980 16490
rect 5980 16438 6032 16490
rect 6032 16438 6034 16490
rect 5978 16436 6034 16438
rect 6082 16490 6138 16492
rect 6082 16438 6084 16490
rect 6084 16438 6136 16490
rect 6136 16438 6138 16490
rect 6082 16436 6138 16438
rect 9884 17836 9940 17892
rect 8988 17052 9044 17108
rect 9716 17106 9772 17108
rect 9716 17054 9718 17106
rect 9718 17054 9770 17106
rect 9770 17054 9772 17106
rect 9716 17052 9772 17054
rect 8652 16268 8708 16324
rect 5874 14922 5930 14924
rect 5874 14870 5876 14922
rect 5876 14870 5928 14922
rect 5928 14870 5930 14922
rect 5874 14868 5930 14870
rect 5978 14922 6034 14924
rect 5978 14870 5980 14922
rect 5980 14870 6032 14922
rect 6032 14870 6034 14922
rect 5978 14868 6034 14870
rect 6082 14922 6138 14924
rect 6082 14870 6084 14922
rect 6084 14870 6136 14922
rect 6136 14870 6138 14922
rect 6082 14868 6138 14870
rect 10536 21978 10592 21980
rect 10536 21926 10538 21978
rect 10538 21926 10590 21978
rect 10590 21926 10592 21978
rect 10536 21924 10592 21926
rect 10640 21978 10696 21980
rect 10640 21926 10642 21978
rect 10642 21926 10694 21978
rect 10694 21926 10696 21978
rect 10640 21924 10696 21926
rect 10744 21978 10800 21980
rect 10744 21926 10746 21978
rect 10746 21926 10798 21978
rect 10798 21926 10800 21978
rect 10744 21924 10800 21926
rect 11900 28364 11956 28420
rect 12740 28812 12796 28868
rect 13356 29372 13412 29428
rect 13356 28140 13412 28196
rect 12124 27916 12180 27972
rect 12124 27132 12180 27188
rect 12852 27186 12908 27188
rect 12852 27134 12854 27186
rect 12854 27134 12906 27186
rect 12906 27134 12908 27186
rect 12852 27132 12908 27134
rect 13356 27132 13412 27188
rect 11788 26796 11844 26852
rect 12348 26012 12404 26068
rect 11788 25452 11844 25508
rect 12460 25506 12516 25508
rect 12460 25454 12462 25506
rect 12462 25454 12514 25506
rect 12514 25454 12516 25506
rect 12460 25452 12516 25454
rect 11788 25228 11844 25284
rect 11004 23100 11060 23156
rect 11116 23378 11172 23380
rect 11116 23326 11118 23378
rect 11118 23326 11170 23378
rect 11170 23326 11172 23378
rect 11116 23324 11172 23326
rect 13076 25228 13132 25284
rect 12236 23938 12292 23940
rect 12236 23886 12238 23938
rect 12238 23886 12290 23938
rect 12290 23886 12292 23938
rect 12236 23884 12292 23886
rect 11788 23660 11844 23716
rect 11452 23212 11508 23268
rect 11564 23324 11620 23380
rect 12012 23324 12068 23380
rect 11116 22316 11172 22372
rect 11900 22370 11956 22372
rect 11900 22318 11902 22370
rect 11902 22318 11954 22370
rect 11954 22318 11956 22370
rect 11900 22316 11956 22318
rect 10892 21756 10948 21812
rect 11564 20972 11620 21028
rect 10536 20410 10592 20412
rect 10536 20358 10538 20410
rect 10538 20358 10590 20410
rect 10590 20358 10592 20410
rect 10536 20356 10592 20358
rect 10640 20410 10696 20412
rect 10640 20358 10642 20410
rect 10642 20358 10694 20410
rect 10694 20358 10696 20410
rect 10640 20356 10696 20358
rect 10744 20410 10800 20412
rect 10744 20358 10746 20410
rect 10746 20358 10798 20410
rect 10798 20358 10800 20410
rect 10744 20356 10800 20358
rect 12236 23660 12292 23716
rect 12908 24668 12964 24724
rect 12740 24108 12796 24164
rect 13356 23324 13412 23380
rect 13636 28812 13692 28868
rect 14010 27298 14066 27300
rect 14010 27246 14012 27298
rect 14012 27246 14064 27298
rect 14064 27246 14066 27298
rect 14010 27244 14066 27246
rect 13636 27186 13692 27188
rect 13636 27134 13638 27186
rect 13638 27134 13690 27186
rect 13690 27134 13692 27186
rect 13636 27132 13692 27134
rect 13804 26908 13860 26964
rect 14140 25452 14196 25508
rect 14812 30044 14868 30100
rect 14476 27580 14532 27636
rect 14588 28140 14644 28196
rect 13636 24444 13692 24500
rect 13636 23884 13692 23940
rect 13580 23660 13636 23716
rect 14252 24444 14308 24500
rect 12236 20860 12292 20916
rect 13916 24108 13972 24164
rect 13804 21644 13860 21700
rect 13692 21084 13748 21140
rect 13562 21026 13618 21028
rect 13562 20974 13564 21026
rect 13564 20974 13616 21026
rect 13616 20974 13618 21026
rect 13562 20972 13618 20974
rect 13356 20748 13412 20804
rect 14140 23996 14196 24052
rect 15260 30380 15316 30436
rect 16716 32620 16772 32676
rect 16492 32284 16548 32340
rect 16380 31836 16436 31892
rect 17500 33180 17556 33236
rect 17836 33516 17892 33572
rect 17948 33852 18004 33908
rect 19180 36706 19236 36708
rect 19180 36654 19182 36706
rect 19182 36654 19234 36706
rect 19234 36654 19236 36706
rect 19180 36652 19236 36654
rect 19964 36652 20020 36708
rect 18620 34802 18676 34804
rect 18620 34750 18622 34802
rect 18622 34750 18674 34802
rect 18674 34750 18676 34802
rect 18620 34748 18676 34750
rect 19068 34748 19124 34804
rect 18788 34636 18844 34692
rect 19860 36090 19916 36092
rect 19860 36038 19862 36090
rect 19862 36038 19914 36090
rect 19914 36038 19916 36090
rect 19860 36036 19916 36038
rect 19964 36090 20020 36092
rect 19964 36038 19966 36090
rect 19966 36038 20018 36090
rect 20018 36038 20020 36090
rect 19964 36036 20020 36038
rect 20068 36090 20124 36092
rect 20068 36038 20070 36090
rect 20070 36038 20122 36090
rect 20122 36038 20124 36090
rect 20068 36036 20124 36038
rect 20300 35868 20356 35924
rect 19628 34914 19684 34916
rect 19628 34862 19630 34914
rect 19630 34862 19682 34914
rect 19682 34862 19684 34914
rect 19628 34860 19684 34862
rect 19180 34300 19236 34356
rect 18284 33628 18340 33684
rect 20076 34860 20132 34916
rect 20972 35868 21028 35924
rect 20860 35644 20916 35700
rect 20580 35586 20636 35588
rect 20580 35534 20582 35586
rect 20582 35534 20634 35586
rect 20634 35534 20636 35586
rect 20580 35532 20636 35534
rect 20804 35084 20860 35140
rect 19860 34522 19916 34524
rect 19860 34470 19862 34522
rect 19862 34470 19914 34522
rect 19914 34470 19916 34522
rect 19860 34468 19916 34470
rect 19964 34522 20020 34524
rect 19964 34470 19966 34522
rect 19966 34470 20018 34522
rect 20018 34470 20020 34522
rect 19964 34468 20020 34470
rect 20068 34522 20124 34524
rect 20068 34470 20070 34522
rect 20070 34470 20122 34522
rect 20122 34470 20124 34522
rect 20068 34468 20124 34470
rect 18396 33740 18452 33796
rect 18172 33068 18228 33124
rect 20412 34354 20468 34356
rect 20412 34302 20414 34354
rect 20414 34302 20466 34354
rect 20466 34302 20468 34354
rect 20412 34300 20468 34302
rect 18060 32620 18116 32676
rect 17612 32396 17668 32452
rect 17500 32060 17556 32116
rect 17836 31948 17892 32004
rect 15932 30380 15988 30436
rect 15484 30156 15540 30212
rect 15372 29820 15428 29876
rect 15596 29820 15652 29876
rect 15198 29034 15254 29036
rect 15198 28982 15200 29034
rect 15200 28982 15252 29034
rect 15252 28982 15254 29034
rect 15198 28980 15254 28982
rect 15302 29034 15358 29036
rect 15302 28982 15304 29034
rect 15304 28982 15356 29034
rect 15356 28982 15358 29034
rect 15302 28980 15358 28982
rect 15406 29034 15462 29036
rect 15406 28982 15408 29034
rect 15408 28982 15460 29034
rect 15460 28982 15462 29034
rect 15406 28980 15462 28982
rect 16286 30604 16342 30660
rect 16940 31164 16996 31220
rect 16940 30994 16996 30996
rect 16940 30942 16942 30994
rect 16942 30942 16994 30994
rect 16994 30942 16996 30994
rect 16940 30940 16996 30942
rect 16772 30380 16828 30436
rect 16604 30268 16660 30324
rect 17500 31836 17556 31892
rect 17836 31164 17892 31220
rect 16940 30156 16996 30212
rect 16156 29932 16212 29988
rect 16268 29820 16324 29876
rect 15820 28812 15876 28868
rect 15198 27466 15254 27468
rect 15198 27414 15200 27466
rect 15200 27414 15252 27466
rect 15252 27414 15254 27466
rect 15198 27412 15254 27414
rect 15302 27466 15358 27468
rect 15302 27414 15304 27466
rect 15304 27414 15356 27466
rect 15356 27414 15358 27466
rect 15302 27412 15358 27414
rect 15406 27466 15462 27468
rect 15406 27414 15408 27466
rect 15408 27414 15460 27466
rect 15460 27414 15462 27466
rect 15406 27412 15462 27414
rect 15260 27074 15316 27076
rect 15260 27022 15262 27074
rect 15262 27022 15314 27074
rect 15314 27022 15316 27074
rect 15260 27020 15316 27022
rect 15428 27074 15484 27076
rect 15428 27022 15430 27074
rect 15430 27022 15482 27074
rect 15482 27022 15484 27074
rect 15428 27020 15484 27022
rect 14924 26962 14980 26964
rect 14924 26910 14926 26962
rect 14926 26910 14978 26962
rect 14978 26910 14980 26962
rect 14924 26908 14980 26910
rect 14980 26012 15036 26068
rect 15198 25898 15254 25900
rect 15198 25846 15200 25898
rect 15200 25846 15252 25898
rect 15252 25846 15254 25898
rect 15198 25844 15254 25846
rect 15302 25898 15358 25900
rect 15302 25846 15304 25898
rect 15304 25846 15356 25898
rect 15356 25846 15358 25898
rect 15302 25844 15358 25846
rect 15406 25898 15462 25900
rect 15406 25846 15408 25898
rect 15408 25846 15460 25898
rect 15460 25846 15462 25898
rect 15406 25844 15462 25846
rect 16604 28642 16660 28644
rect 16604 28590 16606 28642
rect 16606 28590 16658 28642
rect 16658 28590 16660 28642
rect 16604 28588 16660 28590
rect 17164 28476 17220 28532
rect 16492 28364 16548 28420
rect 17052 28364 17108 28420
rect 16604 27804 16660 27860
rect 16604 27356 16660 27412
rect 15820 27020 15876 27076
rect 16174 27074 16230 27076
rect 16174 27022 16176 27074
rect 16176 27022 16228 27074
rect 16228 27022 16230 27074
rect 16174 27020 16230 27022
rect 15260 25506 15316 25508
rect 15260 25454 15262 25506
rect 15262 25454 15314 25506
rect 15314 25454 15316 25506
rect 15260 25452 15316 25454
rect 15484 24444 15540 24500
rect 15198 24330 15254 24332
rect 15198 24278 15200 24330
rect 15200 24278 15252 24330
rect 15252 24278 15254 24330
rect 15198 24276 15254 24278
rect 15302 24330 15358 24332
rect 15302 24278 15304 24330
rect 15304 24278 15356 24330
rect 15356 24278 15358 24330
rect 15302 24276 15358 24278
rect 15406 24330 15462 24332
rect 15406 24278 15408 24330
rect 15408 24278 15460 24330
rect 15460 24278 15462 24330
rect 15406 24276 15462 24278
rect 15036 24108 15092 24164
rect 14812 22988 14868 23044
rect 14028 22876 14084 22932
rect 14812 22652 14868 22708
rect 16716 27244 16772 27300
rect 15820 26348 15876 26404
rect 16828 26348 16884 26404
rect 16380 26290 16436 26292
rect 16380 26238 16382 26290
rect 16382 26238 16434 26290
rect 16434 26238 16436 26290
rect 16380 26236 16436 26238
rect 15820 25564 15876 25620
rect 15932 26124 15988 26180
rect 16380 25452 16436 25508
rect 15652 23378 15708 23380
rect 15652 23326 15654 23378
rect 15654 23326 15706 23378
rect 15706 23326 15708 23378
rect 15652 23324 15708 23326
rect 15092 22930 15148 22932
rect 15092 22878 15094 22930
rect 15094 22878 15146 22930
rect 15146 22878 15148 22930
rect 15092 22876 15148 22878
rect 15198 22762 15254 22764
rect 15198 22710 15200 22762
rect 15200 22710 15252 22762
rect 15252 22710 15254 22762
rect 15198 22708 15254 22710
rect 15302 22762 15358 22764
rect 15302 22710 15304 22762
rect 15304 22710 15356 22762
rect 15356 22710 15358 22762
rect 15302 22708 15358 22710
rect 15406 22762 15462 22764
rect 15406 22710 15408 22762
rect 15408 22710 15460 22762
rect 15460 22710 15462 22762
rect 15406 22708 15462 22710
rect 15484 22370 15540 22372
rect 15484 22318 15486 22370
rect 15486 22318 15538 22370
rect 15538 22318 15540 22370
rect 15484 22316 15540 22318
rect 13916 20748 13972 20804
rect 15932 23324 15988 23380
rect 16604 23378 16660 23380
rect 16604 23326 16606 23378
rect 16606 23326 16658 23378
rect 16658 23326 16660 23378
rect 16604 23324 16660 23326
rect 16100 23042 16156 23044
rect 16100 22990 16102 23042
rect 16102 22990 16154 23042
rect 16154 22990 16156 23042
rect 16100 22988 16156 22990
rect 14812 21868 14868 21924
rect 14476 21644 14532 21700
rect 10668 19852 10724 19908
rect 10668 19404 10724 19460
rect 12236 19852 12292 19908
rect 11900 19292 11956 19348
rect 11284 19010 11340 19012
rect 11284 18958 11286 19010
rect 11286 18958 11338 19010
rect 11338 18958 11340 19010
rect 11284 18956 11340 18958
rect 10536 18842 10592 18844
rect 10536 18790 10538 18842
rect 10538 18790 10590 18842
rect 10590 18790 10592 18842
rect 10536 18788 10592 18790
rect 10640 18842 10696 18844
rect 10640 18790 10642 18842
rect 10642 18790 10694 18842
rect 10694 18790 10696 18842
rect 10640 18788 10696 18790
rect 10744 18842 10800 18844
rect 10744 18790 10746 18842
rect 10746 18790 10798 18842
rect 10798 18790 10800 18842
rect 10744 18788 10800 18790
rect 10892 18396 10948 18452
rect 10724 17836 10780 17892
rect 11116 18450 11172 18452
rect 11116 18398 11118 18450
rect 11118 18398 11170 18450
rect 11170 18398 11172 18450
rect 11116 18396 11172 18398
rect 10536 17274 10592 17276
rect 10536 17222 10538 17274
rect 10538 17222 10590 17274
rect 10590 17222 10592 17274
rect 10536 17220 10592 17222
rect 10640 17274 10696 17276
rect 10640 17222 10642 17274
rect 10642 17222 10694 17274
rect 10694 17222 10696 17274
rect 10640 17220 10696 17222
rect 10744 17274 10800 17276
rect 10744 17222 10746 17274
rect 10746 17222 10798 17274
rect 10798 17222 10800 17274
rect 10744 17220 10800 17222
rect 11900 17724 11956 17780
rect 10332 16044 10388 16100
rect 10892 16044 10948 16100
rect 10536 15706 10592 15708
rect 10536 15654 10538 15706
rect 10538 15654 10590 15706
rect 10590 15654 10592 15706
rect 10536 15652 10592 15654
rect 10640 15706 10696 15708
rect 10640 15654 10642 15706
rect 10642 15654 10694 15706
rect 10694 15654 10696 15706
rect 10640 15652 10696 15654
rect 10744 15706 10800 15708
rect 10744 15654 10746 15706
rect 10746 15654 10798 15706
rect 10798 15654 10800 15706
rect 10744 15652 10800 15654
rect 10220 14700 10276 14756
rect 5874 13354 5930 13356
rect 5874 13302 5876 13354
rect 5876 13302 5928 13354
rect 5928 13302 5930 13354
rect 5874 13300 5930 13302
rect 5978 13354 6034 13356
rect 5978 13302 5980 13354
rect 5980 13302 6032 13354
rect 6032 13302 6034 13354
rect 5978 13300 6034 13302
rect 6082 13354 6138 13356
rect 6082 13302 6084 13354
rect 6084 13302 6136 13354
rect 6136 13302 6138 13354
rect 6082 13300 6138 13302
rect 5874 11786 5930 11788
rect 5874 11734 5876 11786
rect 5876 11734 5928 11786
rect 5928 11734 5930 11786
rect 5874 11732 5930 11734
rect 5978 11786 6034 11788
rect 5978 11734 5980 11786
rect 5980 11734 6032 11786
rect 6032 11734 6034 11786
rect 5978 11732 6034 11734
rect 6082 11786 6138 11788
rect 6082 11734 6084 11786
rect 6084 11734 6136 11786
rect 6136 11734 6138 11786
rect 6082 11732 6138 11734
rect 14700 20748 14756 20804
rect 13916 19740 13972 19796
rect 12572 19628 12628 19684
rect 12460 19292 12516 19348
rect 13412 19404 13468 19460
rect 13916 19404 13972 19460
rect 14028 19292 14084 19348
rect 14252 19628 14308 19684
rect 14252 19292 14308 19348
rect 14364 19964 14420 20020
rect 13692 19180 13748 19236
rect 12908 18450 12964 18452
rect 12908 18398 12910 18450
rect 12910 18398 12962 18450
rect 12962 18398 12964 18450
rect 12908 18396 12964 18398
rect 13580 19122 13636 19124
rect 13580 19070 13582 19122
rect 13582 19070 13634 19122
rect 13634 19070 13636 19122
rect 13580 19068 13636 19070
rect 13244 18396 13300 18452
rect 12124 16940 12180 16996
rect 12684 17778 12740 17780
rect 12684 17726 12686 17778
rect 12686 17726 12738 17778
rect 12738 17726 12740 17778
rect 12684 17724 12740 17726
rect 13412 18450 13468 18452
rect 13412 18398 13414 18450
rect 13414 18398 13466 18450
rect 13466 18398 13468 18450
rect 13412 18396 13468 18398
rect 13580 17052 13636 17108
rect 13020 16940 13076 16996
rect 13804 18732 13860 18788
rect 14476 19234 14532 19236
rect 14476 19182 14478 19234
rect 14478 19182 14530 19234
rect 14530 19182 14532 19234
rect 14476 19180 14532 19182
rect 14028 19068 14084 19124
rect 13804 18450 13860 18452
rect 13804 18398 13806 18450
rect 13806 18398 13858 18450
rect 13858 18398 13860 18450
rect 13804 18396 13860 18398
rect 13860 17052 13916 17108
rect 11340 16098 11396 16100
rect 11340 16046 11342 16098
rect 11342 16046 11394 16098
rect 11394 16046 11396 16098
rect 11340 16044 11396 16046
rect 9212 13244 9268 13300
rect 7308 12402 7364 12404
rect 7308 12350 7310 12402
rect 7310 12350 7362 12402
rect 7362 12350 7364 12402
rect 7308 12348 7364 12350
rect 7644 12236 7700 12292
rect 8652 12348 8708 12404
rect 7084 11676 7140 11732
rect 8036 12178 8092 12180
rect 8036 12126 8038 12178
rect 8038 12126 8090 12178
rect 8090 12126 8092 12178
rect 8036 12124 8092 12126
rect 7868 12012 7924 12068
rect 5852 11564 5908 11620
rect 5874 10218 5930 10220
rect 5874 10166 5876 10218
rect 5876 10166 5928 10218
rect 5928 10166 5930 10218
rect 5874 10164 5930 10166
rect 5978 10218 6034 10220
rect 5978 10166 5980 10218
rect 5980 10166 6032 10218
rect 6032 10166 6034 10218
rect 5978 10164 6034 10166
rect 6082 10218 6138 10220
rect 6082 10166 6084 10218
rect 6084 10166 6136 10218
rect 6136 10166 6138 10218
rect 6082 10164 6138 10166
rect 7980 11228 8036 11284
rect 8316 10668 8372 10724
rect 7868 9884 7924 9940
rect 7084 8764 7140 8820
rect 5874 8650 5930 8652
rect 5874 8598 5876 8650
rect 5876 8598 5928 8650
rect 5928 8598 5930 8650
rect 5874 8596 5930 8598
rect 5978 8650 6034 8652
rect 5978 8598 5980 8650
rect 5980 8598 6032 8650
rect 6032 8598 6034 8650
rect 5978 8596 6034 8598
rect 6082 8650 6138 8652
rect 6082 8598 6084 8650
rect 6084 8598 6136 8650
rect 6136 8598 6138 8650
rect 6082 8596 6138 8598
rect 8204 9772 8260 9828
rect 8092 9660 8148 9716
rect 8428 10220 8484 10276
rect 8782 11340 8838 11396
rect 9044 11282 9100 11284
rect 9044 11230 9046 11282
rect 9046 11230 9098 11282
rect 9098 11230 9100 11282
rect 9044 11228 9100 11230
rect 9548 12738 9604 12740
rect 9548 12686 9550 12738
rect 9550 12686 9602 12738
rect 9602 12686 9604 12738
rect 9548 12684 9604 12686
rect 9884 12348 9940 12404
rect 9604 12178 9660 12180
rect 9604 12126 9606 12178
rect 9606 12126 9658 12178
rect 9658 12126 9660 12178
rect 9604 12124 9660 12126
rect 10536 14138 10592 14140
rect 10536 14086 10538 14138
rect 10538 14086 10590 14138
rect 10590 14086 10592 14138
rect 10536 14084 10592 14086
rect 10640 14138 10696 14140
rect 10640 14086 10642 14138
rect 10642 14086 10694 14138
rect 10694 14086 10696 14138
rect 10640 14084 10696 14086
rect 10744 14138 10800 14140
rect 10744 14086 10746 14138
rect 10746 14086 10798 14138
rect 10798 14086 10800 14138
rect 10744 14084 10800 14086
rect 10332 13468 10388 13524
rect 10220 12796 10276 12852
rect 10668 12684 10724 12740
rect 10536 12570 10592 12572
rect 10536 12518 10538 12570
rect 10538 12518 10590 12570
rect 10590 12518 10592 12570
rect 10536 12516 10592 12518
rect 10640 12570 10696 12572
rect 10640 12518 10642 12570
rect 10642 12518 10694 12570
rect 10694 12518 10696 12570
rect 10640 12516 10696 12518
rect 10744 12570 10800 12572
rect 10744 12518 10746 12570
rect 10746 12518 10798 12570
rect 10798 12518 10800 12570
rect 10744 12516 10800 12518
rect 10108 12236 10164 12292
rect 9324 11394 9380 11396
rect 9324 11342 9326 11394
rect 9326 11342 9378 11394
rect 9378 11342 9380 11394
rect 9324 11340 9380 11342
rect 8652 10610 8708 10612
rect 8652 10558 8654 10610
rect 8654 10558 8706 10610
rect 8706 10558 8708 10610
rect 8652 10556 8708 10558
rect 9436 10668 9492 10724
rect 9884 10444 9940 10500
rect 8746 9714 8802 9716
rect 8746 9662 8748 9714
rect 8748 9662 8800 9714
rect 8800 9662 8802 9714
rect 8746 9660 8802 9662
rect 9660 9884 9716 9940
rect 8988 9826 9044 9828
rect 8988 9774 8990 9826
rect 8990 9774 9042 9826
rect 9042 9774 9044 9826
rect 8988 9772 9044 9774
rect 9548 9100 9604 9156
rect 8204 8764 8260 8820
rect 5874 7082 5930 7084
rect 5874 7030 5876 7082
rect 5876 7030 5928 7082
rect 5928 7030 5930 7082
rect 5874 7028 5930 7030
rect 5978 7082 6034 7084
rect 5978 7030 5980 7082
rect 5980 7030 6032 7082
rect 6032 7030 6034 7082
rect 5978 7028 6034 7030
rect 6082 7082 6138 7084
rect 6082 7030 6084 7082
rect 6084 7030 6136 7082
rect 6136 7030 6138 7082
rect 6082 7028 6138 7030
rect 6524 6748 6580 6804
rect 5852 5906 5908 5908
rect 5852 5854 5854 5906
rect 5854 5854 5906 5906
rect 5906 5854 5908 5906
rect 5852 5852 5908 5854
rect 5874 5514 5930 5516
rect 5874 5462 5876 5514
rect 5876 5462 5928 5514
rect 5928 5462 5930 5514
rect 5874 5460 5930 5462
rect 5978 5514 6034 5516
rect 5978 5462 5980 5514
rect 5980 5462 6032 5514
rect 6032 5462 6034 5514
rect 5978 5460 6034 5462
rect 6082 5514 6138 5516
rect 6082 5462 6084 5514
rect 6084 5462 6136 5514
rect 6136 5462 6138 5514
rect 6082 5460 6138 5462
rect 6188 5180 6244 5236
rect 1148 3388 1204 3444
rect 4172 5094 4228 5124
rect 4172 5068 4174 5094
rect 4174 5068 4226 5094
rect 4226 5068 4228 5094
rect 3500 4956 3556 5012
rect 2772 4562 2828 4564
rect 2772 4510 2774 4562
rect 2774 4510 2826 4562
rect 2826 4510 2828 4562
rect 2772 4508 2828 4510
rect 7308 8316 7364 8372
rect 8316 8092 8372 8148
rect 8316 7532 8372 7588
rect 8148 7474 8204 7476
rect 8148 7422 8150 7474
rect 8150 7422 8202 7474
rect 8202 7422 8204 7474
rect 8148 7420 8204 7422
rect 7980 7196 8036 7252
rect 8652 8540 8708 8596
rect 8428 7196 8484 7252
rect 8540 8092 8596 8148
rect 9436 7980 9492 8036
rect 9044 7532 9100 7588
rect 8540 7308 8596 7364
rect 8540 6748 8596 6804
rect 9436 7308 9492 7364
rect 8894 6636 8950 6692
rect 8652 6524 8708 6580
rect 9660 8316 9716 8372
rect 9548 6524 9604 6580
rect 8316 5234 8372 5236
rect 8316 5182 8318 5234
rect 8318 5182 8370 5234
rect 8370 5182 8372 5234
rect 8316 5180 8372 5182
rect 10668 12290 10724 12292
rect 10668 12238 10670 12290
rect 10670 12238 10722 12290
rect 10722 12238 10724 12290
rect 10668 12236 10724 12238
rect 11004 12962 11060 12964
rect 11004 12910 11006 12962
rect 11006 12910 11058 12962
rect 11058 12910 11060 12962
rect 11004 12908 11060 12910
rect 12460 15314 12516 15316
rect 12460 15262 12462 15314
rect 12462 15262 12514 15314
rect 12514 15262 12516 15314
rect 12460 15260 12516 15262
rect 13468 15260 13524 15316
rect 10892 12236 10948 12292
rect 11004 12348 11060 12404
rect 11004 12178 11060 12180
rect 11004 12126 11006 12178
rect 11006 12126 11058 12178
rect 11058 12126 11060 12178
rect 11004 12124 11060 12126
rect 11452 12908 11508 12964
rect 11900 12684 11956 12740
rect 10668 11564 10724 11620
rect 10388 11394 10444 11396
rect 10388 11342 10390 11394
rect 10390 11342 10442 11394
rect 10442 11342 10444 11394
rect 10388 11340 10444 11342
rect 12068 12178 12124 12180
rect 12068 12126 12070 12178
rect 12070 12126 12122 12178
rect 12122 12126 12124 12178
rect 12068 12124 12124 12126
rect 13132 12066 13188 12068
rect 13132 12014 13134 12066
rect 13134 12014 13186 12066
rect 13186 12014 13188 12066
rect 13132 12012 13188 12014
rect 12236 11564 12292 11620
rect 12068 11394 12124 11396
rect 12068 11342 12070 11394
rect 12070 11342 12122 11394
rect 12122 11342 12124 11394
rect 12068 11340 12124 11342
rect 10536 11002 10592 11004
rect 10536 10950 10538 11002
rect 10538 10950 10590 11002
rect 10590 10950 10592 11002
rect 10536 10948 10592 10950
rect 10640 11002 10696 11004
rect 10640 10950 10642 11002
rect 10642 10950 10694 11002
rect 10694 10950 10696 11002
rect 10640 10948 10696 10950
rect 10744 11002 10800 11004
rect 10744 10950 10746 11002
rect 10746 10950 10798 11002
rect 10798 10950 10800 11002
rect 10744 10948 10800 10950
rect 10108 10780 10164 10836
rect 10220 10444 10276 10500
rect 10164 10220 10220 10276
rect 11228 10108 11284 10164
rect 10462 9996 10518 10052
rect 11788 9996 11844 10052
rect 9996 9100 10052 9156
rect 9940 8034 9996 8036
rect 9940 7982 9942 8034
rect 9942 7982 9994 8034
rect 9994 7982 9996 8034
rect 9940 7980 9996 7982
rect 9940 7474 9996 7476
rect 9940 7422 9942 7474
rect 9942 7422 9994 7474
rect 9994 7422 9996 7474
rect 9940 7420 9996 7422
rect 10536 9434 10592 9436
rect 10536 9382 10538 9434
rect 10538 9382 10590 9434
rect 10590 9382 10592 9434
rect 10536 9380 10592 9382
rect 10640 9434 10696 9436
rect 10640 9382 10642 9434
rect 10642 9382 10694 9434
rect 10694 9382 10696 9434
rect 10640 9380 10696 9382
rect 10744 9434 10800 9436
rect 10744 9382 10746 9434
rect 10746 9382 10798 9434
rect 10798 9382 10800 9434
rect 10744 9380 10800 9382
rect 12572 11452 12628 11508
rect 12814 11394 12870 11396
rect 12814 11342 12816 11394
rect 12816 11342 12868 11394
rect 12868 11342 12870 11394
rect 12814 11340 12870 11342
rect 13580 14754 13636 14756
rect 13580 14702 13582 14754
rect 13582 14702 13634 14754
rect 13634 14702 13636 14754
rect 13580 14700 13636 14702
rect 13580 13804 13636 13860
rect 14364 18732 14420 18788
rect 14140 18396 14196 18452
rect 14252 15260 14308 15316
rect 13692 13356 13748 13412
rect 13636 13132 13692 13188
rect 13636 12348 13692 12404
rect 14476 17164 14532 17220
rect 15198 21194 15254 21196
rect 15198 21142 15200 21194
rect 15200 21142 15252 21194
rect 15252 21142 15254 21194
rect 15198 21140 15254 21142
rect 15302 21194 15358 21196
rect 15302 21142 15304 21194
rect 15304 21142 15356 21194
rect 15356 21142 15358 21194
rect 15302 21140 15358 21142
rect 15406 21194 15462 21196
rect 15406 21142 15408 21194
rect 15408 21142 15460 21194
rect 15460 21142 15462 21194
rect 15406 21140 15462 21142
rect 16940 23154 16996 23156
rect 16940 23102 16942 23154
rect 16942 23102 16994 23154
rect 16994 23102 16996 23154
rect 16940 23100 16996 23102
rect 16828 22370 16884 22372
rect 16828 22318 16830 22370
rect 16830 22318 16882 22370
rect 16882 22318 16884 22370
rect 16828 22316 16884 22318
rect 16604 21868 16660 21924
rect 15596 19852 15652 19908
rect 15764 19740 15820 19796
rect 15198 19626 15254 19628
rect 15198 19574 15200 19626
rect 15200 19574 15252 19626
rect 15252 19574 15254 19626
rect 15198 19572 15254 19574
rect 15302 19626 15358 19628
rect 15302 19574 15304 19626
rect 15304 19574 15356 19626
rect 15356 19574 15358 19626
rect 15302 19572 15358 19574
rect 15406 19626 15462 19628
rect 15406 19574 15408 19626
rect 15408 19574 15460 19626
rect 15460 19574 15462 19626
rect 15406 19572 15462 19574
rect 14924 18732 14980 18788
rect 15198 18058 15254 18060
rect 15198 18006 15200 18058
rect 15200 18006 15252 18058
rect 15252 18006 15254 18058
rect 15198 18004 15254 18006
rect 15302 18058 15358 18060
rect 15302 18006 15304 18058
rect 15304 18006 15356 18058
rect 15356 18006 15358 18058
rect 15302 18004 15358 18006
rect 15406 18058 15462 18060
rect 15406 18006 15408 18058
rect 15408 18006 15460 18058
rect 15460 18006 15462 18058
rect 15406 18004 15462 18006
rect 15596 17164 15652 17220
rect 13916 14252 13972 14308
rect 14308 14306 14364 14308
rect 14308 14254 14310 14306
rect 14310 14254 14362 14306
rect 14362 14254 14364 14306
rect 14308 14252 14364 14254
rect 14476 14140 14532 14196
rect 15198 16490 15254 16492
rect 15198 16438 15200 16490
rect 15200 16438 15252 16490
rect 15252 16438 15254 16490
rect 15198 16436 15254 16438
rect 15302 16490 15358 16492
rect 15302 16438 15304 16490
rect 15304 16438 15356 16490
rect 15356 16438 15358 16490
rect 15302 16436 15358 16438
rect 15406 16490 15462 16492
rect 15406 16438 15408 16490
rect 15408 16438 15460 16490
rect 15460 16438 15462 16490
rect 15406 16436 15462 16438
rect 16380 16994 16436 16996
rect 16380 16942 16382 16994
rect 16382 16942 16434 16994
rect 16434 16942 16436 16994
rect 16380 16940 16436 16942
rect 16716 16380 16772 16436
rect 15198 14922 15254 14924
rect 15198 14870 15200 14922
rect 15200 14870 15252 14922
rect 15252 14870 15254 14922
rect 15198 14868 15254 14870
rect 15302 14922 15358 14924
rect 15302 14870 15304 14922
rect 15304 14870 15356 14922
rect 15356 14870 15358 14922
rect 15302 14868 15358 14870
rect 15406 14922 15462 14924
rect 15406 14870 15408 14922
rect 15408 14870 15460 14922
rect 15460 14870 15462 14922
rect 15406 14868 15462 14870
rect 14700 14140 14756 14196
rect 14924 13804 14980 13860
rect 14140 13356 14196 13412
rect 14028 13132 14084 13188
rect 13916 13020 13972 13076
rect 14196 13074 14252 13076
rect 14196 13022 14198 13074
rect 14198 13022 14250 13074
rect 14250 13022 14252 13074
rect 14196 13020 14252 13022
rect 14532 13356 14588 13412
rect 13804 12796 13860 12852
rect 14084 12178 14140 12180
rect 14084 12126 14086 12178
rect 14086 12126 14138 12178
rect 14138 12126 14140 12178
rect 14084 12124 14140 12126
rect 14140 11788 14196 11844
rect 14028 11394 14084 11396
rect 14028 11342 14030 11394
rect 14030 11342 14082 11394
rect 14082 11342 14084 11394
rect 14028 11340 14084 11342
rect 13748 11282 13804 11284
rect 13748 11230 13750 11282
rect 13750 11230 13802 11282
rect 13802 11230 13804 11282
rect 13748 11228 13804 11230
rect 13468 10556 13524 10612
rect 12572 10220 12628 10276
rect 12964 10108 13020 10164
rect 12964 9938 13020 9940
rect 12964 9886 12966 9938
rect 12966 9886 13018 9938
rect 13018 9886 13020 9938
rect 12964 9884 13020 9886
rect 12796 9660 12852 9716
rect 13524 9714 13580 9716
rect 13524 9662 13526 9714
rect 13526 9662 13578 9714
rect 13578 9662 13580 9714
rect 13524 9660 13580 9662
rect 14588 12684 14644 12740
rect 14364 12236 14420 12292
rect 14700 12348 14756 12404
rect 15708 13804 15764 13860
rect 15036 13356 15092 13412
rect 15198 13354 15254 13356
rect 15198 13302 15200 13354
rect 15200 13302 15252 13354
rect 15252 13302 15254 13354
rect 15198 13300 15254 13302
rect 15302 13354 15358 13356
rect 15302 13302 15304 13354
rect 15304 13302 15356 13354
rect 15356 13302 15358 13354
rect 15302 13300 15358 13302
rect 15406 13354 15462 13356
rect 15406 13302 15408 13354
rect 15408 13302 15460 13354
rect 15460 13302 15462 13354
rect 15406 13300 15462 13302
rect 16940 14530 16996 14532
rect 16940 14478 16942 14530
rect 16942 14478 16994 14530
rect 16994 14478 16996 14530
rect 16940 14476 16996 14478
rect 15036 12796 15092 12852
rect 14700 11788 14756 11844
rect 14588 11506 14644 11508
rect 14588 11454 14590 11506
rect 14590 11454 14642 11506
rect 14642 11454 14644 11506
rect 14588 11452 14644 11454
rect 14364 11228 14420 11284
rect 11060 7980 11116 8036
rect 10536 7866 10592 7868
rect 10536 7814 10538 7866
rect 10538 7814 10590 7866
rect 10590 7814 10592 7866
rect 10536 7812 10592 7814
rect 10640 7866 10696 7868
rect 10640 7814 10642 7866
rect 10642 7814 10694 7866
rect 10694 7814 10696 7866
rect 10640 7812 10696 7814
rect 10744 7866 10800 7868
rect 10744 7814 10746 7866
rect 10746 7814 10798 7866
rect 10798 7814 10800 7866
rect 10744 7812 10800 7814
rect 11060 7756 11116 7812
rect 10668 6690 10724 6692
rect 10668 6638 10670 6690
rect 10670 6638 10722 6690
rect 10722 6638 10724 6690
rect 10668 6636 10724 6638
rect 10892 7420 10948 7476
rect 10108 6412 10164 6468
rect 9996 6076 10052 6132
rect 8988 5180 9044 5236
rect 9100 5068 9156 5124
rect 3500 4508 3556 4564
rect 1932 3388 1988 3444
rect 2940 3388 2996 3444
rect 3500 3388 3556 3444
rect 5874 3946 5930 3948
rect 5874 3894 5876 3946
rect 5876 3894 5928 3946
rect 5928 3894 5930 3946
rect 5874 3892 5930 3894
rect 5978 3946 6034 3948
rect 5978 3894 5980 3946
rect 5980 3894 6032 3946
rect 6032 3894 6034 3946
rect 5978 3892 6034 3894
rect 6082 3946 6138 3948
rect 6082 3894 6084 3946
rect 6084 3894 6136 3946
rect 6136 3894 6138 3946
rect 6082 3892 6138 3894
rect 6524 4060 6580 4116
rect 7644 4898 7700 4900
rect 7644 4846 7646 4898
rect 7646 4846 7698 4898
rect 7698 4846 7700 4898
rect 7644 4844 7700 4846
rect 7532 4114 7588 4116
rect 7532 4062 7534 4114
rect 7534 4062 7586 4114
rect 7586 4062 7588 4114
rect 7532 4060 7588 4062
rect 10220 5234 10276 5236
rect 10220 5182 10222 5234
rect 10222 5182 10274 5234
rect 10274 5182 10276 5234
rect 10220 5180 10276 5182
rect 10536 6298 10592 6300
rect 10536 6246 10538 6298
rect 10538 6246 10590 6298
rect 10590 6246 10592 6298
rect 10536 6244 10592 6246
rect 10640 6298 10696 6300
rect 10640 6246 10642 6298
rect 10642 6246 10694 6298
rect 10694 6246 10696 6298
rect 10640 6244 10696 6246
rect 10744 6298 10800 6300
rect 10744 6246 10746 6298
rect 10746 6246 10798 6298
rect 10798 6246 10800 6298
rect 10744 6244 10800 6246
rect 11900 7474 11956 7476
rect 11900 7422 11902 7474
rect 11902 7422 11954 7474
rect 11954 7422 11956 7474
rect 11900 7420 11956 7422
rect 12124 7474 12180 7476
rect 12124 7422 12126 7474
rect 12126 7422 12178 7474
rect 12178 7422 12180 7474
rect 12124 7420 12180 7422
rect 12460 8204 12516 8260
rect 13804 8258 13860 8260
rect 13804 8206 13806 8258
rect 13806 8206 13858 8258
rect 13858 8206 13860 8258
rect 13804 8204 13860 8206
rect 13916 7644 13972 7700
rect 17612 30210 17668 30212
rect 17612 30158 17614 30210
rect 17614 30158 17666 30210
rect 17666 30158 17668 30210
rect 17612 30156 17668 30158
rect 17388 28588 17444 28644
rect 18956 33570 19012 33572
rect 18956 33518 18958 33570
rect 18958 33518 19010 33570
rect 19010 33518 19012 33570
rect 18956 33516 19012 33518
rect 19404 33180 19460 33236
rect 20076 33180 20132 33236
rect 20412 33180 20468 33236
rect 18396 32284 18452 32340
rect 19860 32954 19916 32956
rect 19860 32902 19862 32954
rect 19862 32902 19914 32954
rect 19914 32902 19916 32954
rect 19860 32900 19916 32902
rect 19964 32954 20020 32956
rect 19964 32902 19966 32954
rect 19966 32902 20018 32954
rect 20018 32902 20020 32954
rect 19964 32900 20020 32902
rect 20068 32954 20124 32956
rect 20068 32902 20070 32954
rect 20070 32902 20122 32954
rect 20122 32902 20124 32954
rect 20068 32900 20124 32902
rect 19628 32674 19684 32676
rect 19628 32622 19630 32674
rect 19630 32622 19682 32674
rect 19682 32622 19684 32674
rect 19628 32620 19684 32622
rect 19292 32284 19348 32340
rect 18844 32060 18900 32116
rect 20020 32562 20076 32564
rect 20020 32510 20022 32562
rect 20022 32510 20074 32562
rect 20074 32510 20076 32562
rect 20020 32508 20076 32510
rect 21084 35196 21140 35252
rect 21756 35532 21812 35588
rect 20076 32060 20132 32116
rect 19740 31836 19796 31892
rect 19964 31890 20020 31892
rect 19964 31838 19966 31890
rect 19966 31838 20018 31890
rect 20018 31838 20020 31890
rect 19964 31836 20020 31838
rect 19516 31164 19572 31220
rect 19516 30994 19572 30996
rect 19516 30942 19518 30994
rect 19518 30942 19570 30994
rect 19570 30942 19572 30994
rect 19516 30940 19572 30942
rect 18284 29484 18340 29540
rect 18396 29372 18452 29428
rect 17388 28364 17444 28420
rect 17276 27132 17332 27188
rect 17388 28140 17444 28196
rect 18676 29036 18732 29092
rect 19860 31386 19916 31388
rect 19860 31334 19862 31386
rect 19862 31334 19914 31386
rect 19914 31334 19916 31386
rect 19860 31332 19916 31334
rect 19964 31386 20020 31388
rect 19964 31334 19966 31386
rect 19966 31334 20018 31386
rect 20018 31334 20020 31386
rect 19964 31332 20020 31334
rect 20068 31386 20124 31388
rect 20068 31334 20070 31386
rect 20070 31334 20122 31386
rect 20122 31334 20124 31386
rect 20068 31332 20124 31334
rect 19852 31164 19908 31220
rect 20076 31052 20132 31108
rect 19964 30716 20020 30772
rect 19628 30210 19684 30212
rect 19628 30158 19630 30210
rect 19630 30158 19682 30210
rect 19682 30158 19684 30210
rect 19628 30156 19684 30158
rect 19516 29426 19572 29428
rect 19516 29374 19518 29426
rect 19518 29374 19570 29426
rect 19570 29374 19572 29426
rect 19516 29372 19572 29374
rect 19404 29148 19460 29204
rect 19124 28588 19180 28644
rect 18396 28476 18452 28532
rect 18060 28140 18116 28196
rect 18732 28140 18788 28196
rect 18284 28082 18340 28084
rect 18284 28030 18286 28082
rect 18286 28030 18338 28082
rect 18338 28030 18340 28082
rect 18284 28028 18340 28030
rect 17500 27804 17556 27860
rect 17500 27468 17556 27524
rect 17948 27858 18004 27860
rect 17948 27806 17950 27858
rect 17950 27806 18002 27858
rect 18002 27806 18004 27858
rect 17948 27804 18004 27806
rect 18956 28140 19012 28196
rect 19010 27858 19066 27860
rect 19010 27806 19012 27858
rect 19012 27806 19064 27858
rect 19064 27806 19066 27858
rect 19010 27804 19066 27806
rect 19628 29148 19684 29204
rect 19516 29036 19572 29092
rect 18396 27356 18452 27412
rect 20524 32562 20580 32564
rect 20524 32510 20526 32562
rect 20526 32510 20578 32562
rect 20578 32510 20580 32562
rect 20524 32508 20580 32510
rect 20636 31554 20692 31556
rect 20636 31502 20638 31554
rect 20638 31502 20690 31554
rect 20690 31502 20692 31554
rect 20636 31500 20692 31502
rect 21308 33180 21364 33236
rect 20860 31164 20916 31220
rect 22316 35196 22372 35252
rect 21868 35084 21924 35140
rect 22764 35756 22820 35812
rect 22652 34972 22708 35028
rect 22148 33346 22204 33348
rect 22148 33294 22150 33346
rect 22150 33294 22202 33346
rect 22202 33294 22204 33346
rect 22148 33292 22204 33294
rect 21756 32732 21812 32788
rect 22876 34860 22932 34916
rect 24522 36874 24578 36876
rect 24522 36822 24524 36874
rect 24524 36822 24576 36874
rect 24576 36822 24578 36874
rect 24522 36820 24578 36822
rect 24626 36874 24682 36876
rect 24626 36822 24628 36874
rect 24628 36822 24680 36874
rect 24680 36822 24682 36874
rect 24626 36820 24682 36822
rect 24730 36874 24786 36876
rect 24730 36822 24732 36874
rect 24732 36822 24784 36874
rect 24784 36822 24786 36874
rect 24730 36820 24786 36822
rect 24332 36540 24388 36596
rect 24556 35868 24612 35924
rect 24332 35756 24388 35812
rect 24052 35084 24108 35140
rect 24444 35474 24500 35476
rect 24444 35422 24446 35474
rect 24446 35422 24498 35474
rect 24498 35422 24500 35474
rect 24444 35420 24500 35422
rect 24522 35306 24578 35308
rect 24522 35254 24524 35306
rect 24524 35254 24576 35306
rect 24576 35254 24578 35306
rect 24522 35252 24578 35254
rect 24626 35306 24682 35308
rect 24626 35254 24628 35306
rect 24628 35254 24680 35306
rect 24680 35254 24682 35306
rect 24626 35252 24682 35254
rect 24730 35306 24786 35308
rect 24730 35254 24732 35306
rect 24732 35254 24784 35306
rect 24784 35254 24786 35306
rect 24730 35252 24786 35254
rect 24892 35084 24948 35140
rect 23324 34860 23380 34916
rect 23996 33740 24052 33796
rect 23996 33180 24052 33236
rect 23156 33068 23212 33124
rect 21532 31948 21588 32004
rect 21756 32172 21812 32228
rect 22372 31948 22428 32004
rect 23324 32620 23380 32676
rect 23996 32956 24052 33012
rect 23660 32396 23716 32452
rect 22764 32172 22820 32228
rect 23100 32284 23156 32340
rect 22092 31612 22148 31668
rect 20972 31052 21028 31108
rect 20188 30994 20244 30996
rect 20188 30942 20190 30994
rect 20190 30942 20242 30994
rect 20242 30942 20244 30994
rect 20188 30940 20244 30942
rect 20188 30492 20244 30548
rect 20188 30210 20244 30212
rect 20188 30158 20190 30210
rect 20190 30158 20242 30210
rect 20242 30158 20244 30210
rect 20188 30156 20244 30158
rect 20636 30492 20692 30548
rect 20412 30156 20468 30212
rect 19860 29818 19916 29820
rect 19860 29766 19862 29818
rect 19862 29766 19914 29818
rect 19914 29766 19916 29818
rect 19860 29764 19916 29766
rect 19964 29818 20020 29820
rect 19964 29766 19966 29818
rect 19966 29766 20018 29818
rect 20018 29766 20020 29818
rect 19964 29764 20020 29766
rect 20068 29818 20124 29820
rect 20068 29766 20070 29818
rect 20070 29766 20122 29818
rect 20122 29766 20124 29818
rect 20068 29764 20124 29766
rect 19908 29538 19964 29540
rect 19908 29486 19910 29538
rect 19910 29486 19962 29538
rect 19962 29486 19964 29538
rect 19908 29484 19964 29486
rect 20412 28642 20468 28644
rect 20412 28590 20414 28642
rect 20414 28590 20466 28642
rect 20466 28590 20468 28642
rect 20412 28588 20468 28590
rect 19860 28250 19916 28252
rect 19860 28198 19862 28250
rect 19862 28198 19914 28250
rect 19914 28198 19916 28250
rect 19860 28196 19916 28198
rect 19964 28250 20020 28252
rect 19964 28198 19966 28250
rect 19966 28198 20018 28250
rect 20018 28198 20020 28250
rect 19964 28196 20020 28198
rect 20068 28250 20124 28252
rect 20068 28198 20070 28250
rect 20070 28198 20122 28250
rect 20122 28198 20124 28250
rect 20068 28196 20124 28198
rect 19740 27804 19796 27860
rect 20076 27916 20132 27972
rect 19628 27580 19684 27636
rect 19292 27356 19348 27412
rect 18844 27074 18900 27076
rect 18844 27022 18846 27074
rect 18846 27022 18898 27074
rect 18898 27022 18900 27074
rect 18844 27020 18900 27022
rect 17388 26908 17444 26964
rect 17948 26908 18004 26964
rect 17276 26290 17332 26292
rect 17276 26238 17278 26290
rect 17278 26238 17330 26290
rect 17330 26238 17332 26290
rect 17276 26236 17332 26238
rect 17612 25788 17668 25844
rect 17836 24722 17892 24724
rect 17836 24670 17838 24722
rect 17838 24670 17890 24722
rect 17890 24670 17892 24722
rect 17836 24668 17892 24670
rect 17500 23938 17556 23940
rect 17500 23886 17502 23938
rect 17502 23886 17554 23938
rect 17554 23886 17556 23938
rect 17500 23884 17556 23886
rect 17836 23660 17892 23716
rect 17164 23324 17220 23380
rect 19068 26908 19124 26964
rect 19516 27020 19572 27076
rect 19180 26796 19236 26852
rect 18732 26236 18788 26292
rect 18620 25506 18676 25508
rect 18620 25454 18622 25506
rect 18622 25454 18674 25506
rect 18674 25454 18676 25506
rect 18620 25452 18676 25454
rect 18452 25282 18508 25284
rect 18452 25230 18454 25282
rect 18454 25230 18506 25282
rect 18506 25230 18508 25282
rect 18452 25228 18508 25230
rect 19180 25900 19236 25956
rect 20188 27858 20244 27860
rect 20188 27806 20190 27858
rect 20190 27806 20242 27858
rect 20242 27806 20244 27858
rect 20188 27804 20244 27806
rect 19572 26572 19628 26628
rect 19516 25900 19572 25956
rect 19292 25676 19348 25732
rect 19404 25788 19460 25844
rect 18116 24668 18172 24724
rect 18284 24780 18340 24836
rect 18956 25228 19012 25284
rect 17948 23324 18004 23380
rect 18060 23212 18116 23268
rect 17164 19346 17220 19348
rect 17164 19294 17166 19346
rect 17166 19294 17218 19346
rect 17218 19294 17220 19346
rect 17164 19292 17220 19294
rect 17500 19180 17556 19236
rect 17780 19234 17836 19236
rect 17780 19182 17782 19234
rect 17782 19182 17834 19234
rect 17834 19182 17836 19234
rect 17780 19180 17836 19182
rect 18340 23548 18396 23604
rect 19292 25228 19348 25284
rect 19124 24498 19180 24500
rect 19124 24446 19126 24498
rect 19126 24446 19178 24498
rect 19178 24446 19180 24498
rect 19124 24444 19180 24446
rect 19180 23938 19236 23940
rect 19180 23886 19182 23938
rect 19182 23886 19234 23938
rect 19234 23886 19236 23938
rect 19180 23884 19236 23886
rect 19860 26682 19916 26684
rect 19860 26630 19862 26682
rect 19862 26630 19914 26682
rect 19914 26630 19916 26682
rect 19860 26628 19916 26630
rect 19964 26682 20020 26684
rect 19964 26630 19966 26682
rect 19966 26630 20018 26682
rect 20018 26630 20020 26682
rect 19964 26628 20020 26630
rect 20068 26682 20124 26684
rect 20068 26630 20070 26682
rect 20070 26630 20122 26682
rect 20122 26630 20124 26682
rect 20068 26628 20124 26630
rect 19852 26348 19908 26404
rect 20076 26290 20132 26292
rect 20076 26238 20078 26290
rect 20078 26238 20130 26290
rect 20130 26238 20132 26290
rect 20076 26236 20132 26238
rect 20748 30380 20804 30436
rect 21028 30716 21084 30772
rect 21420 30604 21476 30660
rect 21532 30492 21588 30548
rect 20860 29484 20916 29540
rect 21196 29820 21252 29876
rect 20860 29314 20916 29316
rect 20860 29262 20862 29314
rect 20862 29262 20914 29314
rect 20914 29262 20916 29314
rect 20860 29260 20916 29262
rect 20972 28028 21028 28084
rect 21084 29484 21140 29540
rect 21196 29426 21252 29428
rect 21196 29374 21198 29426
rect 21198 29374 21250 29426
rect 21250 29374 21252 29426
rect 21196 29372 21252 29374
rect 21084 28700 21140 28756
rect 20524 26796 20580 26852
rect 20636 27804 20692 27860
rect 20300 26572 20356 26628
rect 20524 26348 20580 26404
rect 21420 30210 21476 30212
rect 21420 30158 21422 30210
rect 21422 30158 21474 30210
rect 21474 30158 21476 30210
rect 21420 30156 21476 30158
rect 22652 31724 22708 31780
rect 21700 30380 21756 30436
rect 22316 31500 22372 31556
rect 22876 30981 22878 30996
rect 22878 30981 22930 30996
rect 22930 30981 22932 30996
rect 22540 30380 22596 30436
rect 22876 30940 22932 30981
rect 22988 30268 23044 30324
rect 23324 31948 23380 32004
rect 24522 33738 24578 33740
rect 24522 33686 24524 33738
rect 24524 33686 24576 33738
rect 24576 33686 24578 33738
rect 24522 33684 24578 33686
rect 24626 33738 24682 33740
rect 24626 33686 24628 33738
rect 24628 33686 24680 33738
rect 24680 33686 24682 33738
rect 24626 33684 24682 33686
rect 24730 33738 24786 33740
rect 24730 33686 24732 33738
rect 24732 33686 24784 33738
rect 24784 33686 24786 33738
rect 24730 33684 24786 33686
rect 24276 33234 24332 33236
rect 24276 33182 24278 33234
rect 24278 33182 24330 33234
rect 24330 33182 24332 33234
rect 24276 33180 24332 33182
rect 25228 35673 25230 35700
rect 25230 35673 25282 35700
rect 25282 35673 25284 35700
rect 25228 35644 25284 35673
rect 25788 35420 25844 35476
rect 25564 35084 25620 35140
rect 25676 35196 25732 35252
rect 25116 33740 25172 33796
rect 25116 33404 25172 33460
rect 24612 32508 24668 32564
rect 24780 32620 24836 32676
rect 24108 32396 24164 32452
rect 24332 32396 24388 32452
rect 23996 31948 24052 32004
rect 23772 31778 23828 31780
rect 23772 31726 23774 31778
rect 23774 31726 23826 31778
rect 23826 31726 23828 31778
rect 23772 31724 23828 31726
rect 23436 31500 23492 31556
rect 23660 31052 23716 31108
rect 22708 29372 22764 29428
rect 21532 28812 21588 28868
rect 23100 28924 23156 28980
rect 22260 28866 22316 28868
rect 22260 28814 22262 28866
rect 22262 28814 22314 28866
rect 22314 28814 22316 28866
rect 22260 28812 22316 28814
rect 21308 27916 21364 27972
rect 22764 28754 22820 28756
rect 22764 28702 22766 28754
rect 22766 28702 22818 28754
rect 22818 28702 22820 28754
rect 22764 28700 22820 28702
rect 20748 27746 20804 27748
rect 20748 27694 20750 27746
rect 20750 27694 20802 27746
rect 20802 27694 20804 27746
rect 20748 27692 20804 27694
rect 21868 28530 21924 28532
rect 21868 28478 21870 28530
rect 21870 28478 21922 28530
rect 21922 28478 21924 28530
rect 21868 28476 21924 28478
rect 22148 28364 22204 28420
rect 21532 27692 21588 27748
rect 21756 28028 21812 28084
rect 21084 27132 21140 27188
rect 21644 27468 21700 27524
rect 20804 27074 20860 27076
rect 20804 27022 20806 27074
rect 20806 27022 20858 27074
rect 20858 27022 20860 27074
rect 20804 27020 20860 27022
rect 20748 26348 20804 26404
rect 21420 27132 21476 27188
rect 21644 27074 21700 27076
rect 21644 27022 21646 27074
rect 21646 27022 21698 27074
rect 21698 27022 21700 27074
rect 21644 27020 21700 27022
rect 20076 25452 20132 25508
rect 19852 25228 19908 25284
rect 19860 25114 19916 25116
rect 19860 25062 19862 25114
rect 19862 25062 19914 25114
rect 19914 25062 19916 25114
rect 19860 25060 19916 25062
rect 19964 25114 20020 25116
rect 19964 25062 19966 25114
rect 19966 25062 20018 25114
rect 20018 25062 20020 25114
rect 19964 25060 20020 25062
rect 20068 25114 20124 25116
rect 20068 25062 20070 25114
rect 20070 25062 20122 25114
rect 20122 25062 20124 25114
rect 20068 25060 20124 25062
rect 19516 24780 19572 24836
rect 19740 24668 19796 24724
rect 19404 23884 19460 23940
rect 18844 23548 18900 23604
rect 18956 23772 19012 23828
rect 18732 22482 18788 22484
rect 18732 22430 18734 22482
rect 18734 22430 18786 22482
rect 18786 22430 18788 22482
rect 18732 22428 18788 22430
rect 19292 23660 19348 23716
rect 19068 23154 19124 23156
rect 19068 23102 19070 23154
rect 19070 23102 19122 23154
rect 19122 23102 19124 23154
rect 19068 23100 19124 23102
rect 20692 25730 20748 25732
rect 20692 25678 20694 25730
rect 20694 25678 20746 25730
rect 20746 25678 20748 25730
rect 20692 25676 20748 25678
rect 20524 25340 20580 25396
rect 20412 25228 20468 25284
rect 21476 25282 21532 25284
rect 21476 25230 21478 25282
rect 21478 25230 21530 25282
rect 21530 25230 21532 25282
rect 21476 25228 21532 25230
rect 21308 24722 21364 24724
rect 21308 24670 21310 24722
rect 21310 24670 21362 24722
rect 21362 24670 21364 24722
rect 21308 24668 21364 24670
rect 20972 24610 21028 24612
rect 20972 24558 20974 24610
rect 20974 24558 21026 24610
rect 21026 24558 21028 24610
rect 20972 24556 21028 24558
rect 19860 23546 19916 23548
rect 19860 23494 19862 23546
rect 19862 23494 19914 23546
rect 19914 23494 19916 23546
rect 19860 23492 19916 23494
rect 19964 23546 20020 23548
rect 19964 23494 19966 23546
rect 19966 23494 20018 23546
rect 20018 23494 20020 23546
rect 19964 23492 20020 23494
rect 20068 23546 20124 23548
rect 20068 23494 20070 23546
rect 20070 23494 20122 23546
rect 20122 23494 20124 23546
rect 20068 23492 20124 23494
rect 20076 23266 20132 23268
rect 20076 23214 20078 23266
rect 20078 23214 20130 23266
rect 20130 23214 20132 23266
rect 20076 23212 20132 23214
rect 20524 24444 20580 24500
rect 20300 23100 20356 23156
rect 20748 23884 20804 23940
rect 19404 21586 19460 21588
rect 19404 21534 19406 21586
rect 19406 21534 19458 21586
rect 19458 21534 19460 21586
rect 19404 21532 19460 21534
rect 18956 20076 19012 20132
rect 18172 19292 18228 19348
rect 18844 18620 18900 18676
rect 19068 18620 19124 18676
rect 19180 18284 19236 18340
rect 19404 21026 19460 21028
rect 19404 20974 19406 21026
rect 19406 20974 19458 21026
rect 19458 20974 19460 21026
rect 19404 20972 19460 20974
rect 19516 19234 19572 19236
rect 19516 19182 19518 19234
rect 19518 19182 19570 19234
rect 19570 19182 19572 19234
rect 19516 19180 19572 19182
rect 19860 21978 19916 21980
rect 19860 21926 19862 21978
rect 19862 21926 19914 21978
rect 19914 21926 19916 21978
rect 19860 21924 19916 21926
rect 19964 21978 20020 21980
rect 19964 21926 19966 21978
rect 19966 21926 20018 21978
rect 20018 21926 20020 21978
rect 19964 21924 20020 21926
rect 20068 21978 20124 21980
rect 20068 21926 20070 21978
rect 20070 21926 20122 21978
rect 20122 21926 20124 21978
rect 20068 21924 20124 21926
rect 23100 28364 23156 28420
rect 23548 29932 23604 29988
rect 23436 28812 23492 28868
rect 23548 28588 23604 28644
rect 23772 30994 23828 30996
rect 23772 30942 23774 30994
rect 23774 30942 23826 30994
rect 23826 30942 23828 30994
rect 23772 30940 23828 30942
rect 24108 30994 24164 30996
rect 24108 30942 24110 30994
rect 24110 30942 24162 30994
rect 24162 30942 24164 30994
rect 24108 30940 24164 30942
rect 23996 30716 24052 30772
rect 23772 30210 23828 30212
rect 23772 30158 23774 30210
rect 23774 30158 23826 30210
rect 23826 30158 23828 30210
rect 23772 30156 23828 30158
rect 23772 29650 23828 29652
rect 23772 29598 23774 29650
rect 23774 29598 23826 29650
rect 23826 29598 23828 29650
rect 23772 29596 23828 29598
rect 23660 28700 23716 28756
rect 23492 28418 23548 28420
rect 23492 28366 23494 28418
rect 23494 28366 23546 28418
rect 23546 28366 23548 28418
rect 23492 28364 23548 28366
rect 23212 26572 23268 26628
rect 21756 25228 21812 25284
rect 22204 26012 22260 26068
rect 22092 24610 22148 24612
rect 22092 24558 22094 24610
rect 22094 24558 22146 24610
rect 22146 24558 22148 24610
rect 22092 24556 22148 24558
rect 21980 23938 22036 23940
rect 21980 23886 21982 23938
rect 21982 23886 22034 23938
rect 22034 23886 22036 23938
rect 21980 23884 22036 23886
rect 19796 21586 19852 21588
rect 19796 21534 19798 21586
rect 19798 21534 19850 21586
rect 19850 21534 19852 21586
rect 19796 21532 19852 21534
rect 21644 21586 21700 21588
rect 21644 21534 21646 21586
rect 21646 21534 21698 21586
rect 21698 21534 21700 21586
rect 21644 21532 21700 21534
rect 21980 21362 22036 21364
rect 21980 21310 21982 21362
rect 21982 21310 22034 21362
rect 22034 21310 22036 21362
rect 21980 21308 22036 21310
rect 21532 20972 21588 21028
rect 22316 23324 22372 23380
rect 24522 32170 24578 32172
rect 24522 32118 24524 32170
rect 24524 32118 24576 32170
rect 24576 32118 24578 32170
rect 24522 32116 24578 32118
rect 24626 32170 24682 32172
rect 24626 32118 24628 32170
rect 24628 32118 24680 32170
rect 24680 32118 24682 32170
rect 24626 32116 24682 32118
rect 24730 32170 24786 32172
rect 24730 32118 24732 32170
rect 24732 32118 24784 32170
rect 24784 32118 24786 32170
rect 24730 32116 24786 32118
rect 24724 30882 24780 30884
rect 24724 30830 24726 30882
rect 24726 30830 24778 30882
rect 24778 30830 24780 30882
rect 24724 30828 24780 30830
rect 24220 30604 24276 30660
rect 24522 30602 24578 30604
rect 24522 30550 24524 30602
rect 24524 30550 24576 30602
rect 24576 30550 24578 30602
rect 24522 30548 24578 30550
rect 24626 30602 24682 30604
rect 24626 30550 24628 30602
rect 24628 30550 24680 30602
rect 24680 30550 24682 30602
rect 24626 30548 24682 30550
rect 24730 30602 24786 30604
rect 24730 30550 24732 30602
rect 24732 30550 24784 30602
rect 24784 30550 24786 30602
rect 24730 30548 24786 30550
rect 25282 33346 25338 33348
rect 25282 33294 25284 33346
rect 25284 33294 25336 33346
rect 25336 33294 25338 33346
rect 25282 33292 25338 33294
rect 25116 32620 25172 32676
rect 25228 33068 25284 33124
rect 25004 32284 25060 32340
rect 25900 34972 25956 35028
rect 26684 35308 26740 35364
rect 27244 35196 27300 35252
rect 26012 34860 26068 34916
rect 28588 36540 28644 36596
rect 28028 35532 28084 35588
rect 27804 35196 27860 35252
rect 28140 35420 28196 35476
rect 27244 33740 27300 33796
rect 26292 33068 26348 33124
rect 26292 32620 26348 32676
rect 25564 32284 25620 32340
rect 25452 31052 25508 31108
rect 25564 30828 25620 30884
rect 24892 30492 24948 30548
rect 24668 30380 24724 30436
rect 23548 25564 23604 25620
rect 24332 30156 24388 30212
rect 23212 23212 23268 23268
rect 23548 25340 23604 25396
rect 22428 23154 22484 23156
rect 22428 23102 22430 23154
rect 22430 23102 22482 23154
rect 22482 23102 22484 23154
rect 22428 23100 22484 23102
rect 22652 21532 22708 21588
rect 20188 20914 20244 20916
rect 20188 20862 20190 20914
rect 20190 20862 20242 20914
rect 20242 20862 20244 20914
rect 20188 20860 20244 20862
rect 20188 20636 20244 20692
rect 19860 20410 19916 20412
rect 19860 20358 19862 20410
rect 19862 20358 19914 20410
rect 19914 20358 19916 20410
rect 19860 20356 19916 20358
rect 19964 20410 20020 20412
rect 19964 20358 19966 20410
rect 19966 20358 20018 20410
rect 20018 20358 20020 20410
rect 19964 20356 20020 20358
rect 20068 20410 20124 20412
rect 20068 20358 20070 20410
rect 20070 20358 20122 20410
rect 20122 20358 20124 20410
rect 20068 20356 20124 20358
rect 19908 20076 19964 20132
rect 20300 20524 20356 20580
rect 20188 19964 20244 20020
rect 20300 19404 20356 19460
rect 21756 20748 21812 20804
rect 21420 20524 21476 20580
rect 20524 19516 20580 19572
rect 21140 19794 21196 19796
rect 21140 19742 21142 19794
rect 21142 19742 21194 19794
rect 21194 19742 21196 19794
rect 21140 19740 21196 19742
rect 19740 19068 19796 19124
rect 18172 17836 18228 17892
rect 19404 18620 19460 18676
rect 18172 17666 18228 17668
rect 18172 17614 18174 17666
rect 18174 17614 18226 17666
rect 18226 17614 18228 17666
rect 18172 17612 18228 17614
rect 17724 16940 17780 16996
rect 18396 17052 18452 17108
rect 17276 16380 17332 16436
rect 18060 16604 18116 16660
rect 18788 16604 18844 16660
rect 18844 16156 18900 16212
rect 18060 15314 18116 15316
rect 18060 15262 18062 15314
rect 18062 15262 18114 15314
rect 18114 15262 18116 15314
rect 18060 15260 18116 15262
rect 17276 13356 17332 13412
rect 18172 13356 18228 13412
rect 17724 12962 17780 12964
rect 17724 12910 17726 12962
rect 17726 12910 17778 12962
rect 17778 12910 17780 12962
rect 17724 12908 17780 12910
rect 15198 11786 15254 11788
rect 15198 11734 15200 11786
rect 15200 11734 15252 11786
rect 15252 11734 15254 11786
rect 15198 11732 15254 11734
rect 15302 11786 15358 11788
rect 15302 11734 15304 11786
rect 15304 11734 15356 11786
rect 15356 11734 15358 11786
rect 15302 11732 15358 11734
rect 15406 11786 15462 11788
rect 15406 11734 15408 11786
rect 15408 11734 15460 11786
rect 15460 11734 15462 11786
rect 15406 11732 15462 11734
rect 15198 10218 15254 10220
rect 15198 10166 15200 10218
rect 15200 10166 15252 10218
rect 15252 10166 15254 10218
rect 15198 10164 15254 10166
rect 15302 10218 15358 10220
rect 15302 10166 15304 10218
rect 15304 10166 15356 10218
rect 15356 10166 15358 10218
rect 15302 10164 15358 10166
rect 15406 10218 15462 10220
rect 15406 10166 15408 10218
rect 15408 10166 15460 10218
rect 15460 10166 15462 10218
rect 15406 10164 15462 10166
rect 15484 9884 15540 9940
rect 15484 9212 15540 9268
rect 15198 8650 15254 8652
rect 15198 8598 15200 8650
rect 15200 8598 15252 8650
rect 15252 8598 15254 8650
rect 15198 8596 15254 8598
rect 15302 8650 15358 8652
rect 15302 8598 15304 8650
rect 15304 8598 15356 8650
rect 15356 8598 15358 8650
rect 15302 8596 15358 8598
rect 15406 8650 15462 8652
rect 15406 8598 15408 8650
rect 15408 8598 15460 8650
rect 15460 8598 15462 8650
rect 15406 8596 15462 8598
rect 12460 6748 12516 6804
rect 10444 5964 10500 6020
rect 11004 5906 11060 5908
rect 11004 5854 11006 5906
rect 11006 5854 11058 5906
rect 11058 5854 11060 5906
rect 11004 5852 11060 5854
rect 11004 5122 11060 5124
rect 11004 5070 11006 5122
rect 11006 5070 11058 5122
rect 11058 5070 11060 5122
rect 11004 5068 11060 5070
rect 12572 5068 12628 5124
rect 10108 4732 10164 4788
rect 10332 4956 10388 5012
rect 10536 4730 10592 4732
rect 10536 4678 10538 4730
rect 10538 4678 10590 4730
rect 10590 4678 10592 4730
rect 10536 4676 10592 4678
rect 10640 4730 10696 4732
rect 10640 4678 10642 4730
rect 10642 4678 10694 4730
rect 10694 4678 10696 4730
rect 10640 4676 10696 4678
rect 10744 4730 10800 4732
rect 10744 4678 10746 4730
rect 10746 4678 10798 4730
rect 10798 4678 10800 4730
rect 10744 4676 10800 4678
rect 11900 4284 11956 4340
rect 10536 3162 10592 3164
rect 10536 3110 10538 3162
rect 10538 3110 10590 3162
rect 10590 3110 10592 3162
rect 10536 3108 10592 3110
rect 10640 3162 10696 3164
rect 10640 3110 10642 3162
rect 10642 3110 10694 3162
rect 10694 3110 10696 3162
rect 10640 3108 10696 3110
rect 10744 3162 10800 3164
rect 10744 3110 10746 3162
rect 10746 3110 10798 3162
rect 10798 3110 10800 3162
rect 10744 3108 10800 3110
rect 10108 812 10164 868
rect 13356 4338 13412 4340
rect 13356 4286 13358 4338
rect 13358 4286 13410 4338
rect 13410 4286 13412 4338
rect 13356 4284 13412 4286
rect 13692 6018 13748 6020
rect 13692 5966 13694 6018
rect 13694 5966 13746 6018
rect 13746 5966 13748 6018
rect 13692 5964 13748 5966
rect 13580 5628 13636 5684
rect 14476 6076 14532 6132
rect 14588 7420 14644 7476
rect 14140 5964 14196 6020
rect 14252 5234 14308 5236
rect 14252 5182 14254 5234
rect 14254 5182 14306 5234
rect 14306 5182 14308 5234
rect 14252 5180 14308 5182
rect 13804 4508 13860 4564
rect 13916 3948 13972 4004
rect 13580 3554 13636 3556
rect 13580 3502 13582 3554
rect 13582 3502 13634 3554
rect 13634 3502 13636 3554
rect 13580 3500 13636 3502
rect 10892 812 10948 868
rect 15148 7474 15204 7476
rect 15148 7422 15150 7474
rect 15150 7422 15202 7474
rect 15202 7422 15204 7474
rect 15148 7420 15204 7422
rect 15540 7420 15596 7476
rect 15198 7082 15254 7084
rect 15198 7030 15200 7082
rect 15200 7030 15252 7082
rect 15252 7030 15254 7082
rect 15198 7028 15254 7030
rect 15302 7082 15358 7084
rect 15302 7030 15304 7082
rect 15304 7030 15356 7082
rect 15356 7030 15358 7082
rect 15302 7028 15358 7030
rect 15406 7082 15462 7084
rect 15406 7030 15408 7082
rect 15408 7030 15460 7082
rect 15460 7030 15462 7082
rect 15406 7028 15462 7030
rect 15354 6914 15410 6916
rect 15354 6862 15356 6914
rect 15356 6862 15408 6914
rect 15408 6862 15410 6914
rect 15354 6860 15410 6862
rect 15596 6690 15652 6692
rect 15596 6638 15598 6690
rect 15598 6638 15650 6690
rect 15650 6638 15652 6690
rect 15596 6636 15652 6638
rect 15148 5682 15204 5684
rect 15148 5630 15150 5682
rect 15150 5630 15202 5682
rect 15202 5630 15204 5682
rect 15148 5628 15204 5630
rect 15198 5514 15254 5516
rect 15198 5462 15200 5514
rect 15200 5462 15252 5514
rect 15252 5462 15254 5514
rect 15198 5460 15254 5462
rect 15302 5514 15358 5516
rect 15302 5462 15304 5514
rect 15304 5462 15356 5514
rect 15356 5462 15358 5514
rect 15302 5460 15358 5462
rect 15406 5514 15462 5516
rect 15406 5462 15408 5514
rect 15408 5462 15460 5514
rect 15460 5462 15462 5514
rect 15406 5460 15462 5462
rect 15484 5122 15540 5124
rect 15484 5070 15486 5122
rect 15486 5070 15538 5122
rect 15538 5070 15540 5122
rect 15484 5068 15540 5070
rect 17052 11452 17108 11508
rect 17276 12796 17332 12852
rect 19292 17500 19348 17556
rect 19964 19068 20020 19124
rect 19860 18842 19916 18844
rect 19860 18790 19862 18842
rect 19862 18790 19914 18842
rect 19914 18790 19916 18842
rect 19860 18788 19916 18790
rect 19964 18842 20020 18844
rect 19964 18790 19966 18842
rect 19966 18790 20018 18842
rect 20018 18790 20020 18842
rect 19964 18788 20020 18790
rect 20068 18842 20124 18844
rect 20068 18790 20070 18842
rect 20070 18790 20122 18842
rect 20122 18790 20124 18842
rect 20068 18788 20124 18790
rect 20188 18284 20244 18340
rect 20020 17554 20076 17556
rect 20020 17502 20022 17554
rect 20022 17502 20074 17554
rect 20074 17502 20076 17554
rect 20020 17500 20076 17502
rect 19860 17274 19916 17276
rect 19860 17222 19862 17274
rect 19862 17222 19914 17274
rect 19914 17222 19916 17274
rect 19860 17220 19916 17222
rect 19964 17274 20020 17276
rect 19964 17222 19966 17274
rect 19966 17222 20018 17274
rect 20018 17222 20020 17274
rect 19964 17220 20020 17222
rect 20068 17274 20124 17276
rect 20068 17222 20070 17274
rect 20070 17222 20122 17274
rect 20122 17222 20124 17274
rect 20068 17220 20124 17222
rect 20300 18396 20356 18452
rect 20636 18844 20692 18900
rect 20748 18284 20804 18340
rect 20524 18172 20580 18228
rect 21532 18450 21588 18452
rect 21532 18398 21534 18450
rect 21534 18398 21586 18450
rect 21586 18398 21588 18450
rect 21532 18396 21588 18398
rect 21084 18172 21140 18228
rect 20412 18060 20468 18116
rect 20412 17442 20468 17444
rect 20412 17390 20414 17442
rect 20414 17390 20466 17442
rect 20466 17390 20468 17442
rect 20412 17388 20468 17390
rect 19404 16940 19460 16996
rect 20300 17276 20356 17332
rect 19628 16828 19684 16884
rect 20524 17052 20580 17108
rect 20524 16858 20526 16884
rect 20526 16858 20578 16884
rect 20578 16858 20580 16884
rect 20524 16828 20580 16858
rect 19292 15260 19348 15316
rect 19628 15820 19684 15876
rect 19964 16044 20020 16100
rect 20972 17052 21028 17108
rect 20748 16716 20804 16772
rect 19860 15706 19916 15708
rect 19860 15654 19862 15706
rect 19862 15654 19914 15706
rect 19914 15654 19916 15706
rect 19860 15652 19916 15654
rect 19964 15706 20020 15708
rect 19964 15654 19966 15706
rect 19966 15654 20018 15706
rect 20018 15654 20020 15706
rect 19964 15652 20020 15654
rect 20068 15706 20124 15708
rect 20068 15654 20070 15706
rect 20070 15654 20122 15706
rect 20122 15654 20124 15706
rect 20068 15652 20124 15654
rect 21532 17388 21588 17444
rect 21756 19740 21812 19796
rect 21812 19458 21868 19460
rect 21812 19406 21814 19458
rect 21814 19406 21866 19458
rect 21866 19406 21868 19458
rect 21812 19404 21868 19406
rect 22092 18508 22148 18564
rect 21868 18060 21924 18116
rect 21756 17500 21812 17556
rect 21252 16882 21308 16884
rect 21252 16830 21254 16882
rect 21254 16830 21306 16882
rect 21306 16830 21308 16882
rect 21252 16828 21308 16830
rect 20860 16492 20916 16548
rect 20524 15820 20580 15876
rect 20804 15484 20860 15540
rect 20748 15260 20804 15316
rect 19404 14476 19460 14532
rect 19404 13916 19460 13972
rect 18340 12850 18396 12852
rect 18340 12798 18342 12850
rect 18342 12798 18394 12850
rect 18394 12798 18396 12850
rect 18340 12796 18396 12798
rect 18060 12124 18116 12180
rect 17668 11506 17724 11508
rect 17668 11454 17670 11506
rect 17670 11454 17722 11506
rect 17722 11454 17724 11506
rect 17668 11452 17724 11454
rect 18732 11394 18788 11396
rect 18732 11342 18734 11394
rect 18734 11342 18786 11394
rect 18786 11342 18788 11394
rect 18732 11340 18788 11342
rect 20076 14530 20132 14532
rect 20076 14478 20078 14530
rect 20078 14478 20130 14530
rect 20130 14478 20132 14530
rect 20076 14476 20132 14478
rect 20412 15036 20468 15092
rect 21756 17052 21812 17108
rect 22316 21308 22372 21364
rect 22428 19404 22484 19460
rect 22316 18172 22372 18228
rect 22540 18426 22542 18452
rect 22542 18426 22594 18452
rect 22594 18426 22596 18452
rect 22540 18396 22596 18426
rect 23436 23100 23492 23156
rect 24050 27356 24106 27412
rect 23884 27074 23940 27076
rect 23884 27022 23886 27074
rect 23886 27022 23938 27074
rect 23938 27022 23940 27074
rect 23884 27020 23940 27022
rect 24220 26908 24276 26964
rect 23772 26124 23828 26180
rect 23660 24108 23716 24164
rect 23660 23660 23716 23716
rect 23772 25564 23828 25620
rect 24220 25506 24276 25508
rect 24220 25454 24222 25506
rect 24222 25454 24274 25506
rect 24274 25454 24276 25506
rect 24220 25452 24276 25454
rect 23884 25228 23940 25284
rect 23884 24108 23940 24164
rect 24556 29596 24612 29652
rect 25004 29820 25060 29876
rect 24724 29314 24780 29316
rect 24724 29262 24726 29314
rect 24726 29262 24778 29314
rect 24778 29262 24780 29314
rect 24724 29260 24780 29262
rect 24522 29034 24578 29036
rect 24522 28982 24524 29034
rect 24524 28982 24576 29034
rect 24576 28982 24578 29034
rect 24522 28980 24578 28982
rect 24626 29034 24682 29036
rect 24626 28982 24628 29034
rect 24628 28982 24680 29034
rect 24680 28982 24682 29034
rect 24626 28980 24682 28982
rect 24730 29034 24786 29036
rect 24730 28982 24732 29034
rect 24732 28982 24784 29034
rect 24784 28982 24786 29034
rect 24730 28980 24786 28982
rect 24668 28812 24724 28868
rect 24500 28754 24556 28756
rect 24500 28702 24502 28754
rect 24502 28702 24554 28754
rect 24554 28702 24556 28754
rect 24500 28700 24556 28702
rect 24780 28700 24836 28756
rect 25508 29538 25564 29540
rect 25508 29486 25510 29538
rect 25510 29486 25562 29538
rect 25562 29486 25564 29538
rect 25508 29484 25564 29486
rect 25676 29484 25732 29540
rect 24668 27916 24724 27972
rect 24556 27858 24612 27860
rect 24556 27806 24558 27858
rect 24558 27806 24610 27858
rect 24610 27806 24612 27858
rect 24556 27804 24612 27806
rect 24522 27466 24578 27468
rect 24522 27414 24524 27466
rect 24524 27414 24576 27466
rect 24576 27414 24578 27466
rect 24522 27412 24578 27414
rect 24626 27466 24682 27468
rect 24626 27414 24628 27466
rect 24628 27414 24680 27466
rect 24680 27414 24682 27466
rect 24626 27412 24682 27414
rect 24730 27466 24786 27468
rect 24730 27414 24732 27466
rect 24732 27414 24784 27466
rect 24784 27414 24786 27466
rect 24730 27412 24786 27414
rect 25004 27804 25060 27860
rect 25004 27244 25060 27300
rect 25116 28364 25172 28420
rect 25788 29148 25844 29204
rect 26842 32620 26898 32676
rect 26684 32562 26740 32564
rect 26684 32510 26686 32562
rect 26686 32510 26738 32562
rect 26738 32510 26740 32562
rect 26684 32508 26740 32510
rect 27692 33404 27748 33460
rect 27804 33346 27860 33348
rect 27804 33294 27806 33346
rect 27806 33294 27858 33346
rect 27858 33294 27860 33346
rect 27804 33292 27860 33294
rect 28252 33628 28308 33684
rect 28532 34914 28588 34916
rect 28532 34862 28534 34914
rect 28534 34862 28586 34914
rect 28586 34862 28588 34914
rect 28532 34860 28588 34862
rect 29184 36090 29240 36092
rect 29184 36038 29186 36090
rect 29186 36038 29238 36090
rect 29238 36038 29240 36090
rect 29184 36036 29240 36038
rect 29288 36090 29344 36092
rect 29288 36038 29290 36090
rect 29290 36038 29342 36090
rect 29342 36038 29344 36090
rect 29288 36036 29344 36038
rect 29392 36090 29448 36092
rect 29392 36038 29394 36090
rect 29394 36038 29446 36090
rect 29446 36038 29448 36090
rect 29392 36036 29448 36038
rect 29036 35084 29092 35140
rect 29708 35196 29764 35252
rect 29036 34914 29092 34916
rect 29036 34862 29038 34914
rect 29038 34862 29090 34914
rect 29090 34862 29092 34914
rect 29036 34860 29092 34862
rect 27692 32732 27748 32788
rect 28028 33180 28084 33236
rect 26572 32284 26628 32340
rect 26124 31164 26180 31220
rect 26012 30156 26068 30212
rect 26460 30940 26516 30996
rect 26460 30268 26516 30324
rect 26124 30044 26180 30100
rect 26124 29484 26180 29540
rect 26012 29148 26068 29204
rect 25900 28812 25956 28868
rect 25583 27916 25639 27972
rect 25340 27858 25396 27860
rect 25340 27806 25342 27858
rect 25342 27806 25394 27858
rect 25394 27806 25396 27858
rect 25340 27804 25396 27806
rect 25116 27356 25172 27412
rect 25676 27692 25732 27748
rect 25564 27132 25620 27188
rect 25004 26908 25060 26964
rect 24892 26796 24948 26852
rect 24556 26178 24612 26180
rect 24556 26126 24558 26178
rect 24558 26126 24610 26178
rect 24610 26126 24612 26178
rect 24556 26124 24612 26126
rect 24522 25898 24578 25900
rect 24522 25846 24524 25898
rect 24524 25846 24576 25898
rect 24576 25846 24578 25898
rect 24522 25844 24578 25846
rect 24626 25898 24682 25900
rect 24626 25846 24628 25898
rect 24628 25846 24680 25898
rect 24680 25846 24682 25898
rect 24626 25844 24682 25846
rect 24730 25898 24786 25900
rect 24730 25846 24732 25898
rect 24732 25846 24784 25898
rect 24784 25846 24786 25898
rect 24730 25844 24786 25846
rect 24780 25676 24836 25732
rect 24780 25340 24836 25396
rect 24332 24668 24388 24724
rect 24522 24330 24578 24332
rect 24522 24278 24524 24330
rect 24524 24278 24576 24330
rect 24576 24278 24578 24330
rect 24522 24276 24578 24278
rect 24626 24330 24682 24332
rect 24626 24278 24628 24330
rect 24628 24278 24680 24330
rect 24680 24278 24682 24330
rect 24626 24276 24682 24278
rect 24730 24330 24786 24332
rect 24730 24278 24732 24330
rect 24732 24278 24784 24330
rect 24784 24278 24786 24330
rect 24730 24276 24786 24278
rect 24108 23996 24164 24052
rect 23548 22428 23604 22484
rect 23716 22370 23772 22372
rect 23716 22318 23718 22370
rect 23718 22318 23770 22370
rect 23770 22318 23772 22370
rect 23716 22316 23772 22318
rect 23436 22204 23492 22260
rect 23212 21532 23268 21588
rect 22764 21308 22820 21364
rect 24522 22762 24578 22764
rect 24522 22710 24524 22762
rect 24524 22710 24576 22762
rect 24576 22710 24578 22762
rect 24522 22708 24578 22710
rect 24626 22762 24682 22764
rect 24626 22710 24628 22762
rect 24628 22710 24680 22762
rect 24680 22710 24682 22762
rect 24626 22708 24682 22710
rect 24730 22762 24786 22764
rect 24730 22710 24732 22762
rect 24732 22710 24784 22762
rect 24784 22710 24786 22762
rect 24730 22708 24786 22710
rect 24522 21194 24578 21196
rect 24522 21142 24524 21194
rect 24524 21142 24576 21194
rect 24576 21142 24578 21194
rect 24522 21140 24578 21142
rect 24626 21194 24682 21196
rect 24626 21142 24628 21194
rect 24628 21142 24680 21194
rect 24680 21142 24682 21194
rect 24626 21140 24682 21142
rect 24730 21194 24786 21196
rect 24730 21142 24732 21194
rect 24732 21142 24784 21194
rect 24784 21142 24786 21194
rect 24730 21140 24786 21142
rect 25004 26460 25060 26516
rect 25564 26908 25620 26964
rect 25340 26460 25396 26516
rect 25676 26572 25732 26628
rect 26572 28028 26628 28084
rect 26460 27858 26516 27860
rect 26460 27806 26462 27858
rect 26462 27806 26514 27858
rect 26514 27806 26516 27858
rect 26460 27804 26516 27806
rect 26348 27356 26404 27412
rect 26012 27244 26068 27300
rect 26236 27132 26292 27188
rect 25900 26908 25956 26964
rect 26516 27074 26572 27076
rect 26516 27022 26518 27074
rect 26518 27022 26570 27074
rect 26570 27022 26572 27074
rect 26516 27020 26572 27022
rect 25788 26012 25844 26068
rect 25340 25676 25396 25732
rect 25004 25452 25060 25508
rect 26068 25506 26124 25508
rect 26068 25454 26070 25506
rect 26070 25454 26122 25506
rect 26122 25454 26124 25506
rect 26068 25452 26124 25454
rect 25788 25116 25844 25172
rect 25564 22428 25620 22484
rect 25676 22876 25732 22932
rect 25676 22370 25732 22372
rect 25676 22318 25678 22370
rect 25678 22318 25730 22370
rect 25730 22318 25732 22370
rect 25676 22316 25732 22318
rect 25340 21756 25396 21812
rect 26516 25116 26572 25172
rect 26516 24668 26572 24724
rect 26796 31164 26852 31220
rect 27020 31052 27076 31108
rect 28028 32396 28084 32452
rect 27916 30940 27972 30996
rect 28140 32060 28196 32116
rect 27076 30604 27132 30660
rect 28028 30828 28084 30884
rect 28028 29596 28084 29652
rect 27916 29260 27972 29316
rect 26796 29202 26852 29204
rect 26796 29150 26798 29202
rect 26798 29150 26850 29202
rect 26850 29150 26852 29202
rect 26796 29148 26852 29150
rect 26964 28364 27020 28420
rect 27132 27970 27188 27972
rect 27132 27918 27134 27970
rect 27134 27918 27186 27970
rect 27186 27918 27188 27970
rect 27132 27916 27188 27918
rect 28140 29260 28196 29316
rect 28140 28082 28196 28084
rect 28140 28030 28142 28082
rect 28142 28030 28194 28082
rect 28194 28030 28196 28082
rect 28140 28028 28196 28030
rect 28364 33404 28420 33460
rect 29184 34522 29240 34524
rect 29184 34470 29186 34522
rect 29186 34470 29238 34522
rect 29238 34470 29240 34522
rect 29184 34468 29240 34470
rect 29288 34522 29344 34524
rect 29288 34470 29290 34522
rect 29290 34470 29342 34522
rect 29342 34470 29344 34522
rect 29288 34468 29344 34470
rect 29392 34522 29448 34524
rect 29392 34470 29394 34522
rect 29394 34470 29446 34522
rect 29446 34470 29448 34522
rect 29392 34468 29448 34470
rect 28364 29596 28420 29652
rect 28476 29260 28532 29316
rect 28476 29036 28532 29092
rect 27356 27580 27412 27636
rect 27356 27074 27412 27076
rect 27356 27022 27358 27074
rect 27358 27022 27410 27074
rect 27410 27022 27412 27074
rect 27356 27020 27412 27022
rect 27244 26908 27300 26964
rect 27188 26514 27244 26516
rect 27188 26462 27190 26514
rect 27190 26462 27242 26514
rect 27242 26462 27244 26514
rect 27188 26460 27244 26462
rect 27020 26124 27076 26180
rect 25788 21644 25844 21700
rect 25228 21308 25284 21364
rect 23436 20076 23492 20132
rect 22876 20018 22932 20020
rect 22876 19966 22878 20018
rect 22878 19966 22930 20018
rect 22930 19966 22932 20018
rect 22876 19964 22932 19966
rect 24108 20524 24164 20580
rect 23996 20076 24052 20132
rect 23436 19740 23492 19796
rect 22988 19516 23044 19572
rect 22764 18508 22820 18564
rect 22988 19195 23044 19236
rect 22988 19180 22990 19195
rect 22990 19180 23042 19195
rect 23042 19180 23044 19195
rect 23772 19794 23828 19796
rect 23772 19742 23774 19794
rect 23774 19742 23826 19794
rect 23826 19742 23828 19794
rect 23772 19740 23828 19742
rect 23772 19516 23828 19572
rect 23100 18956 23156 19012
rect 23380 18562 23436 18564
rect 23380 18510 23382 18562
rect 23382 18510 23434 18562
rect 23434 18510 23436 18562
rect 23380 18508 23436 18510
rect 22876 18060 22932 18116
rect 22316 17276 22372 17332
rect 22652 17500 22708 17556
rect 21868 16716 21924 16772
rect 21308 16098 21364 16100
rect 21308 16046 21310 16098
rect 21310 16046 21362 16098
rect 21362 16046 21364 16098
rect 21308 16044 21364 16046
rect 21476 15820 21532 15876
rect 21122 15484 21178 15540
rect 21308 15036 21364 15092
rect 21142 14924 21198 14980
rect 21756 16492 21812 16548
rect 21868 16156 21924 16212
rect 21980 16604 22036 16660
rect 21756 16044 21812 16100
rect 21980 15820 22036 15876
rect 21644 15260 21700 15316
rect 21644 15036 21700 15092
rect 21308 14530 21364 14532
rect 21308 14478 21310 14530
rect 21310 14478 21362 14530
rect 21362 14478 21364 14530
rect 21308 14476 21364 14478
rect 19860 14138 19916 14140
rect 19860 14086 19862 14138
rect 19862 14086 19914 14138
rect 19914 14086 19916 14138
rect 19860 14084 19916 14086
rect 19964 14138 20020 14140
rect 19964 14086 19966 14138
rect 19966 14086 20018 14138
rect 20018 14086 20020 14138
rect 19964 14084 20020 14086
rect 20068 14138 20124 14140
rect 20068 14086 20070 14138
rect 20070 14086 20122 14138
rect 20122 14086 20124 14138
rect 20068 14084 20124 14086
rect 20860 14028 20916 14084
rect 20188 12908 20244 12964
rect 19860 12570 19916 12572
rect 19860 12518 19862 12570
rect 19862 12518 19914 12570
rect 19914 12518 19916 12570
rect 19860 12516 19916 12518
rect 19964 12570 20020 12572
rect 19964 12518 19966 12570
rect 19966 12518 20018 12570
rect 20018 12518 20020 12570
rect 19964 12516 20020 12518
rect 20068 12570 20124 12572
rect 20068 12518 20070 12570
rect 20070 12518 20122 12570
rect 20122 12518 20124 12570
rect 20068 12516 20124 12518
rect 19628 12178 19684 12180
rect 19628 12126 19630 12178
rect 19630 12126 19682 12178
rect 19682 12126 19684 12178
rect 19628 12124 19684 12126
rect 20524 12908 20580 12964
rect 20188 12124 20244 12180
rect 20412 12796 20468 12852
rect 21308 14028 21364 14084
rect 21644 13468 21700 13524
rect 21532 13356 21588 13412
rect 21980 14364 22036 14420
rect 21980 13356 22036 13412
rect 22222 16604 22278 16660
rect 22484 16380 22540 16436
rect 22316 15932 22372 15988
rect 22204 15820 22260 15876
rect 22204 14700 22260 14756
rect 22428 15314 22484 15316
rect 22428 15262 22430 15314
rect 22430 15262 22482 15314
rect 22482 15262 22484 15314
rect 22428 15260 22484 15262
rect 22764 16716 22820 16772
rect 23772 18508 23828 18564
rect 23996 19234 24052 19236
rect 23996 19182 23998 19234
rect 23998 19182 24050 19234
rect 24050 19182 24052 19234
rect 23996 19180 24052 19182
rect 24108 19740 24164 19796
rect 26348 22652 26404 22708
rect 26460 23100 26516 23156
rect 26012 22482 26068 22484
rect 26012 22430 26014 22482
rect 26014 22430 26066 22482
rect 26066 22430 26068 22482
rect 26012 22428 26068 22430
rect 27860 27356 27916 27412
rect 28252 27020 28308 27076
rect 28140 26460 28196 26516
rect 28196 26290 28252 26292
rect 28196 26238 28198 26290
rect 28198 26238 28250 26290
rect 28250 26238 28252 26290
rect 28196 26236 28252 26238
rect 28924 34242 28980 34244
rect 28924 34190 28926 34242
rect 28926 34190 28978 34242
rect 28978 34190 28980 34242
rect 28924 34188 28980 34190
rect 28700 30716 28756 30772
rect 28756 29148 28812 29204
rect 28588 28028 28644 28084
rect 28812 28924 28868 28980
rect 28644 27804 28700 27860
rect 29316 33068 29372 33124
rect 29184 32954 29240 32956
rect 29184 32902 29186 32954
rect 29186 32902 29238 32954
rect 29238 32902 29240 32954
rect 29184 32900 29240 32902
rect 29288 32954 29344 32956
rect 29288 32902 29290 32954
rect 29290 32902 29342 32954
rect 29342 32902 29344 32954
rect 29288 32900 29344 32902
rect 29392 32954 29448 32956
rect 29392 32902 29394 32954
rect 29394 32902 29446 32954
rect 29446 32902 29448 32954
rect 29392 32900 29448 32902
rect 29260 32732 29316 32788
rect 30716 36316 30772 36372
rect 30492 34914 30548 34916
rect 30492 34862 30494 34914
rect 30494 34862 30546 34914
rect 30546 34862 30548 34914
rect 30492 34860 30548 34862
rect 30044 34412 30100 34468
rect 29820 33740 29876 33796
rect 30586 33458 30642 33460
rect 30586 33406 30588 33458
rect 30588 33406 30640 33458
rect 30640 33406 30642 33458
rect 30586 33404 30642 33406
rect 29484 32284 29540 32340
rect 29184 31386 29240 31388
rect 29184 31334 29186 31386
rect 29186 31334 29238 31386
rect 29238 31334 29240 31386
rect 29184 31332 29240 31334
rect 29288 31386 29344 31388
rect 29288 31334 29290 31386
rect 29290 31334 29342 31386
rect 29342 31334 29344 31386
rect 29288 31332 29344 31334
rect 29392 31386 29448 31388
rect 29392 31334 29394 31386
rect 29394 31334 29446 31386
rect 29446 31334 29448 31386
rect 29392 31332 29448 31334
rect 29036 30994 29092 30996
rect 29036 30942 29038 30994
rect 29038 30942 29090 30994
rect 29090 30942 29092 30994
rect 29036 30940 29092 30942
rect 30156 32956 30212 33012
rect 30044 32732 30100 32788
rect 30380 31948 30436 32004
rect 30940 35644 30996 35700
rect 30828 34018 30884 34020
rect 30828 33966 30830 34018
rect 30830 33966 30882 34018
rect 30882 33966 30884 34018
rect 30828 33964 30884 33966
rect 30828 33404 30884 33460
rect 31388 36258 31444 36260
rect 31388 36206 31390 36258
rect 31390 36206 31442 36258
rect 31442 36206 31444 36258
rect 31388 36204 31444 36206
rect 31276 35698 31332 35700
rect 31276 35646 31278 35698
rect 31278 35646 31330 35698
rect 31330 35646 31332 35698
rect 31276 35644 31332 35646
rect 31164 35084 31220 35140
rect 31836 34914 31892 34916
rect 31836 34862 31838 34914
rect 31838 34862 31890 34914
rect 31890 34862 31892 34914
rect 31836 34860 31892 34862
rect 31052 33516 31108 33572
rect 31164 34076 31220 34132
rect 30940 32844 30996 32900
rect 31332 33852 31388 33908
rect 31724 34130 31780 34132
rect 31724 34078 31726 34130
rect 31726 34078 31778 34130
rect 31778 34078 31780 34130
rect 31724 34076 31780 34078
rect 31612 33516 31668 33572
rect 31164 32732 31220 32788
rect 31444 32674 31500 32676
rect 31444 32622 31446 32674
rect 31446 32622 31498 32674
rect 31498 32622 31500 32674
rect 31444 32620 31500 32622
rect 30828 32060 30884 32116
rect 30940 32284 30996 32340
rect 30716 31052 30772 31108
rect 29484 30210 29540 30212
rect 29484 30158 29486 30210
rect 29486 30158 29538 30210
rect 29538 30158 29540 30210
rect 29484 30156 29540 30158
rect 29876 30210 29932 30212
rect 29876 30158 29878 30210
rect 29878 30158 29930 30210
rect 29930 30158 29932 30210
rect 29876 30156 29932 30158
rect 29184 29818 29240 29820
rect 29184 29766 29186 29818
rect 29186 29766 29238 29818
rect 29238 29766 29240 29818
rect 29184 29764 29240 29766
rect 29288 29818 29344 29820
rect 29288 29766 29290 29818
rect 29290 29766 29342 29818
rect 29342 29766 29344 29818
rect 29288 29764 29344 29766
rect 29392 29818 29448 29820
rect 29392 29766 29394 29818
rect 29394 29766 29446 29818
rect 29446 29766 29448 29818
rect 29392 29764 29448 29766
rect 29092 29650 29148 29652
rect 29092 29598 29094 29650
rect 29094 29598 29146 29650
rect 29146 29598 29148 29650
rect 29092 29596 29148 29598
rect 29260 29484 29316 29540
rect 29372 29426 29428 29428
rect 29372 29374 29374 29426
rect 29374 29374 29426 29426
rect 29426 29374 29428 29426
rect 29372 29372 29428 29374
rect 29036 29148 29092 29204
rect 29372 29148 29428 29204
rect 29596 28642 29652 28644
rect 29596 28590 29598 28642
rect 29598 28590 29650 28642
rect 29650 28590 29652 28642
rect 29596 28588 29652 28590
rect 29184 28250 29240 28252
rect 29184 28198 29186 28250
rect 29186 28198 29238 28250
rect 29238 28198 29240 28250
rect 29184 28196 29240 28198
rect 29288 28250 29344 28252
rect 29288 28198 29290 28250
rect 29290 28198 29342 28250
rect 29342 28198 29344 28250
rect 29288 28196 29344 28198
rect 29392 28250 29448 28252
rect 29392 28198 29394 28250
rect 29394 28198 29446 28250
rect 29446 28198 29448 28250
rect 29392 28196 29448 28198
rect 29652 27746 29708 27748
rect 29652 27694 29654 27746
rect 29654 27694 29706 27746
rect 29706 27694 29708 27746
rect 29652 27692 29708 27694
rect 28476 26236 28532 26292
rect 30940 29596 30996 29652
rect 30380 29372 30436 29428
rect 30604 28924 30660 28980
rect 30156 27692 30212 27748
rect 30380 28476 30436 28532
rect 30492 27858 30548 27860
rect 30492 27806 30494 27858
rect 30494 27806 30546 27858
rect 30546 27806 30548 27858
rect 30492 27804 30548 27806
rect 31388 32396 31444 32452
rect 31500 31724 31556 31780
rect 33068 36204 33124 36260
rect 33180 34972 33236 35028
rect 32172 34076 32228 34132
rect 32060 34018 32116 34020
rect 32060 33966 32062 34018
rect 32062 33966 32114 34018
rect 32114 33966 32116 34018
rect 32060 33964 32116 33966
rect 32172 33404 32228 33460
rect 31836 32620 31892 32676
rect 31948 32284 32004 32340
rect 31724 31948 31780 32004
rect 30716 27580 30772 27636
rect 30828 27074 30884 27076
rect 30828 27022 30830 27074
rect 30830 27022 30882 27074
rect 30882 27022 30884 27074
rect 30828 27020 30884 27022
rect 28364 26124 28420 26180
rect 27916 25564 27972 25620
rect 28588 25564 28644 25620
rect 28028 25228 28084 25284
rect 27580 23938 27636 23940
rect 27580 23886 27582 23938
rect 27582 23886 27634 23938
rect 27634 23886 27636 23938
rect 27580 23884 27636 23886
rect 27132 23154 27188 23156
rect 27132 23102 27134 23154
rect 27134 23102 27186 23154
rect 27186 23102 27188 23154
rect 27132 23100 27188 23102
rect 27804 23324 27860 23380
rect 26012 22204 26068 22260
rect 24556 20076 24612 20132
rect 24444 19964 24500 20020
rect 24332 19516 24388 19572
rect 24522 19626 24578 19628
rect 24522 19574 24524 19626
rect 24524 19574 24576 19626
rect 24576 19574 24578 19626
rect 24522 19572 24578 19574
rect 24626 19626 24682 19628
rect 24626 19574 24628 19626
rect 24628 19574 24680 19626
rect 24680 19574 24682 19626
rect 24626 19572 24682 19574
rect 24730 19626 24786 19628
rect 24730 19574 24732 19626
rect 24732 19574 24784 19626
rect 24784 19574 24786 19626
rect 24730 19572 24786 19574
rect 25284 19404 25340 19460
rect 24108 18508 24164 18564
rect 23660 17500 23716 17556
rect 23044 17106 23100 17108
rect 23044 17054 23046 17106
rect 23046 17054 23098 17106
rect 23098 17054 23100 17106
rect 23044 17052 23100 17054
rect 23772 17052 23828 17108
rect 23660 16940 23716 16996
rect 23100 16098 23156 16100
rect 23100 16046 23102 16098
rect 23102 16046 23154 16098
rect 23154 16046 23156 16098
rect 23100 16044 23156 16046
rect 22876 15932 22932 15988
rect 23492 15874 23548 15876
rect 23492 15822 23494 15874
rect 23494 15822 23546 15874
rect 23546 15822 23548 15874
rect 23492 15820 23548 15822
rect 23940 16044 23996 16100
rect 23436 15260 23492 15316
rect 22764 14924 22820 14980
rect 22652 14530 22708 14532
rect 22652 14478 22654 14530
rect 22654 14478 22706 14530
rect 22706 14478 22708 14530
rect 22652 14476 22708 14478
rect 24612 18450 24668 18452
rect 24612 18398 24614 18450
rect 24614 18398 24666 18450
rect 24666 18398 24668 18450
rect 24612 18396 24668 18398
rect 25004 18620 25060 18676
rect 25452 19180 25508 19236
rect 25564 18620 25620 18676
rect 25228 18284 25284 18340
rect 24780 18172 24836 18228
rect 25564 18172 25620 18228
rect 24332 18060 24388 18116
rect 24522 18058 24578 18060
rect 24522 18006 24524 18058
rect 24524 18006 24576 18058
rect 24576 18006 24578 18058
rect 24522 18004 24578 18006
rect 24626 18058 24682 18060
rect 24626 18006 24628 18058
rect 24628 18006 24680 18058
rect 24680 18006 24682 18058
rect 24626 18004 24682 18006
rect 24730 18058 24786 18060
rect 24730 18006 24732 18058
rect 24732 18006 24784 18058
rect 24784 18006 24786 18058
rect 24730 18004 24786 18006
rect 24332 17836 24388 17892
rect 24220 17500 24276 17556
rect 25172 17666 25228 17668
rect 25172 17614 25174 17666
rect 25174 17614 25226 17666
rect 25226 17614 25228 17666
rect 25172 17612 25228 17614
rect 25452 17666 25508 17668
rect 25452 17614 25454 17666
rect 25454 17614 25506 17666
rect 25506 17614 25508 17666
rect 25452 17612 25508 17614
rect 25788 20972 25844 21028
rect 26796 21644 26852 21700
rect 26124 20802 26180 20804
rect 26124 20750 26126 20802
rect 26126 20750 26178 20802
rect 26178 20750 26180 20802
rect 26124 20748 26180 20750
rect 26236 20636 26292 20692
rect 26460 20972 26516 21028
rect 25900 19068 25956 19124
rect 26572 19234 26628 19236
rect 25788 18284 25844 18340
rect 25900 17388 25956 17444
rect 26012 17724 26068 17780
rect 25732 17164 25788 17220
rect 24332 16940 24388 16996
rect 25564 16940 25620 16996
rect 25732 16940 25788 16996
rect 26012 16882 26068 16884
rect 26012 16830 26014 16882
rect 26014 16830 26066 16882
rect 26066 16830 26068 16882
rect 26012 16828 26068 16830
rect 24522 16490 24578 16492
rect 24522 16438 24524 16490
rect 24524 16438 24576 16490
rect 24576 16438 24578 16490
rect 24522 16436 24578 16438
rect 24626 16490 24682 16492
rect 24626 16438 24628 16490
rect 24628 16438 24680 16490
rect 24680 16438 24682 16490
rect 24626 16436 24682 16438
rect 24730 16490 24786 16492
rect 24730 16438 24732 16490
rect 24732 16438 24784 16490
rect 24784 16438 24786 16490
rect 24730 16436 24786 16438
rect 24575 16098 24631 16100
rect 24575 16046 24577 16098
rect 24577 16046 24629 16098
rect 24629 16046 24631 16098
rect 24575 16044 24631 16046
rect 25452 16098 25508 16100
rect 25452 16046 25454 16098
rect 25454 16046 25506 16098
rect 25506 16046 25508 16098
rect 25452 16044 25508 16046
rect 24388 15260 24444 15316
rect 22876 13916 22932 13972
rect 23100 14364 23156 14420
rect 22316 13356 22372 13412
rect 21308 12962 21364 12964
rect 21308 12910 21310 12962
rect 21310 12910 21362 12962
rect 21362 12910 21364 12962
rect 21308 12908 21364 12910
rect 21084 11788 21140 11844
rect 20524 11340 20580 11396
rect 19860 11002 19916 11004
rect 19860 10950 19862 11002
rect 19862 10950 19914 11002
rect 19914 10950 19916 11002
rect 19860 10948 19916 10950
rect 19964 11002 20020 11004
rect 19964 10950 19966 11002
rect 19966 10950 20018 11002
rect 20018 10950 20020 11002
rect 19964 10948 20020 10950
rect 20068 11002 20124 11004
rect 20068 10950 20070 11002
rect 20070 10950 20122 11002
rect 20122 10950 20124 11002
rect 20068 10948 20124 10950
rect 22184 12796 22240 12852
rect 21980 11452 22036 11508
rect 19292 10610 19348 10612
rect 19292 10558 19294 10610
rect 19294 10558 19346 10610
rect 19346 10558 19348 10610
rect 19292 10556 19348 10558
rect 20524 10780 20580 10836
rect 21028 10834 21084 10836
rect 21028 10782 21030 10834
rect 21030 10782 21082 10834
rect 21082 10782 21084 10834
rect 21028 10780 21084 10782
rect 19740 10610 19796 10612
rect 19740 10558 19742 10610
rect 19742 10558 19794 10610
rect 19794 10558 19796 10610
rect 19740 10556 19796 10558
rect 16940 9548 16996 9604
rect 17556 9548 17612 9604
rect 18228 9266 18284 9268
rect 18228 9214 18230 9266
rect 18230 9214 18282 9266
rect 18282 9214 18284 9266
rect 18228 9212 18284 9214
rect 18732 8764 18788 8820
rect 16604 7756 16660 7812
rect 17164 7980 17220 8036
rect 17780 8034 17836 8036
rect 17780 7982 17782 8034
rect 17782 7982 17834 8034
rect 17834 7982 17836 8034
rect 17780 7980 17836 7982
rect 16268 6690 16324 6692
rect 15820 6076 15876 6132
rect 15372 4396 15428 4452
rect 16268 6638 16270 6690
rect 16270 6638 16322 6690
rect 16322 6638 16324 6690
rect 16268 6636 16324 6638
rect 16716 6860 16772 6916
rect 20076 9548 20132 9604
rect 19860 9434 19916 9436
rect 19860 9382 19862 9434
rect 19862 9382 19914 9434
rect 19914 9382 19916 9434
rect 19860 9380 19916 9382
rect 19964 9434 20020 9436
rect 19964 9382 19966 9434
rect 19966 9382 20018 9434
rect 20018 9382 20020 9434
rect 19964 9380 20020 9382
rect 20068 9434 20124 9436
rect 20068 9382 20070 9434
rect 20070 9382 20122 9434
rect 20122 9382 20124 9434
rect 20068 9380 20124 9382
rect 20468 9938 20524 9940
rect 20468 9886 20470 9938
rect 20470 9886 20522 9938
rect 20522 9886 20524 9938
rect 20468 9884 20524 9886
rect 20468 9548 20524 9604
rect 21868 9772 21924 9828
rect 19180 8818 19236 8820
rect 19180 8766 19182 8818
rect 19182 8766 19234 8818
rect 19234 8766 19236 8818
rect 19180 8764 19236 8766
rect 20076 8204 20132 8260
rect 22876 13468 22932 13524
rect 22988 13356 23044 13412
rect 23230 13746 23286 13748
rect 23230 13694 23232 13746
rect 23232 13694 23284 13746
rect 23284 13694 23286 13746
rect 23230 13692 23286 13694
rect 23100 13132 23156 13188
rect 23100 12908 23156 12964
rect 23212 13244 23268 13300
rect 22764 12796 22820 12852
rect 23324 13132 23380 13188
rect 23548 14028 23604 14084
rect 23940 13970 23996 13972
rect 23940 13918 23942 13970
rect 23942 13918 23994 13970
rect 23994 13918 23996 13970
rect 23940 13916 23996 13918
rect 23772 13746 23828 13748
rect 23772 13694 23774 13746
rect 23774 13694 23826 13746
rect 23826 13694 23828 13746
rect 23772 13692 23828 13694
rect 24108 13132 24164 13188
rect 23436 12796 23492 12852
rect 24522 14922 24578 14924
rect 24522 14870 24524 14922
rect 24524 14870 24576 14922
rect 24576 14870 24578 14922
rect 24522 14868 24578 14870
rect 24626 14922 24682 14924
rect 24626 14870 24628 14922
rect 24628 14870 24680 14922
rect 24680 14870 24682 14922
rect 24626 14868 24682 14870
rect 24730 14922 24786 14924
rect 24730 14870 24732 14922
rect 24732 14870 24784 14922
rect 24784 14870 24786 14922
rect 24730 14868 24786 14870
rect 26572 19182 26574 19234
rect 26574 19182 26626 19234
rect 26626 19182 26628 19234
rect 26572 19180 26628 19182
rect 26460 18172 26516 18228
rect 27132 21586 27188 21588
rect 27132 21534 27134 21586
rect 27134 21534 27186 21586
rect 27186 21534 27188 21586
rect 27132 21532 27188 21534
rect 26908 20972 26964 21028
rect 27580 22428 27636 22484
rect 29184 26682 29240 26684
rect 29184 26630 29186 26682
rect 29186 26630 29238 26682
rect 29238 26630 29240 26682
rect 29184 26628 29240 26630
rect 29288 26682 29344 26684
rect 29288 26630 29290 26682
rect 29290 26630 29342 26682
rect 29342 26630 29344 26682
rect 29288 26628 29344 26630
rect 29392 26682 29448 26684
rect 29392 26630 29394 26682
rect 29394 26630 29446 26682
rect 29446 26630 29448 26682
rect 29392 26628 29448 26630
rect 29428 25452 29484 25508
rect 29184 25114 29240 25116
rect 29184 25062 29186 25114
rect 29186 25062 29238 25114
rect 29238 25062 29240 25114
rect 29184 25060 29240 25062
rect 29288 25114 29344 25116
rect 29288 25062 29290 25114
rect 29290 25062 29342 25114
rect 29342 25062 29344 25114
rect 29288 25060 29344 25062
rect 29392 25114 29448 25116
rect 29392 25062 29394 25114
rect 29394 25062 29446 25114
rect 29446 25062 29448 25114
rect 29392 25060 29448 25062
rect 29932 25506 29988 25508
rect 29932 25454 29934 25506
rect 29934 25454 29986 25506
rect 29986 25454 29988 25506
rect 29932 25452 29988 25454
rect 29820 25004 29876 25060
rect 29036 24892 29092 24948
rect 29820 24722 29876 24724
rect 29820 24670 29822 24722
rect 29822 24670 29874 24722
rect 29874 24670 29876 24722
rect 29820 24668 29876 24670
rect 28028 23436 28084 23492
rect 29036 24108 29092 24164
rect 28252 23938 28308 23940
rect 28252 23886 28254 23938
rect 28254 23886 28306 23938
rect 28306 23886 28308 23938
rect 28252 23884 28308 23886
rect 28644 23436 28700 23492
rect 28924 23436 28980 23492
rect 29036 23884 29092 23940
rect 29652 24108 29708 24164
rect 29820 23996 29876 24052
rect 29372 23884 29428 23940
rect 29184 23546 29240 23548
rect 29184 23494 29186 23546
rect 29186 23494 29238 23546
rect 29238 23494 29240 23546
rect 29184 23492 29240 23494
rect 29288 23546 29344 23548
rect 29288 23494 29290 23546
rect 29290 23494 29342 23546
rect 29342 23494 29344 23546
rect 29288 23492 29344 23494
rect 29392 23546 29448 23548
rect 29392 23494 29394 23546
rect 29394 23494 29446 23546
rect 29446 23494 29448 23546
rect 29392 23492 29448 23494
rect 27468 20972 27524 21028
rect 27076 20578 27132 20580
rect 27076 20526 27078 20578
rect 27078 20526 27130 20578
rect 27130 20526 27132 20578
rect 27076 20524 27132 20526
rect 26908 18284 26964 18340
rect 26684 17836 26740 17892
rect 27076 17836 27132 17892
rect 26572 17724 26628 17780
rect 27188 17724 27244 17780
rect 26684 17500 26740 17556
rect 26292 16882 26348 16884
rect 26292 16830 26294 16882
rect 26294 16830 26346 16882
rect 26346 16830 26348 16882
rect 26292 16828 26348 16830
rect 26684 17164 26740 17220
rect 27412 16380 27468 16436
rect 27692 18338 27748 18340
rect 27692 18286 27694 18338
rect 27694 18286 27746 18338
rect 27746 18286 27748 18338
rect 27692 18284 27748 18286
rect 28084 21474 28140 21476
rect 28084 21422 28086 21474
rect 28086 21422 28138 21474
rect 28138 21422 28140 21474
rect 28084 21420 28140 21422
rect 28700 21644 28756 21700
rect 29148 22652 29204 22708
rect 28588 21586 28644 21588
rect 28588 21534 28590 21586
rect 28590 21534 28642 21586
rect 28642 21534 28644 21586
rect 28588 21532 28644 21534
rect 28924 21644 28980 21700
rect 30324 26402 30380 26404
rect 30324 26350 30326 26402
rect 30326 26350 30378 26402
rect 30378 26350 30380 26402
rect 30324 26348 30380 26350
rect 30604 26684 30660 26740
rect 30380 25228 30436 25284
rect 30156 24834 30212 24836
rect 30156 24782 30158 24834
rect 30158 24782 30210 24834
rect 30210 24782 30212 24834
rect 30156 24780 30212 24782
rect 30268 24668 30324 24724
rect 31164 27244 31220 27300
rect 30940 26348 30996 26404
rect 31052 26908 31108 26964
rect 31276 27132 31332 27188
rect 31276 26796 31332 26852
rect 31668 27858 31724 27860
rect 31668 27806 31670 27858
rect 31670 27806 31722 27858
rect 31722 27806 31724 27858
rect 31668 27804 31724 27806
rect 31500 27020 31556 27076
rect 31500 26796 31556 26852
rect 31612 26684 31668 26740
rect 30828 25116 30884 25172
rect 30716 23996 30772 24052
rect 30380 23324 30436 23380
rect 30156 23212 30212 23268
rect 30044 22204 30100 22260
rect 29184 21978 29240 21980
rect 29184 21926 29186 21978
rect 29186 21926 29238 21978
rect 29238 21926 29240 21978
rect 29184 21924 29240 21926
rect 29288 21978 29344 21980
rect 29288 21926 29290 21978
rect 29290 21926 29342 21978
rect 29342 21926 29344 21978
rect 29288 21924 29344 21926
rect 29392 21978 29448 21980
rect 29392 21926 29394 21978
rect 29394 21926 29446 21978
rect 29446 21926 29448 21978
rect 29392 21924 29448 21926
rect 29036 21532 29092 21588
rect 30156 21586 30212 21588
rect 30156 21534 30158 21586
rect 30158 21534 30210 21586
rect 30210 21534 30212 21586
rect 30492 23212 30548 23268
rect 30940 23938 30996 23940
rect 30940 23886 30942 23938
rect 30942 23886 30994 23938
rect 30994 23886 30996 23938
rect 30940 23884 30996 23886
rect 31164 25900 31220 25956
rect 30492 22370 30548 22372
rect 30492 22318 30494 22370
rect 30494 22318 30546 22370
rect 30546 22318 30548 22370
rect 30492 22316 30548 22318
rect 31052 23154 31108 23156
rect 31052 23102 31054 23154
rect 31054 23102 31106 23154
rect 31106 23102 31108 23154
rect 31052 23100 31108 23102
rect 30716 22092 30772 22148
rect 30492 21980 30548 22036
rect 30156 21532 30212 21534
rect 30604 21196 30660 21252
rect 29184 20410 29240 20412
rect 29184 20358 29186 20410
rect 29186 20358 29238 20410
rect 29238 20358 29240 20410
rect 29184 20356 29240 20358
rect 29288 20410 29344 20412
rect 29288 20358 29290 20410
rect 29290 20358 29342 20410
rect 29342 20358 29344 20410
rect 29288 20356 29344 20358
rect 29392 20410 29448 20412
rect 29392 20358 29394 20410
rect 29394 20358 29446 20410
rect 29446 20358 29448 20410
rect 29392 20356 29448 20358
rect 28812 20188 28868 20244
rect 29036 20018 29092 20020
rect 29036 19966 29038 20018
rect 29038 19966 29090 20018
rect 29090 19966 29092 20018
rect 29036 19964 29092 19966
rect 29540 20018 29596 20020
rect 29540 19966 29542 20018
rect 29542 19966 29594 20018
rect 29594 19966 29596 20018
rect 29540 19964 29596 19966
rect 29932 19852 29988 19908
rect 29260 19516 29316 19572
rect 29484 19740 29540 19796
rect 29820 19740 29876 19796
rect 29820 19516 29876 19572
rect 29148 19234 29204 19236
rect 29148 19182 29150 19234
rect 29150 19182 29202 19234
rect 29202 19182 29204 19234
rect 29148 19180 29204 19182
rect 29036 18844 29092 18900
rect 29184 18842 29240 18844
rect 29184 18790 29186 18842
rect 29186 18790 29238 18842
rect 29238 18790 29240 18842
rect 29184 18788 29240 18790
rect 29288 18842 29344 18844
rect 29288 18790 29290 18842
rect 29290 18790 29342 18842
rect 29342 18790 29344 18842
rect 29288 18788 29344 18790
rect 29392 18842 29448 18844
rect 29392 18790 29394 18842
rect 29394 18790 29446 18842
rect 29446 18790 29448 18842
rect 29392 18788 29448 18790
rect 30268 20076 30324 20132
rect 30604 19740 30660 19796
rect 30492 19516 30548 19572
rect 30548 19234 30604 19236
rect 30548 19182 30550 19234
rect 30550 19182 30602 19234
rect 30602 19182 30604 19234
rect 30548 19180 30604 19182
rect 31052 22092 31108 22148
rect 31276 25228 31332 25284
rect 31724 26124 31780 26180
rect 31500 26012 31556 26068
rect 32284 32284 32340 32340
rect 32172 31164 32228 31220
rect 32284 31052 32340 31108
rect 32732 33964 32788 34020
rect 32956 33628 33012 33684
rect 33846 36874 33902 36876
rect 33846 36822 33848 36874
rect 33848 36822 33900 36874
rect 33900 36822 33902 36874
rect 33846 36820 33902 36822
rect 33950 36874 34006 36876
rect 33950 36822 33952 36874
rect 33952 36822 34004 36874
rect 34004 36822 34006 36874
rect 33950 36820 34006 36822
rect 34054 36874 34110 36876
rect 34054 36822 34056 36874
rect 34056 36822 34108 36874
rect 34108 36822 34110 36874
rect 34054 36820 34110 36822
rect 33846 35306 33902 35308
rect 33846 35254 33848 35306
rect 33848 35254 33900 35306
rect 33900 35254 33902 35306
rect 33846 35252 33902 35254
rect 33950 35306 34006 35308
rect 33950 35254 33952 35306
rect 33952 35254 34004 35306
rect 34004 35254 34006 35306
rect 33950 35252 34006 35254
rect 34054 35306 34110 35308
rect 34054 35254 34056 35306
rect 34056 35254 34108 35306
rect 34108 35254 34110 35306
rect 34054 35252 34110 35254
rect 34412 35084 34468 35140
rect 33740 34860 33796 34916
rect 33964 34412 34020 34468
rect 33628 33852 33684 33908
rect 35084 36258 35140 36260
rect 35084 36206 35086 36258
rect 35086 36206 35138 36258
rect 35138 36206 35140 36258
rect 35084 36204 35140 36206
rect 35532 34972 35588 35028
rect 35420 34914 35476 34916
rect 35420 34862 35422 34914
rect 35422 34862 35474 34914
rect 35474 34862 35476 34914
rect 35420 34860 35476 34862
rect 35308 34748 35364 34804
rect 33964 33852 34020 33908
rect 33846 33738 33902 33740
rect 33846 33686 33848 33738
rect 33848 33686 33900 33738
rect 33900 33686 33902 33738
rect 33846 33684 33902 33686
rect 33950 33738 34006 33740
rect 33950 33686 33952 33738
rect 33952 33686 34004 33738
rect 34004 33686 34006 33738
rect 33950 33684 34006 33686
rect 34054 33738 34110 33740
rect 34054 33686 34056 33738
rect 34056 33686 34108 33738
rect 34108 33686 34110 33738
rect 34054 33684 34110 33686
rect 34188 33740 34244 33796
rect 33404 33068 33460 33124
rect 33404 32396 33460 32452
rect 32620 30268 32676 30324
rect 32396 30044 32452 30100
rect 32060 29932 32116 29988
rect 32508 29708 32564 29764
rect 32060 29596 32116 29652
rect 32060 28924 32116 28980
rect 32060 28642 32116 28644
rect 32060 28590 32062 28642
rect 32062 28590 32114 28642
rect 32114 28590 32116 28642
rect 32060 28588 32116 28590
rect 32302 28530 32358 28532
rect 32302 28478 32304 28530
rect 32304 28478 32356 28530
rect 32356 28478 32358 28530
rect 32302 28476 32358 28478
rect 32172 28364 32228 28420
rect 32844 29036 32900 29092
rect 32844 28812 32900 28868
rect 32732 28700 32788 28756
rect 33162 31164 33218 31220
rect 33404 30994 33460 30996
rect 33404 30942 33406 30994
rect 33406 30942 33458 30994
rect 33458 30942 33460 30994
rect 33404 30940 33460 30942
rect 33404 30716 33460 30772
rect 33236 30044 33292 30100
rect 34076 32450 34132 32452
rect 34076 32398 34078 32450
rect 34078 32398 34130 32450
rect 34130 32398 34132 32450
rect 34076 32396 34132 32398
rect 33846 32170 33902 32172
rect 33846 32118 33848 32170
rect 33848 32118 33900 32170
rect 33900 32118 33902 32170
rect 33846 32116 33902 32118
rect 33950 32170 34006 32172
rect 33950 32118 33952 32170
rect 33952 32118 34004 32170
rect 34004 32118 34006 32170
rect 33950 32116 34006 32118
rect 34054 32170 34110 32172
rect 34054 32118 34056 32170
rect 34056 32118 34108 32170
rect 34108 32118 34110 32170
rect 34054 32116 34110 32118
rect 34412 33234 34468 33236
rect 34412 33182 34414 33234
rect 34414 33182 34466 33234
rect 34466 33182 34468 33234
rect 34412 33180 34468 33182
rect 34412 32620 34468 32676
rect 34300 32508 34356 32564
rect 34300 31948 34356 32004
rect 33908 30828 33964 30884
rect 33846 30602 33902 30604
rect 33846 30550 33848 30602
rect 33848 30550 33900 30602
rect 33900 30550 33902 30602
rect 33846 30548 33902 30550
rect 33950 30602 34006 30604
rect 33950 30550 33952 30602
rect 33952 30550 34004 30602
rect 34004 30550 34006 30602
rect 33950 30548 34006 30550
rect 34054 30602 34110 30604
rect 34054 30550 34056 30602
rect 34056 30550 34108 30602
rect 34108 30550 34110 30602
rect 34054 30548 34110 30550
rect 33068 28642 33124 28644
rect 33068 28590 33070 28642
rect 33070 28590 33122 28642
rect 33122 28590 33124 28642
rect 33068 28588 33124 28590
rect 32396 27244 32452 27300
rect 32060 26908 32116 26964
rect 31836 25900 31892 25956
rect 31836 25676 31892 25732
rect 31500 25340 31556 25396
rect 31388 24892 31444 24948
rect 31724 25228 31780 25284
rect 32508 27132 32564 27188
rect 32284 25228 32340 25284
rect 32396 26124 32452 26180
rect 31388 24722 31444 24724
rect 31388 24670 31390 24722
rect 31390 24670 31442 24722
rect 31442 24670 31444 24722
rect 31388 24668 31444 24670
rect 32060 24668 32116 24724
rect 31724 24610 31780 24612
rect 31724 24558 31726 24610
rect 31726 24558 31778 24610
rect 31778 24558 31780 24610
rect 31724 24556 31780 24558
rect 31724 24332 31780 24388
rect 31388 23324 31444 23380
rect 31276 22876 31332 22932
rect 31612 23154 31668 23156
rect 31612 23102 31614 23154
rect 31614 23102 31666 23154
rect 31666 23102 31668 23154
rect 31612 23100 31668 23102
rect 31388 22370 31444 22372
rect 31388 22318 31390 22370
rect 31390 22318 31442 22370
rect 31442 22318 31444 22370
rect 31388 22316 31444 22318
rect 31164 21420 31220 21476
rect 31332 21532 31388 21588
rect 31164 21196 31220 21252
rect 31332 20972 31388 21028
rect 30940 20300 30996 20356
rect 31052 20188 31108 20244
rect 31276 19964 31332 20020
rect 31052 19180 31108 19236
rect 31164 19516 31220 19572
rect 30268 18732 30324 18788
rect 31388 19852 31444 19908
rect 31612 21586 31668 21588
rect 31612 21534 31614 21586
rect 31614 21534 31666 21586
rect 31666 21534 31668 21586
rect 31612 21532 31668 21534
rect 32508 25004 32564 25060
rect 34188 29986 34244 29988
rect 34188 29934 34190 29986
rect 34190 29934 34242 29986
rect 34242 29934 34244 29986
rect 34188 29932 34244 29934
rect 33846 29034 33902 29036
rect 33846 28982 33848 29034
rect 33848 28982 33900 29034
rect 33900 28982 33902 29034
rect 33846 28980 33902 28982
rect 33950 29034 34006 29036
rect 33950 28982 33952 29034
rect 33952 28982 34004 29034
rect 34004 28982 34006 29034
rect 33950 28980 34006 28982
rect 34054 29034 34110 29036
rect 34054 28982 34056 29034
rect 34056 28982 34108 29034
rect 34108 28982 34110 29034
rect 34054 28980 34110 28982
rect 33740 28476 33796 28532
rect 34188 27916 34244 27972
rect 34412 30828 34468 30884
rect 34412 29932 34468 29988
rect 34412 29148 34468 29204
rect 35084 34188 35140 34244
rect 35084 33404 35140 33460
rect 34748 30044 34804 30100
rect 35028 33180 35084 33236
rect 36148 36370 36204 36372
rect 36148 36318 36150 36370
rect 36150 36318 36202 36370
rect 36202 36318 36204 36370
rect 36148 36316 36204 36318
rect 35980 36204 36036 36260
rect 35644 34412 35700 34468
rect 35420 33852 35476 33908
rect 35644 33852 35700 33908
rect 35868 33404 35924 33460
rect 35420 32844 35476 32900
rect 35308 32562 35364 32564
rect 35308 32510 35310 32562
rect 35310 32510 35362 32562
rect 35362 32510 35364 32562
rect 35308 32508 35364 32510
rect 35196 31836 35252 31892
rect 35084 30882 35140 30884
rect 35084 30830 35086 30882
rect 35086 30830 35138 30882
rect 35138 30830 35140 30882
rect 35084 30828 35140 30830
rect 35644 32284 35700 32340
rect 35868 32956 35924 33012
rect 38332 37436 38388 37492
rect 37604 36988 37660 37044
rect 38332 36988 38388 37044
rect 36372 34802 36428 34804
rect 36372 34750 36374 34802
rect 36374 34750 36426 34802
rect 36426 34750 36428 34802
rect 36372 34748 36428 34750
rect 36204 34300 36260 34356
rect 36260 34130 36316 34132
rect 36260 34078 36262 34130
rect 36262 34078 36314 34130
rect 36314 34078 36316 34130
rect 36260 34076 36316 34078
rect 36372 33122 36428 33124
rect 36372 33070 36374 33122
rect 36374 33070 36426 33122
rect 36426 33070 36428 33122
rect 36372 33068 36428 33070
rect 36652 33068 36708 33124
rect 36540 32844 36596 32900
rect 38508 36090 38564 36092
rect 38508 36038 38510 36090
rect 38510 36038 38562 36090
rect 38562 36038 38564 36090
rect 38508 36036 38564 36038
rect 38612 36090 38668 36092
rect 38612 36038 38614 36090
rect 38614 36038 38666 36090
rect 38666 36038 38668 36090
rect 38612 36036 38668 36038
rect 38716 36090 38772 36092
rect 38716 36038 38718 36090
rect 38718 36038 38770 36090
rect 38770 36038 38772 36090
rect 38716 36036 38772 36038
rect 37996 35420 38052 35476
rect 37324 34018 37380 34020
rect 37324 33966 37326 34018
rect 37326 33966 37378 34018
rect 37378 33966 37380 34018
rect 37324 33964 37380 33966
rect 38508 34522 38564 34524
rect 38508 34470 38510 34522
rect 38510 34470 38562 34522
rect 38562 34470 38564 34522
rect 38508 34468 38564 34470
rect 38612 34522 38668 34524
rect 38612 34470 38614 34522
rect 38614 34470 38666 34522
rect 38666 34470 38668 34522
rect 38612 34468 38668 34470
rect 38716 34522 38772 34524
rect 38716 34470 38718 34522
rect 38718 34470 38770 34522
rect 38770 34470 38772 34522
rect 38716 34468 38772 34470
rect 36988 33234 37044 33236
rect 36988 33182 36990 33234
rect 36990 33182 37042 33234
rect 37042 33182 37044 33234
rect 36988 33180 37044 33182
rect 36876 32732 36932 32788
rect 36092 32450 36148 32452
rect 36092 32398 36094 32450
rect 36094 32398 36146 32450
rect 36146 32398 36148 32450
rect 36092 32396 36148 32398
rect 35868 32060 35924 32116
rect 35924 31890 35980 31892
rect 35924 31838 35926 31890
rect 35926 31838 35978 31890
rect 35978 31838 35980 31890
rect 35924 31836 35980 31838
rect 35756 31164 35812 31220
rect 36204 32060 36260 32116
rect 36652 32172 36708 32228
rect 34972 29148 35028 29204
rect 34860 28028 34916 28084
rect 33846 27466 33902 27468
rect 33846 27414 33848 27466
rect 33848 27414 33900 27466
rect 33900 27414 33902 27466
rect 33846 27412 33902 27414
rect 33950 27466 34006 27468
rect 33950 27414 33952 27466
rect 33952 27414 34004 27466
rect 34004 27414 34006 27466
rect 33950 27412 34006 27414
rect 34054 27466 34110 27468
rect 34054 27414 34056 27466
rect 34056 27414 34108 27466
rect 34108 27414 34110 27466
rect 34054 27412 34110 27414
rect 34412 27580 34468 27636
rect 33628 26012 33684 26068
rect 33516 25506 33572 25508
rect 33516 25454 33518 25506
rect 33518 25454 33570 25506
rect 33570 25454 33572 25506
rect 33516 25452 33572 25454
rect 33846 25898 33902 25900
rect 33846 25846 33848 25898
rect 33848 25846 33900 25898
rect 33900 25846 33902 25898
rect 33846 25844 33902 25846
rect 33950 25898 34006 25900
rect 33950 25846 33952 25898
rect 33952 25846 34004 25898
rect 34004 25846 34006 25898
rect 33950 25844 34006 25846
rect 34054 25898 34110 25900
rect 34054 25846 34056 25898
rect 34056 25846 34108 25898
rect 34108 25846 34110 25898
rect 34054 25844 34110 25846
rect 33852 25340 33908 25396
rect 34188 25228 34244 25284
rect 32732 24556 32788 24612
rect 31836 23938 31892 23940
rect 31836 23886 31838 23938
rect 31838 23886 31890 23938
rect 31890 23886 31892 23938
rect 31836 23884 31892 23886
rect 31948 23548 32004 23604
rect 31836 21980 31892 22036
rect 32060 22876 32116 22932
rect 31612 20018 31668 20020
rect 31612 19966 31614 20018
rect 31614 19966 31666 20018
rect 31666 19966 31668 20018
rect 31612 19964 31668 19966
rect 29484 18562 29540 18564
rect 29484 18510 29486 18562
rect 29486 18510 29538 18562
rect 29538 18510 29540 18562
rect 29484 18508 29540 18510
rect 30268 18508 30324 18564
rect 28028 18450 28084 18452
rect 28028 18398 28030 18450
rect 28030 18398 28082 18450
rect 28082 18398 28084 18450
rect 28028 18396 28084 18398
rect 29820 18450 29876 18452
rect 27804 17164 27860 17220
rect 27804 16940 27860 16996
rect 25340 14530 25396 14532
rect 25340 14478 25342 14530
rect 25342 14478 25394 14530
rect 25394 14478 25396 14530
rect 25340 14476 25396 14478
rect 25900 14588 25956 14644
rect 26404 14476 26460 14532
rect 24836 14418 24892 14420
rect 24836 14366 24838 14418
rect 24838 14366 24890 14418
rect 24890 14366 24892 14418
rect 24836 14364 24892 14366
rect 25788 14364 25844 14420
rect 27076 14642 27132 14644
rect 27076 14590 27078 14642
rect 27078 14590 27130 14642
rect 27130 14590 27132 14642
rect 27076 14588 27132 14590
rect 24332 13468 24388 13524
rect 24522 13354 24578 13356
rect 24522 13302 24524 13354
rect 24524 13302 24576 13354
rect 24576 13302 24578 13354
rect 24522 13300 24578 13302
rect 24626 13354 24682 13356
rect 24626 13302 24628 13354
rect 24628 13302 24680 13354
rect 24680 13302 24682 13354
rect 24626 13300 24682 13302
rect 24730 13354 24786 13356
rect 24730 13302 24732 13354
rect 24732 13302 24784 13354
rect 24784 13302 24786 13354
rect 24730 13300 24786 13302
rect 25340 13522 25396 13524
rect 25340 13470 25342 13522
rect 25342 13470 25394 13522
rect 25394 13470 25396 13522
rect 25340 13468 25396 13470
rect 24892 13244 24948 13300
rect 23212 11788 23268 11844
rect 22428 9826 22484 9828
rect 22428 9774 22430 9826
rect 22430 9774 22482 9826
rect 22482 9774 22484 9826
rect 22428 9772 22484 9774
rect 21980 9212 22036 9268
rect 23884 10108 23940 10164
rect 22764 9212 22820 9268
rect 21868 8428 21924 8484
rect 25116 12178 25172 12180
rect 25116 12126 25118 12178
rect 25118 12126 25170 12178
rect 25170 12126 25172 12178
rect 25116 12124 25172 12126
rect 27244 14140 27300 14196
rect 28644 17778 28700 17780
rect 28644 17726 28646 17778
rect 28646 17726 28698 17778
rect 28698 17726 28700 17778
rect 28644 17724 28700 17726
rect 28140 17500 28196 17556
rect 28588 16882 28644 16884
rect 28588 16830 28590 16882
rect 28590 16830 28642 16882
rect 28642 16830 28644 16882
rect 28588 16828 28644 16830
rect 29372 18172 29428 18228
rect 29820 18398 29822 18450
rect 29822 18398 29874 18450
rect 29874 18398 29876 18450
rect 29820 18396 29876 18398
rect 29372 17724 29428 17780
rect 29596 17724 29652 17780
rect 30268 18172 30324 18228
rect 29820 17666 29876 17668
rect 29820 17614 29822 17666
rect 29822 17614 29874 17666
rect 29874 17614 29876 17666
rect 29820 17612 29876 17614
rect 30098 17388 30154 17444
rect 29036 17164 29092 17220
rect 29184 17274 29240 17276
rect 29184 17222 29186 17274
rect 29186 17222 29238 17274
rect 29238 17222 29240 17274
rect 29184 17220 29240 17222
rect 29288 17274 29344 17276
rect 29288 17222 29290 17274
rect 29290 17222 29342 17274
rect 29342 17222 29344 17274
rect 29288 17220 29344 17222
rect 29392 17274 29448 17276
rect 29392 17222 29394 17274
rect 29394 17222 29446 17274
rect 29446 17222 29448 17274
rect 29392 17220 29448 17222
rect 29372 16828 29428 16884
rect 28588 16492 28644 16548
rect 28252 16380 28308 16436
rect 28364 16210 28420 16212
rect 28364 16158 28366 16210
rect 28366 16158 28418 16210
rect 28418 16158 28420 16210
rect 28364 16156 28420 16158
rect 28140 15314 28196 15316
rect 28140 15262 28142 15314
rect 28142 15262 28194 15314
rect 28194 15262 28196 15314
rect 28140 15260 28196 15262
rect 29036 16044 29092 16100
rect 29184 15706 29240 15708
rect 29184 15654 29186 15706
rect 29186 15654 29238 15706
rect 29238 15654 29240 15706
rect 29184 15652 29240 15654
rect 29288 15706 29344 15708
rect 29288 15654 29290 15706
rect 29290 15654 29342 15706
rect 29342 15654 29344 15706
rect 29288 15652 29344 15654
rect 29392 15706 29448 15708
rect 29392 15654 29394 15706
rect 29394 15654 29446 15706
rect 29446 15654 29448 15706
rect 29392 15652 29448 15654
rect 28588 15260 28644 15316
rect 27804 13020 27860 13076
rect 24522 11786 24578 11788
rect 24522 11734 24524 11786
rect 24524 11734 24576 11786
rect 24576 11734 24578 11786
rect 24522 11732 24578 11734
rect 24626 11786 24682 11788
rect 24626 11734 24628 11786
rect 24628 11734 24680 11786
rect 24680 11734 24682 11786
rect 24626 11732 24682 11734
rect 24730 11786 24786 11788
rect 24730 11734 24732 11786
rect 24732 11734 24784 11786
rect 24784 11734 24786 11786
rect 24730 11732 24786 11734
rect 25116 11676 25172 11732
rect 24522 10218 24578 10220
rect 24522 10166 24524 10218
rect 24524 10166 24576 10218
rect 24576 10166 24578 10218
rect 24522 10164 24578 10166
rect 24626 10218 24682 10220
rect 24626 10166 24628 10218
rect 24628 10166 24680 10218
rect 24680 10166 24682 10218
rect 24626 10164 24682 10166
rect 24730 10218 24786 10220
rect 24730 10166 24732 10218
rect 24732 10166 24784 10218
rect 24784 10166 24786 10218
rect 24730 10164 24786 10166
rect 24522 8650 24578 8652
rect 24522 8598 24524 8650
rect 24524 8598 24576 8650
rect 24576 8598 24578 8650
rect 24522 8596 24578 8598
rect 24626 8650 24682 8652
rect 24626 8598 24628 8650
rect 24628 8598 24680 8650
rect 24680 8598 24682 8650
rect 24626 8596 24682 8598
rect 24730 8650 24786 8652
rect 24730 8598 24732 8650
rect 24732 8598 24784 8650
rect 24784 8598 24786 8650
rect 24730 8596 24786 8598
rect 17108 7420 17164 7476
rect 17276 7474 17332 7476
rect 17276 7422 17278 7474
rect 17278 7422 17330 7474
rect 17330 7422 17332 7474
rect 17276 7420 17332 7422
rect 19012 6748 19068 6804
rect 18844 6690 18900 6692
rect 18844 6638 18846 6690
rect 18846 6638 18898 6690
rect 18898 6638 18900 6690
rect 18844 6636 18900 6638
rect 18060 6524 18116 6580
rect 16940 6412 16996 6468
rect 17948 6412 18004 6468
rect 16100 6076 16156 6132
rect 16492 6076 16548 6132
rect 16268 5234 16324 5236
rect 16268 5182 16270 5234
rect 16270 5182 16322 5234
rect 16322 5182 16324 5234
rect 16268 5180 16324 5182
rect 15260 4338 15316 4340
rect 15260 4286 15262 4338
rect 15262 4286 15314 4338
rect 15314 4286 15316 4338
rect 15260 4284 15316 4286
rect 15988 4338 16044 4340
rect 15988 4286 15990 4338
rect 15990 4286 16042 4338
rect 16042 4286 16044 4338
rect 15988 4284 16044 4286
rect 17500 6076 17556 6132
rect 17388 5628 17444 5684
rect 16734 4338 16790 4340
rect 16734 4286 16736 4338
rect 16736 4286 16788 4338
rect 16788 4286 16790 4338
rect 16734 4284 16790 4286
rect 15198 3946 15254 3948
rect 15198 3894 15200 3946
rect 15200 3894 15252 3946
rect 15252 3894 15254 3946
rect 15198 3892 15254 3894
rect 15302 3946 15358 3948
rect 15302 3894 15304 3946
rect 15304 3894 15356 3946
rect 15356 3894 15358 3946
rect 15302 3892 15358 3894
rect 15406 3946 15462 3948
rect 15406 3894 15408 3946
rect 15408 3894 15460 3946
rect 15460 3894 15462 3946
rect 15406 3892 15462 3894
rect 14588 3500 14644 3556
rect 17444 4450 17500 4452
rect 17444 4398 17446 4450
rect 17446 4398 17498 4450
rect 17498 4398 17500 4450
rect 17444 4396 17500 4398
rect 17724 4338 17780 4340
rect 17724 4286 17726 4338
rect 17726 4286 17778 4338
rect 17778 4286 17780 4338
rect 17724 4284 17780 4286
rect 19012 6524 19068 6580
rect 19180 6636 19236 6692
rect 18172 6076 18228 6132
rect 19516 6524 19572 6580
rect 19180 5964 19236 6020
rect 18508 5682 18564 5684
rect 18508 5630 18510 5682
rect 18510 5630 18562 5682
rect 18562 5630 18564 5682
rect 18508 5628 18564 5630
rect 19860 7866 19916 7868
rect 19860 7814 19862 7866
rect 19862 7814 19914 7866
rect 19914 7814 19916 7866
rect 19860 7812 19916 7814
rect 19964 7866 20020 7868
rect 19964 7814 19966 7866
rect 19966 7814 20018 7866
rect 20018 7814 20020 7866
rect 19964 7812 20020 7814
rect 20068 7866 20124 7868
rect 20068 7814 20070 7866
rect 20070 7814 20122 7866
rect 20122 7814 20124 7866
rect 20068 7812 20124 7814
rect 21756 8204 21812 8260
rect 19964 6748 20020 6804
rect 19758 6690 19814 6692
rect 19758 6638 19760 6690
rect 19760 6638 19812 6690
rect 19812 6638 19814 6690
rect 19758 6636 19814 6638
rect 20076 6412 20132 6468
rect 20300 6690 20356 6692
rect 20300 6638 20302 6690
rect 20302 6638 20354 6690
rect 20354 6638 20356 6690
rect 20300 6636 20356 6638
rect 20300 6412 20356 6468
rect 19860 6298 19916 6300
rect 19860 6246 19862 6298
rect 19862 6246 19914 6298
rect 19914 6246 19916 6298
rect 19860 6244 19916 6246
rect 19964 6298 20020 6300
rect 19964 6246 19966 6298
rect 19966 6246 20018 6298
rect 20018 6246 20020 6298
rect 19964 6244 20020 6246
rect 20068 6298 20124 6300
rect 20068 6246 20070 6298
rect 20070 6246 20122 6298
rect 20122 6246 20124 6298
rect 20068 6244 20124 6246
rect 19628 5180 19684 5236
rect 18788 4956 18844 5012
rect 19860 4730 19916 4732
rect 19860 4678 19862 4730
rect 19862 4678 19914 4730
rect 19914 4678 19916 4730
rect 19860 4676 19916 4678
rect 19964 4730 20020 4732
rect 19964 4678 19966 4730
rect 19966 4678 20018 4730
rect 20018 4678 20020 4730
rect 19964 4676 20020 4678
rect 20068 4730 20124 4732
rect 20068 4678 20070 4730
rect 20070 4678 20122 4730
rect 20122 4678 20124 4730
rect 20068 4676 20124 4678
rect 20972 3724 21028 3780
rect 21084 6524 21140 6580
rect 20860 3612 20916 3668
rect 19860 3162 19916 3164
rect 19860 3110 19862 3162
rect 19862 3110 19914 3162
rect 19914 3110 19916 3162
rect 19860 3108 19916 3110
rect 19964 3162 20020 3164
rect 19964 3110 19966 3162
rect 19966 3110 20018 3162
rect 20018 3110 20020 3162
rect 19964 3108 20020 3110
rect 20068 3162 20124 3164
rect 20068 3110 20070 3162
rect 20070 3110 20122 3162
rect 20122 3110 20124 3162
rect 20068 3108 20124 3110
rect 21420 6466 21476 6468
rect 21420 6414 21422 6466
rect 21422 6414 21474 6466
rect 21474 6414 21476 6466
rect 21420 6412 21476 6414
rect 25900 11116 25956 11172
rect 26012 10780 26068 10836
rect 26348 10780 26404 10836
rect 26908 11170 26964 11172
rect 26908 11118 26910 11170
rect 26910 11118 26962 11170
rect 26962 11118 26964 11170
rect 26908 11116 26964 11118
rect 26012 10108 26068 10164
rect 25676 9996 25732 10052
rect 25116 9826 25172 9828
rect 25116 9774 25118 9826
rect 25118 9774 25170 9826
rect 25170 9774 25172 9826
rect 25116 9772 25172 9774
rect 24892 8428 24948 8484
rect 26124 9826 26180 9828
rect 26124 9774 26126 9826
rect 26126 9774 26178 9826
rect 26178 9774 26180 9826
rect 26124 9772 26180 9774
rect 25994 8818 26050 8820
rect 25994 8766 25996 8818
rect 25996 8766 26048 8818
rect 26048 8766 26050 8818
rect 25994 8764 26050 8766
rect 26796 9714 26852 9716
rect 26796 9662 26798 9714
rect 26798 9662 26850 9714
rect 26850 9662 26852 9714
rect 26796 9660 26852 9662
rect 26460 9100 26516 9156
rect 22204 8258 22260 8260
rect 22204 8206 22206 8258
rect 22206 8206 22258 8258
rect 22258 8206 22260 8258
rect 22204 8204 22260 8206
rect 21420 6018 21476 6020
rect 21420 5966 21422 6018
rect 21422 5966 21474 6018
rect 21474 5966 21476 6018
rect 21420 5964 21476 5966
rect 21756 5964 21812 6020
rect 22092 5964 22148 6020
rect 23324 7644 23380 7700
rect 22876 6636 22932 6692
rect 22764 5906 22820 5908
rect 22764 5854 22766 5906
rect 22766 5854 22818 5906
rect 22818 5854 22820 5906
rect 22764 5852 22820 5854
rect 23996 6690 24052 6692
rect 23996 6638 23998 6690
rect 23998 6638 24050 6690
rect 24050 6638 24052 6690
rect 23996 6636 24052 6638
rect 23772 5740 23828 5796
rect 24108 5740 24164 5796
rect 23156 5068 23212 5124
rect 23660 5122 23716 5124
rect 23660 5070 23662 5122
rect 23662 5070 23714 5122
rect 23714 5070 23716 5122
rect 23660 5068 23716 5070
rect 22540 4284 22596 4340
rect 23660 4338 23716 4340
rect 23660 4286 23662 4338
rect 23662 4286 23714 4338
rect 23714 4286 23716 4338
rect 23660 4284 23716 4286
rect 21196 3724 21252 3780
rect 22092 3666 22148 3668
rect 22092 3614 22094 3666
rect 22094 3614 22146 3666
rect 22146 3614 22148 3666
rect 22092 3612 22148 3614
rect 22652 3612 22708 3668
rect 24556 7474 24612 7476
rect 24556 7422 24558 7474
rect 24558 7422 24610 7474
rect 24610 7422 24612 7474
rect 24556 7420 24612 7422
rect 24522 7082 24578 7084
rect 24522 7030 24524 7082
rect 24524 7030 24576 7082
rect 24576 7030 24578 7082
rect 24522 7028 24578 7030
rect 24626 7082 24682 7084
rect 24626 7030 24628 7082
rect 24628 7030 24680 7082
rect 24680 7030 24682 7082
rect 24626 7028 24682 7030
rect 24730 7082 24786 7084
rect 24730 7030 24732 7082
rect 24732 7030 24784 7082
rect 24784 7030 24786 7082
rect 24730 7028 24786 7030
rect 24332 5906 24388 5908
rect 24332 5854 24334 5906
rect 24334 5854 24386 5906
rect 24386 5854 24388 5906
rect 24332 5852 24388 5854
rect 24332 5628 24388 5684
rect 24522 5514 24578 5516
rect 24522 5462 24524 5514
rect 24524 5462 24576 5514
rect 24576 5462 24578 5514
rect 24522 5460 24578 5462
rect 24626 5514 24682 5516
rect 24626 5462 24628 5514
rect 24628 5462 24680 5514
rect 24680 5462 24682 5514
rect 24626 5460 24682 5462
rect 24730 5514 24786 5516
rect 24730 5462 24732 5514
rect 24732 5462 24784 5514
rect 24784 5462 24786 5514
rect 24730 5460 24786 5462
rect 29316 14642 29372 14644
rect 29316 14590 29318 14642
rect 29318 14590 29370 14642
rect 29370 14590 29372 14642
rect 29316 14588 29372 14590
rect 28812 14140 28868 14196
rect 29184 14138 29240 14140
rect 29184 14086 29186 14138
rect 29186 14086 29238 14138
rect 29238 14086 29240 14138
rect 29184 14084 29240 14086
rect 29288 14138 29344 14140
rect 29288 14086 29290 14138
rect 29290 14086 29342 14138
rect 29342 14086 29344 14138
rect 29288 14084 29344 14086
rect 29392 14138 29448 14140
rect 29392 14086 29394 14138
rect 29394 14086 29446 14138
rect 29446 14086 29448 14138
rect 29392 14084 29448 14086
rect 30380 16828 30436 16884
rect 30492 16940 30548 16996
rect 30156 16604 30212 16660
rect 29708 13916 29764 13972
rect 29820 16492 29876 16548
rect 29932 16156 29988 16212
rect 30380 16156 30436 16212
rect 31164 18732 31220 18788
rect 32284 22876 32340 22932
rect 32172 22482 32228 22484
rect 32172 22430 32174 22482
rect 32174 22430 32226 22482
rect 32226 22430 32228 22482
rect 32172 22428 32228 22430
rect 32172 22092 32228 22148
rect 32396 22764 32452 22820
rect 32508 22540 32564 22596
rect 32284 21980 32340 22036
rect 32396 22316 32452 22372
rect 32284 21586 32340 21588
rect 32284 21534 32286 21586
rect 32286 21534 32338 21586
rect 32338 21534 32340 21586
rect 32284 21532 32340 21534
rect 32732 22764 32788 22820
rect 32844 23548 32900 23604
rect 33404 24780 33460 24836
rect 32956 23436 33012 23492
rect 33846 24330 33902 24332
rect 33846 24278 33848 24330
rect 33848 24278 33900 24330
rect 33900 24278 33902 24330
rect 33846 24276 33902 24278
rect 33950 24330 34006 24332
rect 33950 24278 33952 24330
rect 33952 24278 34004 24330
rect 34004 24278 34006 24330
rect 33950 24276 34006 24278
rect 34054 24330 34110 24332
rect 34054 24278 34056 24330
rect 34056 24278 34108 24330
rect 34108 24278 34110 24330
rect 34054 24276 34110 24278
rect 33846 22762 33902 22764
rect 33846 22710 33848 22762
rect 33848 22710 33900 22762
rect 33900 22710 33902 22762
rect 33846 22708 33902 22710
rect 33950 22762 34006 22764
rect 33950 22710 33952 22762
rect 33952 22710 34004 22762
rect 34004 22710 34006 22762
rect 33950 22708 34006 22710
rect 34054 22762 34110 22764
rect 34054 22710 34056 22762
rect 34056 22710 34108 22762
rect 34108 22710 34110 22762
rect 34054 22708 34110 22710
rect 34412 25676 34468 25732
rect 34692 25340 34748 25396
rect 36036 30322 36092 30324
rect 36036 30270 36038 30322
rect 36038 30270 36090 30322
rect 36090 30270 36092 30322
rect 36036 30268 36092 30270
rect 36316 29708 36372 29764
rect 36540 32060 36596 32116
rect 36540 30268 36596 30324
rect 36484 27074 36540 27076
rect 36484 27022 36486 27074
rect 36486 27022 36538 27074
rect 36538 27022 36540 27074
rect 36484 27020 36540 27022
rect 37156 31388 37212 31444
rect 37996 33906 38052 33908
rect 37996 33854 37998 33906
rect 37998 33854 38050 33906
rect 38050 33854 38052 33906
rect 37996 33852 38052 33854
rect 37660 33346 37716 33348
rect 37660 33294 37662 33346
rect 37662 33294 37714 33346
rect 37714 33294 37716 33346
rect 37660 33292 37716 33294
rect 38220 33292 38276 33348
rect 38108 33180 38164 33236
rect 37436 31612 37492 31668
rect 36988 30994 37044 30996
rect 36988 30942 36990 30994
rect 36990 30942 37042 30994
rect 37042 30942 37044 30994
rect 36988 30940 37044 30942
rect 37212 31164 37268 31220
rect 37324 31052 37380 31108
rect 37156 30210 37212 30212
rect 37156 30158 37158 30210
rect 37158 30158 37210 30210
rect 37210 30158 37212 30210
rect 37156 30156 37212 30158
rect 36764 29202 36820 29204
rect 36764 29150 36766 29202
rect 36766 29150 36818 29202
rect 36818 29150 36820 29202
rect 36764 29148 36820 29150
rect 36988 28700 37044 28756
rect 37436 28588 37492 28644
rect 37660 32396 37716 32452
rect 37996 32450 38052 32452
rect 37996 32398 37998 32450
rect 37998 32398 38050 32450
rect 38050 32398 38052 32450
rect 37996 32396 38052 32398
rect 37660 31052 37716 31108
rect 37660 30882 37716 30884
rect 37660 30830 37662 30882
rect 37662 30830 37714 30882
rect 37714 30830 37716 30882
rect 37660 30828 37716 30830
rect 37660 29932 37716 29988
rect 37902 30098 37958 30100
rect 37902 30046 37904 30098
rect 37904 30046 37956 30098
rect 37956 30046 37958 30098
rect 37902 30044 37958 30046
rect 38220 30940 38276 30996
rect 39004 33852 39060 33908
rect 38508 32954 38564 32956
rect 38508 32902 38510 32954
rect 38510 32902 38562 32954
rect 38562 32902 38564 32954
rect 38508 32900 38564 32902
rect 38612 32954 38668 32956
rect 38612 32902 38614 32954
rect 38614 32902 38666 32954
rect 38666 32902 38668 32954
rect 38612 32900 38668 32902
rect 38716 32954 38772 32956
rect 38716 32902 38718 32954
rect 38718 32902 38770 32954
rect 38770 32902 38772 32954
rect 38716 32900 38772 32902
rect 38508 31386 38564 31388
rect 38508 31334 38510 31386
rect 38510 31334 38562 31386
rect 38562 31334 38564 31386
rect 38508 31332 38564 31334
rect 38612 31386 38668 31388
rect 38612 31334 38614 31386
rect 38614 31334 38666 31386
rect 38666 31334 38668 31386
rect 38612 31332 38668 31334
rect 38716 31386 38772 31388
rect 38716 31334 38718 31386
rect 38718 31334 38770 31386
rect 38770 31334 38772 31386
rect 38716 31332 38772 31334
rect 38508 29818 38564 29820
rect 38508 29766 38510 29818
rect 38510 29766 38562 29818
rect 38562 29766 38564 29818
rect 38508 29764 38564 29766
rect 38612 29818 38668 29820
rect 38612 29766 38614 29818
rect 38614 29766 38666 29818
rect 38666 29766 38668 29818
rect 38612 29764 38668 29766
rect 38716 29818 38772 29820
rect 38716 29766 38718 29818
rect 38718 29766 38770 29818
rect 38770 29766 38772 29818
rect 38716 29764 38772 29766
rect 38332 29372 38388 29428
rect 38508 28250 38564 28252
rect 38508 28198 38510 28250
rect 38510 28198 38562 28250
rect 38562 28198 38564 28250
rect 38508 28196 38564 28198
rect 38612 28250 38668 28252
rect 38612 28198 38614 28250
rect 38614 28198 38666 28250
rect 38666 28198 38668 28250
rect 38612 28196 38668 28198
rect 38716 28250 38772 28252
rect 38716 28198 38718 28250
rect 38718 28198 38770 28250
rect 38770 28198 38772 28250
rect 38716 28196 38772 28198
rect 36876 26908 36932 26964
rect 35756 25506 35812 25508
rect 35756 25454 35758 25506
rect 35758 25454 35810 25506
rect 35810 25454 35812 25506
rect 35756 25452 35812 25454
rect 35364 25340 35420 25396
rect 35532 25394 35588 25396
rect 35532 25342 35534 25394
rect 35534 25342 35586 25394
rect 35586 25342 35588 25394
rect 35532 25340 35588 25342
rect 37996 26962 38052 26964
rect 37996 26910 37998 26962
rect 37998 26910 38050 26962
rect 38050 26910 38052 26962
rect 37996 26908 38052 26910
rect 35980 25004 36036 25060
rect 34972 24722 35028 24724
rect 34972 24670 34974 24722
rect 34974 24670 35026 24722
rect 35026 24670 35028 24722
rect 34972 24668 35028 24670
rect 35196 24780 35252 24836
rect 34580 24108 34636 24164
rect 34972 23772 35028 23828
rect 36876 24780 36932 24836
rect 37212 24722 37268 24724
rect 37212 24670 37214 24722
rect 37214 24670 37266 24722
rect 37266 24670 37268 24722
rect 37212 24668 37268 24670
rect 37436 24668 37492 24724
rect 36204 24556 36260 24612
rect 35308 24108 35364 24164
rect 35420 23996 35476 24052
rect 35196 23548 35252 23604
rect 34860 23324 34916 23380
rect 35644 23996 35700 24052
rect 35980 23938 36036 23940
rect 35980 23886 35982 23938
rect 35982 23886 36034 23938
rect 36034 23886 36036 23938
rect 35980 23884 36036 23886
rect 34524 23154 34580 23156
rect 34524 23102 34526 23154
rect 34526 23102 34578 23154
rect 34578 23102 34580 23154
rect 34524 23100 34580 23102
rect 35420 23154 35476 23156
rect 35420 23102 35422 23154
rect 35422 23102 35474 23154
rect 35474 23102 35476 23154
rect 35420 23100 35476 23102
rect 34860 22930 34916 22932
rect 34860 22878 34862 22930
rect 34862 22878 34914 22930
rect 34914 22878 34916 22930
rect 34860 22876 34916 22878
rect 33516 22540 33572 22596
rect 33404 22428 33460 22484
rect 32732 21756 32788 21812
rect 33740 22316 33796 22372
rect 32620 21532 32676 21588
rect 33516 21308 33572 21364
rect 33964 22204 34020 22260
rect 34636 22370 34692 22372
rect 34636 22318 34638 22370
rect 34638 22318 34690 22370
rect 34690 22318 34692 22370
rect 34636 22316 34692 22318
rect 34318 22258 34374 22260
rect 34318 22206 34320 22258
rect 34320 22206 34372 22258
rect 34372 22206 34374 22258
rect 34318 22204 34374 22206
rect 33846 21194 33902 21196
rect 33846 21142 33848 21194
rect 33848 21142 33900 21194
rect 33900 21142 33902 21194
rect 33846 21140 33902 21142
rect 33950 21194 34006 21196
rect 33950 21142 33952 21194
rect 33952 21142 34004 21194
rect 34004 21142 34006 21194
rect 33950 21140 34006 21142
rect 34054 21194 34110 21196
rect 34054 21142 34056 21194
rect 34056 21142 34108 21194
rect 34108 21142 34110 21194
rect 34054 21140 34110 21142
rect 35868 23548 35924 23604
rect 36372 23938 36428 23940
rect 36372 23886 36374 23938
rect 36374 23886 36426 23938
rect 36426 23886 36428 23938
rect 36372 23884 36428 23886
rect 37324 23938 37380 23940
rect 37324 23886 37326 23938
rect 37326 23886 37378 23938
rect 37378 23886 37380 23938
rect 37324 23884 37380 23886
rect 37548 24610 37604 24612
rect 37548 24558 37550 24610
rect 37550 24558 37602 24610
rect 37602 24558 37604 24610
rect 37548 24556 37604 24558
rect 37884 24780 37940 24836
rect 37996 24556 38052 24612
rect 37996 24108 38052 24164
rect 37436 23772 37492 23828
rect 35644 22876 35700 22932
rect 34972 21308 35028 21364
rect 34860 21084 34916 21140
rect 35644 21084 35700 21140
rect 33852 20802 33908 20804
rect 33852 20750 33854 20802
rect 33854 20750 33906 20802
rect 33906 20750 33908 20802
rect 33852 20748 33908 20750
rect 32564 20300 32620 20356
rect 34206 20300 34262 20356
rect 32060 19852 32116 19908
rect 31892 19628 31948 19684
rect 31164 18172 31220 18228
rect 31108 17778 31164 17780
rect 31108 17726 31110 17778
rect 31110 17726 31162 17778
rect 31162 17726 31164 17778
rect 31108 17724 31164 17726
rect 31108 16940 31164 16996
rect 30716 16492 30772 16548
rect 30828 16380 30884 16436
rect 31388 16210 31444 16212
rect 31388 16158 31390 16210
rect 31390 16158 31442 16210
rect 31442 16158 31444 16210
rect 31388 16156 31444 16158
rect 30994 16098 31050 16100
rect 30994 16046 30996 16098
rect 30996 16046 31048 16098
rect 31048 16046 31050 16098
rect 30994 16044 31050 16046
rect 29932 13468 29988 13524
rect 28588 12236 28644 12292
rect 28084 11506 28140 11508
rect 28084 11454 28086 11506
rect 28086 11454 28138 11506
rect 28138 11454 28140 11506
rect 28084 11452 28140 11454
rect 29596 12962 29652 12964
rect 29596 12910 29598 12962
rect 29598 12910 29650 12962
rect 29650 12910 29652 12962
rect 29596 12908 29652 12910
rect 30156 13356 30212 13412
rect 29184 12570 29240 12572
rect 29184 12518 29186 12570
rect 29186 12518 29238 12570
rect 29238 12518 29240 12570
rect 29184 12516 29240 12518
rect 29288 12570 29344 12572
rect 29288 12518 29290 12570
rect 29290 12518 29342 12570
rect 29342 12518 29344 12570
rect 29288 12516 29344 12518
rect 29392 12570 29448 12572
rect 29392 12518 29394 12570
rect 29394 12518 29446 12570
rect 29446 12518 29448 12570
rect 29392 12516 29448 12518
rect 28700 11676 28756 11732
rect 30660 13634 30716 13636
rect 30660 13582 30662 13634
rect 30662 13582 30714 13634
rect 30714 13582 30716 13634
rect 30660 13580 30716 13582
rect 31388 15484 31444 15540
rect 31500 15426 31556 15428
rect 31500 15374 31502 15426
rect 31502 15374 31554 15426
rect 31554 15374 31556 15426
rect 31500 15372 31556 15374
rect 30996 13522 31052 13524
rect 30996 13470 30998 13522
rect 30998 13470 31050 13522
rect 31050 13470 31052 13522
rect 30996 13468 31052 13470
rect 31164 13468 31220 13524
rect 30492 12348 30548 12404
rect 31388 13580 31444 13636
rect 31724 16828 31780 16884
rect 31836 19068 31892 19124
rect 31724 16604 31780 16660
rect 34636 19852 34692 19908
rect 32340 19628 32396 19684
rect 33846 19626 33902 19628
rect 33846 19574 33848 19626
rect 33848 19574 33900 19626
rect 33900 19574 33902 19626
rect 33846 19572 33902 19574
rect 33950 19626 34006 19628
rect 33950 19574 33952 19626
rect 33952 19574 34004 19626
rect 34004 19574 34006 19626
rect 33950 19572 34006 19574
rect 34054 19626 34110 19628
rect 34054 19574 34056 19626
rect 34056 19574 34108 19626
rect 34108 19574 34110 19626
rect 34054 19572 34110 19574
rect 32060 17724 32116 17780
rect 32172 16828 32228 16884
rect 32004 16604 32060 16660
rect 32004 16380 32060 16436
rect 31836 15484 31892 15540
rect 31724 15372 31780 15428
rect 31612 13692 31668 13748
rect 31612 13468 31668 13524
rect 31500 13356 31556 13412
rect 31276 13244 31332 13300
rect 29372 11676 29428 11732
rect 28588 11452 28644 11508
rect 29184 11002 29240 11004
rect 29184 10950 29186 11002
rect 29186 10950 29238 11002
rect 29238 10950 29240 11002
rect 29184 10948 29240 10950
rect 29288 11002 29344 11004
rect 29288 10950 29290 11002
rect 29290 10950 29342 11002
rect 29342 10950 29344 11002
rect 29288 10948 29344 10950
rect 29392 11002 29448 11004
rect 29392 10950 29394 11002
rect 29394 10950 29446 11002
rect 29446 10950 29448 11002
rect 29392 10948 29448 10950
rect 30492 11170 30548 11172
rect 30492 11118 30494 11170
rect 30494 11118 30546 11170
rect 30546 11118 30548 11170
rect 30492 11116 30548 11118
rect 27916 9996 27972 10052
rect 27132 9548 27188 9604
rect 27804 9100 27860 9156
rect 28122 9042 28178 9044
rect 28122 8990 28124 9042
rect 28124 8990 28176 9042
rect 28176 8990 28178 9042
rect 28122 8988 28178 8990
rect 28364 9772 28420 9828
rect 28364 9212 28420 9268
rect 27020 8764 27076 8820
rect 26908 8316 26964 8372
rect 25434 7644 25490 7700
rect 25676 7474 25732 7476
rect 25676 7422 25678 7474
rect 25678 7422 25730 7474
rect 25730 7422 25732 7474
rect 26348 7586 26404 7588
rect 26348 7534 26350 7586
rect 26350 7534 26402 7586
rect 26402 7534 26404 7586
rect 26348 7532 26404 7534
rect 25676 7420 25732 7422
rect 26852 7308 26908 7364
rect 27020 6860 27076 6916
rect 25228 5964 25284 6020
rect 25788 5740 25844 5796
rect 24444 4338 24500 4340
rect 24444 4286 24446 4338
rect 24446 4286 24498 4338
rect 24498 4286 24500 4338
rect 24444 4284 24500 4286
rect 26236 5682 26292 5684
rect 26236 5630 26238 5682
rect 26238 5630 26290 5682
rect 26290 5630 26292 5682
rect 26236 5628 26292 5630
rect 26236 4844 26292 4900
rect 26908 4338 26964 4340
rect 26908 4286 26910 4338
rect 26910 4286 26962 4338
rect 26962 4286 26964 4338
rect 26908 4284 26964 4286
rect 24522 3946 24578 3948
rect 24522 3894 24524 3946
rect 24524 3894 24576 3946
rect 24576 3894 24578 3946
rect 24522 3892 24578 3894
rect 24626 3946 24682 3948
rect 24626 3894 24628 3946
rect 24628 3894 24680 3946
rect 24680 3894 24682 3946
rect 24626 3892 24682 3894
rect 24730 3946 24786 3948
rect 24730 3894 24732 3946
rect 24732 3894 24784 3946
rect 24784 3894 24786 3946
rect 24730 3892 24786 3894
rect 24556 3724 24612 3780
rect 27468 8316 27524 8372
rect 27356 7474 27412 7476
rect 27356 7422 27358 7474
rect 27358 7422 27410 7474
rect 27410 7422 27412 7474
rect 27356 7420 27412 7422
rect 29036 10108 29092 10164
rect 29260 10332 29316 10388
rect 29148 9772 29204 9828
rect 29708 10332 29764 10388
rect 29184 9434 29240 9436
rect 29184 9382 29186 9434
rect 29186 9382 29238 9434
rect 29238 9382 29240 9434
rect 29184 9380 29240 9382
rect 29288 9434 29344 9436
rect 29288 9382 29290 9434
rect 29290 9382 29342 9434
rect 29342 9382 29344 9434
rect 29288 9380 29344 9382
rect 29392 9434 29448 9436
rect 29392 9382 29394 9434
rect 29394 9382 29446 9434
rect 29446 9382 29448 9434
rect 29392 9380 29448 9382
rect 30604 10332 30660 10388
rect 30828 12962 30884 12964
rect 30828 12910 30830 12962
rect 30830 12910 30882 12962
rect 30882 12910 30884 12962
rect 30828 12908 30884 12910
rect 32844 16828 32900 16884
rect 33846 18058 33902 18060
rect 33846 18006 33848 18058
rect 33848 18006 33900 18058
rect 33900 18006 33902 18058
rect 33846 18004 33902 18006
rect 33950 18058 34006 18060
rect 33950 18006 33952 18058
rect 33952 18006 34004 18058
rect 34004 18006 34006 18058
rect 33950 18004 34006 18006
rect 34054 18058 34110 18060
rect 34054 18006 34056 18058
rect 34056 18006 34108 18058
rect 34108 18006 34110 18058
rect 34054 18004 34110 18006
rect 34468 18450 34524 18452
rect 34468 18398 34470 18450
rect 34470 18398 34522 18450
rect 34522 18398 34524 18450
rect 34468 18396 34524 18398
rect 34412 18172 34468 18228
rect 34188 17276 34244 17332
rect 34076 16770 34132 16772
rect 34076 16718 34078 16770
rect 34078 16718 34130 16770
rect 34130 16718 34132 16770
rect 34076 16716 34132 16718
rect 33846 16490 33902 16492
rect 33846 16438 33848 16490
rect 33848 16438 33900 16490
rect 33900 16438 33902 16490
rect 33846 16436 33902 16438
rect 33950 16490 34006 16492
rect 33950 16438 33952 16490
rect 33952 16438 34004 16490
rect 34004 16438 34006 16490
rect 33950 16436 34006 16438
rect 34054 16490 34110 16492
rect 34054 16438 34056 16490
rect 34056 16438 34108 16490
rect 34108 16438 34110 16490
rect 34054 16436 34110 16438
rect 35252 19906 35308 19908
rect 35252 19854 35254 19906
rect 35254 19854 35306 19906
rect 35306 19854 35308 19906
rect 35252 19852 35308 19854
rect 37156 23436 37212 23492
rect 37996 23548 38052 23604
rect 35980 20300 36036 20356
rect 34748 18450 34804 18452
rect 34748 18398 34750 18450
rect 34750 18398 34802 18450
rect 34802 18398 34804 18450
rect 34748 18396 34804 18398
rect 35084 18226 35140 18228
rect 35084 18174 35086 18226
rect 35086 18174 35138 18226
rect 35138 18174 35140 18226
rect 35084 18172 35140 18174
rect 36988 20860 37044 20916
rect 37156 20802 37212 20804
rect 37156 20750 37158 20802
rect 37158 20750 37210 20802
rect 37210 20750 37212 20802
rect 37156 20748 37212 20750
rect 36428 19852 36484 19908
rect 36428 19404 36484 19460
rect 37156 19404 37212 19460
rect 35084 17276 35140 17332
rect 35308 16770 35364 16772
rect 35308 16718 35310 16770
rect 35310 16718 35362 16770
rect 35362 16718 35364 16770
rect 35308 16716 35364 16718
rect 33516 16268 33572 16324
rect 33180 15874 33236 15876
rect 33180 15822 33182 15874
rect 33182 15822 33234 15874
rect 33234 15822 33236 15874
rect 33180 15820 33236 15822
rect 32956 15036 33012 15092
rect 34412 16268 34468 16324
rect 33852 15820 33908 15876
rect 33852 15148 33908 15204
rect 33628 15036 33684 15092
rect 31948 13020 32004 13076
rect 32060 13244 32116 13300
rect 31612 12684 31668 12740
rect 31164 11116 31220 11172
rect 29932 10108 29988 10164
rect 28588 8204 28644 8260
rect 28588 7532 28644 7588
rect 27468 7308 27524 7364
rect 27580 5964 27636 6020
rect 27468 5234 27524 5236
rect 27468 5182 27470 5234
rect 27470 5182 27522 5234
rect 27522 5182 27524 5234
rect 27468 5180 27524 5182
rect 28364 6636 28420 6692
rect 28122 5906 28178 5908
rect 28122 5854 28124 5906
rect 28124 5854 28176 5906
rect 28176 5854 28178 5906
rect 28122 5852 28178 5854
rect 28364 5906 28420 5908
rect 28364 5854 28366 5906
rect 28366 5854 28418 5906
rect 28418 5854 28420 5906
rect 28364 5852 28420 5854
rect 29036 8258 29092 8260
rect 29036 8206 29038 8258
rect 29038 8206 29090 8258
rect 29090 8206 29092 8258
rect 29036 8204 29092 8206
rect 29184 7866 29240 7868
rect 29184 7814 29186 7866
rect 29186 7814 29238 7866
rect 29238 7814 29240 7866
rect 29184 7812 29240 7814
rect 29288 7866 29344 7868
rect 29288 7814 29290 7866
rect 29290 7814 29342 7866
rect 29342 7814 29344 7866
rect 29288 7812 29344 7814
rect 29392 7866 29448 7868
rect 29392 7814 29394 7866
rect 29394 7814 29446 7866
rect 29446 7814 29448 7866
rect 29392 7812 29448 7814
rect 29036 7586 29092 7588
rect 29036 7534 29038 7586
rect 29038 7534 29090 7586
rect 29090 7534 29092 7586
rect 29036 7532 29092 7534
rect 29484 6860 29540 6916
rect 28700 6076 28756 6132
rect 29596 6412 29652 6468
rect 29184 6298 29240 6300
rect 29184 6246 29186 6298
rect 29186 6246 29238 6298
rect 29238 6246 29240 6298
rect 29184 6244 29240 6246
rect 29288 6298 29344 6300
rect 29288 6246 29290 6298
rect 29290 6246 29342 6298
rect 29342 6246 29344 6298
rect 29288 6244 29344 6246
rect 29392 6298 29448 6300
rect 29392 6246 29394 6298
rect 29394 6246 29446 6298
rect 29446 6246 29448 6298
rect 29392 6244 29448 6246
rect 28868 5964 28924 6020
rect 28364 5180 28420 5236
rect 27916 5068 27972 5124
rect 29184 4730 29240 4732
rect 29184 4678 29186 4730
rect 29186 4678 29238 4730
rect 29238 4678 29240 4730
rect 29184 4676 29240 4678
rect 29288 4730 29344 4732
rect 29288 4678 29290 4730
rect 29290 4678 29342 4730
rect 29342 4678 29344 4730
rect 29288 4676 29344 4678
rect 29392 4730 29448 4732
rect 29392 4678 29394 4730
rect 29394 4678 29446 4730
rect 29446 4678 29448 4730
rect 29392 4676 29448 4678
rect 29820 6524 29876 6580
rect 29708 6300 29764 6356
rect 30380 9548 30436 9604
rect 30380 9154 30436 9156
rect 30380 9102 30382 9154
rect 30382 9102 30434 9154
rect 30434 9102 30436 9154
rect 30380 9100 30436 9102
rect 30212 9042 30268 9044
rect 30212 8990 30214 9042
rect 30214 8990 30266 9042
rect 30266 8990 30268 9042
rect 30212 8988 30268 8990
rect 30716 9042 30772 9044
rect 30716 8990 30718 9042
rect 30718 8990 30770 9042
rect 30770 8990 30772 9042
rect 30716 8988 30772 8990
rect 31500 9100 31556 9156
rect 34020 15036 34076 15092
rect 33846 14922 33902 14924
rect 33846 14870 33848 14922
rect 33848 14870 33900 14922
rect 33900 14870 33902 14922
rect 33846 14868 33902 14870
rect 33950 14922 34006 14924
rect 33950 14870 33952 14922
rect 33952 14870 34004 14922
rect 34004 14870 34006 14922
rect 33950 14868 34006 14870
rect 34054 14922 34110 14924
rect 34054 14870 34056 14922
rect 34056 14870 34108 14922
rect 34108 14870 34110 14922
rect 34054 14868 34110 14870
rect 33068 13746 33124 13748
rect 33068 13694 33070 13746
rect 33070 13694 33122 13746
rect 33122 13694 33124 13746
rect 33068 13692 33124 13694
rect 33628 13692 33684 13748
rect 33180 13020 33236 13076
rect 32620 12236 32676 12292
rect 32732 12908 32788 12964
rect 31836 12178 31892 12180
rect 31836 12126 31838 12178
rect 31838 12126 31890 12178
rect 31890 12126 31892 12178
rect 31836 12124 31892 12126
rect 32732 12124 32788 12180
rect 32620 9826 32676 9828
rect 32620 9774 32622 9826
rect 32622 9774 32674 9826
rect 32674 9774 32676 9826
rect 32620 9772 32676 9774
rect 32844 9826 32900 9828
rect 32844 9774 32846 9826
rect 32846 9774 32898 9826
rect 32898 9774 32900 9826
rect 32844 9772 32900 9774
rect 31948 9548 32004 9604
rect 32340 9602 32396 9604
rect 32340 9550 32342 9602
rect 32342 9550 32394 9602
rect 32394 9550 32396 9602
rect 32340 9548 32396 9550
rect 32956 9548 33012 9604
rect 31612 8988 31668 9044
rect 32060 8988 32116 9044
rect 30940 8204 30996 8260
rect 30268 7532 30324 7588
rect 29932 6300 29988 6356
rect 30044 6860 30100 6916
rect 30156 6690 30212 6692
rect 30156 6638 30158 6690
rect 30158 6638 30210 6690
rect 30210 6638 30212 6690
rect 30156 6636 30212 6638
rect 30604 7532 30660 7588
rect 32172 8818 32228 8820
rect 32172 8766 32174 8818
rect 32174 8766 32226 8818
rect 32226 8766 32228 8818
rect 32172 8764 32228 8766
rect 32172 8258 32228 8260
rect 32172 8206 32174 8258
rect 32174 8206 32226 8258
rect 32226 8206 32228 8258
rect 32172 8204 32228 8206
rect 32508 7420 32564 7476
rect 30604 6860 30660 6916
rect 30212 6076 30268 6132
rect 30716 6524 30772 6580
rect 29708 5906 29764 5908
rect 29708 5854 29710 5906
rect 29710 5854 29762 5906
rect 29762 5854 29764 5906
rect 29708 5852 29764 5854
rect 29932 4284 29988 4340
rect 31388 5404 31444 5460
rect 31948 6524 32004 6580
rect 32172 6524 32228 6580
rect 32284 6300 32340 6356
rect 32620 5404 32676 5460
rect 33852 14364 33908 14420
rect 34300 14364 34356 14420
rect 35980 15820 36036 15876
rect 36484 16210 36540 16212
rect 36484 16158 36486 16210
rect 36486 16158 36538 16210
rect 36538 16158 36540 16210
rect 36484 16156 36540 16158
rect 36316 16044 36372 16100
rect 35532 15314 35588 15316
rect 35532 15262 35534 15314
rect 35534 15262 35586 15314
rect 35586 15262 35588 15314
rect 35532 15260 35588 15262
rect 35308 15148 35364 15204
rect 34524 14028 34580 14084
rect 34412 13916 34468 13972
rect 33846 13354 33902 13356
rect 33846 13302 33848 13354
rect 33848 13302 33900 13354
rect 33900 13302 33902 13354
rect 33846 13300 33902 13302
rect 33950 13354 34006 13356
rect 33950 13302 33952 13354
rect 33952 13302 34004 13354
rect 34004 13302 34006 13354
rect 33950 13300 34006 13302
rect 34054 13354 34110 13356
rect 34054 13302 34056 13354
rect 34056 13302 34108 13354
rect 34108 13302 34110 13354
rect 34054 13300 34110 13302
rect 34300 13356 34356 13412
rect 33852 12962 33908 12964
rect 33852 12910 33854 12962
rect 33854 12910 33906 12962
rect 33906 12910 33908 12962
rect 33852 12908 33908 12910
rect 34094 12850 34150 12852
rect 34094 12798 34096 12850
rect 34096 12798 34148 12850
rect 34148 12798 34150 12850
rect 34094 12796 34150 12798
rect 33908 12684 33964 12740
rect 35308 14028 35364 14084
rect 34636 13132 34692 13188
rect 34636 12962 34692 12964
rect 34636 12910 34638 12962
rect 34638 12910 34690 12962
rect 34690 12910 34692 12962
rect 35588 14140 35644 14196
rect 35756 13746 35812 13748
rect 35756 13694 35758 13746
rect 35758 13694 35810 13746
rect 35810 13694 35812 13746
rect 35756 13692 35812 13694
rect 35420 13356 35476 13412
rect 34636 12908 34692 12910
rect 35550 12962 35606 12964
rect 35550 12910 35552 12962
rect 35552 12910 35604 12962
rect 35604 12910 35606 12962
rect 35550 12908 35606 12910
rect 36204 15426 36260 15428
rect 36204 15374 36206 15426
rect 36206 15374 36258 15426
rect 36258 15374 36260 15426
rect 36204 15372 36260 15374
rect 36204 15036 36260 15092
rect 36298 14140 36354 14196
rect 34636 12684 34692 12740
rect 35868 12796 35924 12852
rect 36092 12796 36148 12852
rect 35252 12684 35308 12740
rect 33846 11786 33902 11788
rect 33846 11734 33848 11786
rect 33848 11734 33900 11786
rect 33900 11734 33902 11786
rect 33846 11732 33902 11734
rect 33950 11786 34006 11788
rect 33950 11734 33952 11786
rect 33952 11734 34004 11786
rect 34004 11734 34006 11786
rect 33950 11732 34006 11734
rect 34054 11786 34110 11788
rect 34054 11734 34056 11786
rect 34056 11734 34108 11786
rect 34108 11734 34110 11786
rect 34054 11732 34110 11734
rect 35644 12684 35700 12740
rect 33846 10218 33902 10220
rect 33846 10166 33848 10218
rect 33848 10166 33900 10218
rect 33900 10166 33902 10218
rect 33846 10164 33902 10166
rect 33950 10218 34006 10220
rect 33950 10166 33952 10218
rect 33952 10166 34004 10218
rect 34004 10166 34006 10218
rect 33950 10164 34006 10166
rect 34054 10218 34110 10220
rect 34054 10166 34056 10218
rect 34056 10166 34108 10218
rect 34108 10166 34110 10218
rect 34054 10164 34110 10166
rect 33628 9548 33684 9604
rect 33292 8764 33348 8820
rect 33846 8650 33902 8652
rect 33846 8598 33848 8650
rect 33848 8598 33900 8650
rect 33900 8598 33902 8650
rect 33846 8596 33902 8598
rect 33950 8650 34006 8652
rect 33950 8598 33952 8650
rect 33952 8598 34004 8650
rect 34004 8598 34006 8650
rect 33950 8596 34006 8598
rect 34054 8650 34110 8652
rect 34054 8598 34056 8650
rect 34056 8598 34108 8650
rect 34108 8598 34110 8650
rect 34054 8596 34110 8598
rect 34412 8316 34468 8372
rect 33846 7082 33902 7084
rect 33846 7030 33848 7082
rect 33848 7030 33900 7082
rect 33900 7030 33902 7082
rect 33846 7028 33902 7030
rect 33950 7082 34006 7084
rect 33950 7030 33952 7082
rect 33952 7030 34004 7082
rect 34004 7030 34006 7082
rect 33950 7028 34006 7030
rect 34054 7082 34110 7084
rect 34054 7030 34056 7082
rect 34056 7030 34108 7082
rect 34108 7030 34110 7082
rect 34054 7028 34110 7030
rect 34972 9548 35028 9604
rect 35252 9548 35308 9604
rect 35980 9212 36036 9268
rect 35756 8258 35812 8260
rect 34692 8146 34748 8148
rect 34692 8094 34694 8146
rect 34694 8094 34746 8146
rect 34746 8094 34748 8146
rect 34692 8092 34748 8094
rect 34300 7474 34356 7476
rect 34300 7422 34302 7474
rect 34302 7422 34354 7474
rect 34354 7422 34356 7474
rect 34300 7420 34356 7422
rect 33964 6690 34020 6692
rect 33964 6638 33966 6690
rect 33966 6638 34018 6690
rect 34018 6638 34020 6690
rect 33964 6636 34020 6638
rect 34468 7308 34524 7364
rect 34206 6578 34262 6580
rect 34206 6526 34208 6578
rect 34208 6526 34260 6578
rect 34260 6526 34262 6578
rect 34206 6524 34262 6526
rect 33404 5404 33460 5460
rect 34076 6412 34132 6468
rect 34188 5852 34244 5908
rect 35756 8206 35758 8258
rect 35758 8206 35810 8258
rect 35810 8206 35812 8258
rect 35756 8204 35812 8206
rect 35252 7980 35308 8036
rect 35532 8092 35588 8148
rect 35214 7644 35270 7700
rect 35084 7420 35140 7476
rect 36372 13468 36428 13524
rect 36540 12684 36596 12740
rect 36988 16716 37044 16772
rect 36876 16156 36932 16212
rect 36876 15372 36932 15428
rect 37212 16770 37268 16772
rect 37212 16718 37214 16770
rect 37214 16718 37266 16770
rect 37266 16718 37268 16770
rect 37212 16716 37268 16718
rect 37660 21084 37716 21140
rect 38332 27020 38388 27076
rect 38508 26682 38564 26684
rect 38508 26630 38510 26682
rect 38510 26630 38562 26682
rect 38562 26630 38564 26682
rect 38508 26628 38564 26630
rect 38612 26682 38668 26684
rect 38612 26630 38614 26682
rect 38614 26630 38666 26682
rect 38666 26630 38668 26682
rect 38612 26628 38668 26630
rect 38716 26682 38772 26684
rect 38716 26630 38718 26682
rect 38718 26630 38770 26682
rect 38770 26630 38772 26682
rect 38716 26628 38772 26630
rect 38332 25788 38388 25844
rect 38508 25114 38564 25116
rect 38508 25062 38510 25114
rect 38510 25062 38562 25114
rect 38562 25062 38564 25114
rect 38508 25060 38564 25062
rect 38612 25114 38668 25116
rect 38612 25062 38614 25114
rect 38614 25062 38666 25114
rect 38666 25062 38668 25114
rect 38612 25060 38668 25062
rect 38716 25114 38772 25116
rect 38716 25062 38718 25114
rect 38718 25062 38770 25114
rect 38770 25062 38772 25114
rect 38716 25060 38772 25062
rect 38220 24780 38276 24836
rect 38276 24610 38332 24612
rect 38276 24558 38278 24610
rect 38278 24558 38330 24610
rect 38330 24558 38332 24610
rect 38276 24556 38332 24558
rect 38276 24108 38332 24164
rect 38508 23546 38564 23548
rect 38508 23494 38510 23546
rect 38510 23494 38562 23546
rect 38562 23494 38564 23546
rect 38508 23492 38564 23494
rect 38612 23546 38668 23548
rect 38612 23494 38614 23546
rect 38614 23494 38666 23546
rect 38666 23494 38668 23546
rect 38612 23492 38668 23494
rect 38716 23546 38772 23548
rect 38716 23494 38718 23546
rect 38718 23494 38770 23546
rect 38770 23494 38772 23546
rect 38716 23492 38772 23494
rect 38332 22876 38388 22932
rect 38508 21978 38564 21980
rect 38508 21926 38510 21978
rect 38510 21926 38562 21978
rect 38562 21926 38564 21978
rect 38508 21924 38564 21926
rect 38612 21978 38668 21980
rect 38612 21926 38614 21978
rect 38614 21926 38666 21978
rect 38666 21926 38668 21978
rect 38612 21924 38668 21926
rect 38716 21978 38772 21980
rect 38716 21926 38718 21978
rect 38718 21926 38770 21978
rect 38770 21926 38772 21978
rect 38716 21924 38772 21926
rect 39004 24556 39060 24612
rect 38892 20860 38948 20916
rect 37996 20748 38052 20804
rect 38508 20410 38564 20412
rect 38508 20358 38510 20410
rect 38510 20358 38562 20410
rect 38562 20358 38564 20410
rect 38508 20356 38564 20358
rect 38612 20410 38668 20412
rect 38612 20358 38614 20410
rect 38614 20358 38666 20410
rect 38666 20358 38668 20410
rect 38612 20356 38668 20358
rect 38716 20410 38772 20412
rect 38716 20358 38718 20410
rect 38718 20358 38770 20410
rect 38770 20358 38772 20410
rect 38716 20356 38772 20358
rect 38332 19404 38388 19460
rect 38444 19964 38500 20020
rect 37604 19234 37660 19236
rect 37604 19182 37606 19234
rect 37606 19182 37658 19234
rect 37658 19182 37660 19234
rect 37604 19180 37660 19182
rect 38332 19234 38388 19236
rect 38332 19182 38334 19234
rect 38334 19182 38386 19234
rect 38386 19182 38388 19234
rect 38332 19180 38388 19182
rect 38508 18842 38564 18844
rect 38508 18790 38510 18842
rect 38510 18790 38562 18842
rect 38562 18790 38564 18842
rect 38508 18788 38564 18790
rect 38612 18842 38668 18844
rect 38612 18790 38614 18842
rect 38614 18790 38666 18842
rect 38666 18790 38668 18842
rect 38612 18788 38668 18790
rect 38716 18842 38772 18844
rect 38716 18790 38718 18842
rect 38718 18790 38770 18842
rect 38770 18790 38772 18842
rect 38716 18788 38772 18790
rect 37996 17164 38052 17220
rect 37604 17052 37660 17108
rect 38508 17274 38564 17276
rect 38508 17222 38510 17274
rect 38510 17222 38562 17274
rect 38562 17222 38564 17274
rect 38508 17220 38564 17222
rect 38612 17274 38668 17276
rect 38612 17222 38614 17274
rect 38614 17222 38666 17274
rect 38666 17222 38668 17274
rect 38612 17220 38668 17222
rect 38716 17274 38772 17276
rect 38716 17222 38718 17274
rect 38718 17222 38770 17274
rect 38770 17222 38772 17274
rect 38716 17220 38772 17222
rect 38332 17052 38388 17108
rect 37324 16604 37380 16660
rect 37100 16098 37156 16100
rect 37100 16046 37102 16098
rect 37102 16046 37154 16098
rect 37154 16046 37156 16098
rect 37100 16044 37156 16046
rect 36988 15260 37044 15316
rect 37380 16322 37436 16324
rect 37380 16270 37382 16322
rect 37382 16270 37434 16322
rect 37434 16270 37436 16322
rect 37380 16268 37436 16270
rect 38508 15706 38564 15708
rect 38508 15654 38510 15706
rect 38510 15654 38562 15706
rect 38562 15654 38564 15706
rect 38508 15652 38564 15654
rect 38612 15706 38668 15708
rect 38612 15654 38614 15706
rect 38614 15654 38666 15706
rect 38666 15654 38668 15706
rect 38612 15652 38668 15654
rect 38716 15706 38772 15708
rect 38716 15654 38718 15706
rect 38718 15654 38770 15706
rect 38770 15654 38772 15706
rect 38716 15652 38772 15654
rect 37996 14418 38052 14420
rect 37996 14366 37998 14418
rect 37998 14366 38050 14418
rect 38050 14366 38052 14418
rect 37996 14364 38052 14366
rect 37604 14306 37660 14308
rect 37604 14254 37606 14306
rect 37606 14254 37658 14306
rect 37658 14254 37660 14306
rect 37604 14252 37660 14254
rect 36876 13244 36932 13300
rect 36988 13356 37044 13412
rect 37212 13356 37268 13412
rect 37436 13468 37492 13524
rect 37156 12962 37212 12964
rect 37156 12910 37158 12962
rect 37158 12910 37210 12962
rect 37210 12910 37212 12962
rect 37156 12908 37212 12910
rect 37268 10834 37324 10836
rect 37268 10782 37270 10834
rect 37270 10782 37322 10834
rect 37322 10782 37324 10834
rect 37268 10780 37324 10782
rect 36652 10722 36708 10724
rect 36652 10670 36654 10722
rect 36654 10670 36706 10722
rect 36706 10670 36708 10722
rect 36652 10668 36708 10670
rect 37156 9212 37212 9268
rect 37324 8764 37380 8820
rect 36988 8652 37044 8708
rect 36204 7980 36260 8036
rect 36652 8428 36708 8484
rect 34860 5964 34916 6020
rect 34636 5906 34692 5908
rect 34636 5854 34638 5906
rect 34638 5854 34690 5906
rect 34690 5854 34692 5906
rect 34636 5852 34692 5854
rect 35196 6524 35252 6580
rect 35644 6636 35700 6692
rect 33846 5514 33902 5516
rect 33846 5462 33848 5514
rect 33848 5462 33900 5514
rect 33900 5462 33902 5514
rect 33846 5460 33902 5462
rect 33950 5514 34006 5516
rect 33950 5462 33952 5514
rect 33952 5462 34004 5514
rect 34004 5462 34006 5514
rect 33950 5460 34006 5462
rect 34054 5514 34110 5516
rect 34054 5462 34056 5514
rect 34056 5462 34108 5514
rect 34108 5462 34110 5514
rect 34054 5460 34110 5462
rect 35420 5180 35476 5236
rect 37156 7644 37212 7700
rect 37324 7980 37380 8036
rect 33846 3946 33902 3948
rect 33846 3894 33848 3946
rect 33848 3894 33900 3946
rect 33900 3894 33902 3946
rect 33846 3892 33902 3894
rect 33950 3946 34006 3948
rect 33950 3894 33952 3946
rect 33952 3894 34004 3946
rect 34004 3894 34006 3946
rect 33950 3892 34006 3894
rect 34054 3946 34110 3948
rect 34054 3894 34056 3946
rect 34056 3894 34108 3946
rect 34108 3894 34110 3946
rect 34054 3892 34110 3894
rect 35980 6076 36036 6132
rect 37156 6076 37212 6132
rect 36260 5234 36316 5236
rect 36260 5182 36262 5234
rect 36262 5182 36314 5234
rect 36314 5182 36316 5234
rect 36260 5180 36316 5182
rect 37156 5234 37212 5236
rect 37156 5182 37158 5234
rect 37158 5182 37210 5234
rect 37210 5182 37212 5234
rect 37156 5180 37212 5182
rect 35252 3724 35308 3780
rect 36204 3778 36260 3780
rect 36204 3726 36206 3778
rect 36206 3726 36258 3778
rect 36258 3726 36260 3778
rect 36204 3724 36260 3726
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
rect 26236 3500 26292 3556
rect 24220 2492 24276 2548
rect 27804 3554 27860 3556
rect 27804 3502 27806 3554
rect 27806 3502 27858 3554
rect 27858 3502 27860 3554
rect 27804 3500 27860 3502
rect 28028 3500 28084 3556
rect 28812 3554 28868 3556
rect 28812 3502 28814 3554
rect 28814 3502 28866 3554
rect 28866 3502 28868 3554
rect 28812 3500 28868 3502
rect 29652 3554 29708 3556
rect 29652 3502 29654 3554
rect 29654 3502 29706 3554
rect 29706 3502 29708 3554
rect 29652 3500 29708 3502
rect 29820 3500 29876 3556
rect 29204 3442 29260 3444
rect 29204 3390 29206 3442
rect 29206 3390 29258 3442
rect 29258 3390 29260 3442
rect 29204 3388 29260 3390
rect 29184 3162 29240 3164
rect 29184 3110 29186 3162
rect 29186 3110 29238 3162
rect 29238 3110 29240 3162
rect 29184 3108 29240 3110
rect 29288 3162 29344 3164
rect 29288 3110 29290 3162
rect 29290 3110 29342 3162
rect 29342 3110 29344 3162
rect 29288 3108 29344 3110
rect 29392 3162 29448 3164
rect 29392 3110 29394 3162
rect 29394 3110 29446 3162
rect 29446 3110 29448 3162
rect 29392 3108 29448 3110
rect 30492 3554 30548 3556
rect 30492 3502 30494 3554
rect 30494 3502 30546 3554
rect 30546 3502 30548 3554
rect 30492 3500 30548 3502
rect 30884 3554 30940 3556
rect 30884 3502 30886 3554
rect 30886 3502 30938 3554
rect 30938 3502 30940 3554
rect 30884 3500 30940 3502
rect 38108 13020 38164 13076
rect 37902 12850 37958 12852
rect 37902 12798 37904 12850
rect 37904 12798 37956 12850
rect 37956 12798 37958 12850
rect 37902 12796 37958 12798
rect 37660 12684 37716 12740
rect 38332 14252 38388 14308
rect 38508 14138 38564 14140
rect 38508 14086 38510 14138
rect 38510 14086 38562 14138
rect 38562 14086 38564 14138
rect 38508 14084 38564 14086
rect 38612 14138 38668 14140
rect 38612 14086 38614 14138
rect 38614 14086 38666 14138
rect 38666 14086 38668 14138
rect 38612 14084 38668 14086
rect 38716 14138 38772 14140
rect 38716 14086 38718 14138
rect 38718 14086 38770 14138
rect 38770 14086 38772 14138
rect 38716 14084 38772 14086
rect 38508 12570 38564 12572
rect 38508 12518 38510 12570
rect 38510 12518 38562 12570
rect 38562 12518 38564 12570
rect 38508 12516 38564 12518
rect 38612 12570 38668 12572
rect 38612 12518 38614 12570
rect 38614 12518 38666 12570
rect 38666 12518 38668 12570
rect 38612 12516 38668 12518
rect 38716 12570 38772 12572
rect 38716 12518 38718 12570
rect 38718 12518 38770 12570
rect 38770 12518 38772 12570
rect 38716 12516 38772 12518
rect 37604 11282 37660 11284
rect 37604 11230 37606 11282
rect 37606 11230 37658 11282
rect 37658 11230 37660 11282
rect 37604 11228 37660 11230
rect 38332 11228 38388 11284
rect 38508 11002 38564 11004
rect 38508 10950 38510 11002
rect 38510 10950 38562 11002
rect 38562 10950 38564 11002
rect 38508 10948 38564 10950
rect 38612 11002 38668 11004
rect 38612 10950 38614 11002
rect 38614 10950 38666 11002
rect 38666 10950 38668 11002
rect 38612 10948 38668 10950
rect 38716 11002 38772 11004
rect 38716 10950 38718 11002
rect 38718 10950 38770 11002
rect 38770 10950 38772 11002
rect 38716 10948 38772 10950
rect 38220 10780 38276 10836
rect 37660 10668 37716 10724
rect 37902 9826 37958 9828
rect 37902 9774 37904 9826
rect 37904 9774 37956 9826
rect 37956 9774 37958 9826
rect 37902 9772 37958 9774
rect 38108 9100 38164 9156
rect 37548 8428 37604 8484
rect 37902 8370 37958 8372
rect 37902 8318 37904 8370
rect 37904 8318 37956 8370
rect 37956 8318 37958 8370
rect 37902 8316 37958 8318
rect 37660 8258 37716 8260
rect 37660 8206 37662 8258
rect 37662 8206 37714 8258
rect 37714 8206 37716 8258
rect 37660 8204 37716 8206
rect 38508 9434 38564 9436
rect 38508 9382 38510 9434
rect 38510 9382 38562 9434
rect 38562 9382 38564 9434
rect 38508 9380 38564 9382
rect 38612 9434 38668 9436
rect 38612 9382 38614 9434
rect 38614 9382 38666 9434
rect 38666 9382 38668 9434
rect 38612 9380 38668 9382
rect 38716 9434 38772 9436
rect 38716 9382 38718 9434
rect 38718 9382 38770 9434
rect 38770 9382 38772 9434
rect 38716 9380 38772 9382
rect 37436 7308 37492 7364
rect 37772 7420 37828 7476
rect 37660 6524 37716 6580
rect 37902 5964 37958 6020
rect 38108 6524 38164 6580
rect 37996 5346 38052 5348
rect 37996 5294 37998 5346
rect 37998 5294 38050 5346
rect 38050 5294 38052 5346
rect 37996 5292 38052 5294
rect 38332 8316 38388 8372
rect 38508 7866 38564 7868
rect 38508 7814 38510 7866
rect 38510 7814 38562 7866
rect 38562 7814 38564 7866
rect 38508 7812 38564 7814
rect 38612 7866 38668 7868
rect 38612 7814 38614 7866
rect 38614 7814 38666 7866
rect 38666 7814 38668 7866
rect 38612 7812 38668 7814
rect 38716 7866 38772 7868
rect 38716 7814 38718 7866
rect 38718 7814 38770 7866
rect 38770 7814 38772 7866
rect 38716 7812 38772 7814
rect 38332 7474 38388 7476
rect 38332 7422 38334 7474
rect 38334 7422 38386 7474
rect 38386 7422 38388 7474
rect 38332 7420 38388 7422
rect 38508 6298 38564 6300
rect 38508 6246 38510 6298
rect 38510 6246 38562 6298
rect 38562 6246 38564 6298
rect 38508 6244 38564 6246
rect 38612 6298 38668 6300
rect 38612 6246 38614 6298
rect 38614 6246 38666 6298
rect 38666 6246 38668 6298
rect 38612 6244 38668 6246
rect 38716 6298 38772 6300
rect 38716 6246 38718 6298
rect 38718 6246 38770 6298
rect 38770 6246 38772 6298
rect 38716 6244 38772 6246
rect 38220 5180 38276 5236
rect 38332 5404 38388 5460
rect 38508 4730 38564 4732
rect 38508 4678 38510 4730
rect 38510 4678 38562 4730
rect 38562 4678 38564 4730
rect 38508 4676 38564 4678
rect 38612 4730 38668 4732
rect 38612 4678 38614 4730
rect 38614 4678 38666 4730
rect 38666 4678 38668 4730
rect 38612 4676 38668 4678
rect 38716 4730 38772 4732
rect 38716 4678 38718 4730
rect 38718 4678 38770 4730
rect 38770 4678 38772 4730
rect 38716 4676 38772 4678
rect 38508 3162 38564 3164
rect 38508 3110 38510 3162
rect 38510 3110 38562 3162
rect 38562 3110 38564 3162
rect 38508 3108 38564 3110
rect 38612 3162 38668 3164
rect 38612 3110 38614 3162
rect 38614 3110 38666 3162
rect 38666 3110 38668 3162
rect 38612 3108 38668 3110
rect 38716 3162 38772 3164
rect 38716 3110 38718 3162
rect 38718 3110 38770 3162
rect 38770 3110 38772 3162
rect 38716 3108 38772 3110
<< metal3 >>
rect 39200 37492 40000 37520
rect 38322 37436 38332 37492
rect 38388 37436 40000 37492
rect 39200 37408 40000 37436
rect 37594 36988 37604 37044
rect 37660 36988 38332 37044
rect 38388 36988 38398 37044
rect 5864 36820 5874 36876
rect 5930 36820 5978 36876
rect 6034 36820 6082 36876
rect 6138 36820 6148 36876
rect 15188 36820 15198 36876
rect 15254 36820 15302 36876
rect 15358 36820 15406 36876
rect 15462 36820 15472 36876
rect 24512 36820 24522 36876
rect 24578 36820 24626 36876
rect 24682 36820 24730 36876
rect 24786 36820 24796 36876
rect 33836 36820 33846 36876
rect 33902 36820 33950 36876
rect 34006 36820 34054 36876
rect 34110 36820 34120 36876
rect 19170 36652 19180 36708
rect 19236 36652 19964 36708
rect 20020 36652 20030 36708
rect 24322 36540 24332 36596
rect 24388 36540 28588 36596
rect 28644 36540 28654 36596
rect 12338 36428 12348 36484
rect 12404 36428 13244 36484
rect 13300 36428 13310 36484
rect 30706 36316 30716 36372
rect 30772 36316 36148 36372
rect 36204 36316 36214 36372
rect 8866 36204 8876 36260
rect 8932 36204 13916 36260
rect 13972 36204 13982 36260
rect 31378 36204 31388 36260
rect 31444 36204 33068 36260
rect 33124 36204 33134 36260
rect 35074 36204 35084 36260
rect 35140 36204 35980 36260
rect 36036 36204 36046 36260
rect 10526 36036 10536 36092
rect 10592 36036 10640 36092
rect 10696 36036 10744 36092
rect 10800 36036 10810 36092
rect 19850 36036 19860 36092
rect 19916 36036 19964 36092
rect 20020 36036 20068 36092
rect 20124 36036 20134 36092
rect 29174 36036 29184 36092
rect 29240 36036 29288 36092
rect 29344 36036 29392 36092
rect 29448 36036 29458 36092
rect 38498 36036 38508 36092
rect 38564 36036 38612 36092
rect 38668 36036 38716 36092
rect 38772 36036 38782 36092
rect 20290 35868 20300 35924
rect 20356 35868 20972 35924
rect 21028 35868 24556 35924
rect 24612 35868 24622 35924
rect 22754 35756 22764 35812
rect 22820 35756 24332 35812
rect 24388 35756 24398 35812
rect 5506 35644 5516 35700
rect 5572 35644 5796 35700
rect 5852 35644 6188 35700
rect 6244 35644 9548 35700
rect 9604 35644 9614 35700
rect 13346 35644 13356 35700
rect 13412 35644 16268 35700
rect 16324 35644 16334 35700
rect 20850 35644 20860 35700
rect 20916 35644 25228 35700
rect 25284 35644 25294 35700
rect 30930 35644 30940 35700
rect 30996 35644 31276 35700
rect 31332 35644 31342 35700
rect 6962 35532 6972 35588
rect 7028 35532 8764 35588
rect 8820 35532 8830 35588
rect 15586 35532 15596 35588
rect 15652 35532 18060 35588
rect 18116 35532 18126 35588
rect 20570 35532 20580 35588
rect 20636 35532 21756 35588
rect 21812 35532 28028 35588
rect 28084 35532 28094 35588
rect 5170 35420 5180 35476
rect 5236 35420 7588 35476
rect 12226 35420 12236 35476
rect 12292 35420 12796 35476
rect 12852 35420 15820 35476
rect 15876 35420 15886 35476
rect 24434 35420 24444 35476
rect 24500 35420 25788 35476
rect 25844 35420 25854 35476
rect 28130 35420 28140 35476
rect 28196 35420 37996 35476
rect 38052 35420 38062 35476
rect 7532 35364 7588 35420
rect 7522 35308 7532 35364
rect 7588 35308 7598 35364
rect 26674 35308 26684 35364
rect 26740 35308 26908 35364
rect 26964 35308 26974 35364
rect 5864 35252 5874 35308
rect 5930 35252 5978 35308
rect 6034 35252 6082 35308
rect 6138 35252 6148 35308
rect 15188 35252 15198 35308
rect 15254 35252 15302 35308
rect 15358 35252 15406 35308
rect 15462 35252 15472 35308
rect 24512 35252 24522 35308
rect 24578 35252 24626 35308
rect 24682 35252 24730 35308
rect 24786 35252 24796 35308
rect 33836 35252 33846 35308
rect 33902 35252 33950 35308
rect 34006 35252 34054 35308
rect 34110 35252 34120 35308
rect 10098 35196 10108 35252
rect 10164 35196 10948 35252
rect 11004 35196 12348 35252
rect 12404 35196 12414 35252
rect 14242 35196 14252 35252
rect 14308 35196 15036 35252
rect 15092 35196 15102 35252
rect 21074 35196 21084 35252
rect 21140 35196 22316 35252
rect 22372 35196 22382 35252
rect 25666 35196 25676 35252
rect 25732 35196 27244 35252
rect 27300 35196 27310 35252
rect 27794 35196 27804 35252
rect 27860 35196 29708 35252
rect 29764 35196 29774 35252
rect 14354 35084 14364 35140
rect 14420 35084 15708 35140
rect 15764 35084 15774 35140
rect 20794 35084 20804 35140
rect 20860 35084 21868 35140
rect 21924 35084 24052 35140
rect 24108 35084 24892 35140
rect 24948 35084 24958 35140
rect 25554 35084 25564 35140
rect 25620 35084 29036 35140
rect 29092 35084 29102 35140
rect 31154 35084 31164 35140
rect 31220 35084 34412 35140
rect 34468 35084 34478 35140
rect 22642 34972 22652 35028
rect 22708 34972 25900 35028
rect 25956 34972 25966 35028
rect 26898 34972 26908 35028
rect 26964 34972 33180 35028
rect 33236 34972 33246 35028
rect 35522 34972 35532 35028
rect 35588 34972 35644 35028
rect 35700 34972 35710 35028
rect 12338 34860 12348 34916
rect 12404 34860 13748 34916
rect 13804 34860 15932 34916
rect 15988 34860 15998 34916
rect 19618 34860 19628 34916
rect 19684 34860 20076 34916
rect 20132 34860 22876 34916
rect 22932 34860 22942 34916
rect 23314 34860 23324 34916
rect 23380 34860 26012 34916
rect 26068 34860 26078 34916
rect 28522 34860 28532 34916
rect 28588 34860 29036 34916
rect 29092 34860 29102 34916
rect 30482 34860 30492 34916
rect 30548 34860 31836 34916
rect 31892 34860 31902 34916
rect 33730 34860 33740 34916
rect 33796 34860 35420 34916
rect 35476 34860 35486 34916
rect 8194 34748 8204 34804
rect 8260 34748 10220 34804
rect 10276 34748 10286 34804
rect 16594 34748 16604 34804
rect 16660 34748 18620 34804
rect 18676 34748 19068 34804
rect 19124 34748 19134 34804
rect 35270 34748 35308 34804
rect 35364 34748 36372 34804
rect 36428 34748 36438 34804
rect 15922 34636 15932 34692
rect 15988 34636 16940 34692
rect 16996 34636 17276 34692
rect 17332 34636 18788 34692
rect 18844 34636 18854 34692
rect 39200 34580 40000 34608
rect 38892 34524 40000 34580
rect 10526 34468 10536 34524
rect 10592 34468 10640 34524
rect 10696 34468 10744 34524
rect 10800 34468 10810 34524
rect 19850 34468 19860 34524
rect 19916 34468 19964 34524
rect 20020 34468 20068 34524
rect 20124 34468 20134 34524
rect 29174 34468 29184 34524
rect 29240 34468 29288 34524
rect 29344 34468 29392 34524
rect 29448 34468 29458 34524
rect 38498 34468 38508 34524
rect 38564 34468 38612 34524
rect 38668 34468 38716 34524
rect 38772 34468 38782 34524
rect 30034 34412 30044 34468
rect 30100 34412 33964 34468
rect 34020 34412 34030 34468
rect 35410 34412 35420 34468
rect 35476 34412 35644 34468
rect 35700 34412 35710 34468
rect 15922 34300 15932 34356
rect 15988 34300 16604 34356
rect 16660 34300 16670 34356
rect 19170 34300 19180 34356
rect 19236 34300 20412 34356
rect 20468 34300 20478 34356
rect 29820 34300 36204 34356
rect 36260 34300 36270 34356
rect 29820 34244 29876 34300
rect 38892 34244 38948 34524
rect 39200 34496 40000 34524
rect 28914 34188 28924 34244
rect 28980 34188 29876 34244
rect 35074 34188 35084 34244
rect 35140 34188 38948 34244
rect 8586 34076 8596 34132
rect 8652 34076 9436 34132
rect 9492 34076 9502 34132
rect 15026 33852 15036 33908
rect 15092 33852 17948 33908
rect 18004 33852 18014 33908
rect 29820 33796 29876 34188
rect 31154 34076 31164 34132
rect 31220 34076 31724 34132
rect 31780 34076 31790 34132
rect 32162 34076 32172 34132
rect 32228 34076 36260 34132
rect 36316 34076 36326 34132
rect 30818 33964 30828 34020
rect 30884 33964 32060 34020
rect 32116 33964 32126 34020
rect 32722 33964 32732 34020
rect 32788 33964 37324 34020
rect 37380 33964 37390 34020
rect 31322 33852 31332 33908
rect 31388 33852 33628 33908
rect 33684 33852 33694 33908
rect 33954 33852 33964 33908
rect 34020 33852 34244 33908
rect 35410 33852 35420 33908
rect 35476 33852 35644 33908
rect 35700 33852 35710 33908
rect 37986 33852 37996 33908
rect 38052 33852 39004 33908
rect 39060 33852 39070 33908
rect 34188 33796 34244 33852
rect 8978 33740 8988 33796
rect 9044 33740 9436 33796
rect 9492 33740 9502 33796
rect 14354 33740 14364 33796
rect 14420 33740 14430 33796
rect 18386 33740 18396 33796
rect 18452 33740 23996 33796
rect 24052 33740 24062 33796
rect 25106 33740 25116 33796
rect 25172 33740 27244 33796
rect 27300 33740 27310 33796
rect 29810 33740 29820 33796
rect 29876 33740 29886 33796
rect 34178 33740 34188 33796
rect 34244 33740 34254 33796
rect 5864 33684 5874 33740
rect 5930 33684 5978 33740
rect 6034 33684 6082 33740
rect 6138 33684 6148 33740
rect 14364 33572 14420 33740
rect 15188 33684 15198 33740
rect 15254 33684 15302 33740
rect 15358 33684 15406 33740
rect 15462 33684 15472 33740
rect 24512 33684 24522 33740
rect 24578 33684 24626 33740
rect 24682 33684 24730 33740
rect 24786 33684 24796 33740
rect 33836 33684 33846 33740
rect 33902 33684 33950 33740
rect 34006 33684 34054 33740
rect 34110 33684 34120 33740
rect 18274 33628 18284 33684
rect 18340 33628 19012 33684
rect 28242 33628 28252 33684
rect 28308 33628 28318 33684
rect 32946 33628 32956 33684
rect 33012 33628 33022 33684
rect 18956 33572 19012 33628
rect 28252 33572 28308 33628
rect 32956 33572 33012 33628
rect 11218 33516 11228 33572
rect 11284 33516 12012 33572
rect 12068 33516 12078 33572
rect 12450 33516 12460 33572
rect 12516 33516 14420 33572
rect 16818 33516 16828 33572
rect 16884 33516 17836 33572
rect 17892 33516 17902 33572
rect 18946 33516 18956 33572
rect 19012 33516 19022 33572
rect 28252 33516 31052 33572
rect 31108 33516 31612 33572
rect 31668 33516 33012 33572
rect 9426 33404 9436 33460
rect 9492 33404 10444 33460
rect 10500 33404 13972 33460
rect 25106 33404 25116 33460
rect 25172 33404 27692 33460
rect 27748 33404 27758 33460
rect 28354 33404 28364 33460
rect 28420 33404 30586 33460
rect 30642 33404 30652 33460
rect 30818 33404 30828 33460
rect 30884 33404 32172 33460
rect 32228 33404 32238 33460
rect 35074 33404 35084 33460
rect 35140 33404 35150 33460
rect 35858 33404 35868 33460
rect 35924 33404 35934 33460
rect 13916 33348 13972 33404
rect 35084 33348 35140 33404
rect 10042 33292 10052 33348
rect 10108 33292 10780 33348
rect 10836 33292 11340 33348
rect 11396 33292 11406 33348
rect 13906 33292 13916 33348
rect 13972 33292 14252 33348
rect 14308 33292 14318 33348
rect 22138 33292 22148 33348
rect 22204 33292 25282 33348
rect 25338 33292 26180 33348
rect 27794 33292 27804 33348
rect 27860 33292 35140 33348
rect 26124 33236 26180 33292
rect 35868 33236 35924 33404
rect 37650 33292 37660 33348
rect 37716 33292 38220 33348
rect 38276 33292 38286 33348
rect 7522 33180 7532 33236
rect 7588 33180 12460 33236
rect 12516 33180 12526 33236
rect 17490 33180 17500 33236
rect 17556 33180 19404 33236
rect 19460 33180 20076 33236
rect 20132 33180 20142 33236
rect 20402 33180 20412 33236
rect 20468 33180 21308 33236
rect 21364 33180 21374 33236
rect 23986 33180 23996 33236
rect 24052 33180 24276 33236
rect 24332 33180 24342 33236
rect 26124 33180 28028 33236
rect 28084 33180 28094 33236
rect 34402 33180 34412 33236
rect 34468 33180 35028 33236
rect 35084 33180 35924 33236
rect 36978 33180 36988 33236
rect 37044 33180 38108 33236
rect 38164 33180 38174 33236
rect 8754 33068 8764 33124
rect 8820 33068 11116 33124
rect 11172 33068 11182 33124
rect 18162 33068 18172 33124
rect 18228 33068 23156 33124
rect 23212 33068 25228 33124
rect 25284 33068 26292 33124
rect 26348 33068 26358 33124
rect 26852 33068 29316 33124
rect 29372 33068 29382 33124
rect 33394 33068 33404 33124
rect 33460 33068 36372 33124
rect 36428 33068 36652 33124
rect 36708 33068 36718 33124
rect 26852 33012 26908 33068
rect 35868 33012 35924 33068
rect 12226 32956 12236 33012
rect 12292 32956 12908 33012
rect 12964 32956 12974 33012
rect 23986 32956 23996 33012
rect 24052 32956 26908 33012
rect 30146 32956 30156 33012
rect 30212 32956 35644 33012
rect 35700 32956 35710 33012
rect 35858 32956 35868 33012
rect 35924 32956 35934 33012
rect 10526 32900 10536 32956
rect 10592 32900 10640 32956
rect 10696 32900 10744 32956
rect 10800 32900 10810 32956
rect 19850 32900 19860 32956
rect 19916 32900 19964 32956
rect 20020 32900 20068 32956
rect 20124 32900 20134 32956
rect 29174 32900 29184 32956
rect 29240 32900 29288 32956
rect 29344 32900 29392 32956
rect 29448 32900 29458 32956
rect 38498 32900 38508 32956
rect 38564 32900 38612 32956
rect 38668 32900 38716 32956
rect 38772 32900 38782 32956
rect 10882 32844 10892 32900
rect 10948 32844 16044 32900
rect 16100 32844 16110 32900
rect 30930 32844 30940 32900
rect 30996 32844 31724 32900
rect 31780 32844 31790 32900
rect 35410 32844 35420 32900
rect 35476 32844 36540 32900
rect 36596 32844 36606 32900
rect 7746 32732 7756 32788
rect 7812 32732 8428 32788
rect 8484 32732 9940 32788
rect 21718 32732 21756 32788
rect 21812 32732 21822 32788
rect 27682 32732 27692 32788
rect 27748 32732 29260 32788
rect 29316 32732 29326 32788
rect 30034 32732 30044 32788
rect 30100 32732 31164 32788
rect 31220 32732 31230 32788
rect 36652 32732 36876 32788
rect 36932 32732 36942 32788
rect 9884 32676 9940 32732
rect 9874 32620 9884 32676
rect 9940 32620 10892 32676
rect 10948 32620 10958 32676
rect 11666 32620 11676 32676
rect 11732 32620 12348 32676
rect 12404 32620 16716 32676
rect 16772 32620 18060 32676
rect 18116 32620 18126 32676
rect 19618 32620 19628 32676
rect 19684 32620 23324 32676
rect 23380 32620 23390 32676
rect 24770 32620 24780 32676
rect 24836 32620 25116 32676
rect 25172 32620 25182 32676
rect 26282 32620 26292 32676
rect 26348 32620 26842 32676
rect 26898 32620 26908 32676
rect 31434 32620 31444 32676
rect 31500 32620 31836 32676
rect 31892 32620 31902 32676
rect 34076 32620 34412 32676
rect 34468 32620 34478 32676
rect 34076 32564 34132 32620
rect 7354 32508 7364 32564
rect 7420 32508 8428 32564
rect 8484 32508 8494 32564
rect 9986 32508 9996 32564
rect 10052 32508 11116 32564
rect 11172 32508 11182 32564
rect 13346 32508 13356 32564
rect 13412 32508 14364 32564
rect 14420 32508 14430 32564
rect 20010 32508 20020 32564
rect 20076 32508 20524 32564
rect 20580 32508 20590 32564
rect 24602 32508 24612 32564
rect 24668 32508 26684 32564
rect 26740 32508 26750 32564
rect 31388 32508 34132 32564
rect 34290 32508 34300 32564
rect 34356 32508 35308 32564
rect 35364 32508 35374 32564
rect 9996 32452 10052 32508
rect 7186 32396 7196 32452
rect 7252 32396 7644 32452
rect 7700 32396 10052 32452
rect 11218 32396 11228 32452
rect 11284 32396 11900 32452
rect 11956 32396 11966 32452
rect 14028 32340 14084 32508
rect 31388 32452 31444 32508
rect 16034 32396 16044 32452
rect 16100 32396 17612 32452
rect 17668 32396 17678 32452
rect 23650 32396 23660 32452
rect 23716 32396 24108 32452
rect 24164 32396 24332 32452
rect 24388 32396 28028 32452
rect 28084 32396 28094 32452
rect 31378 32396 31388 32452
rect 31444 32396 31454 32452
rect 31948 32396 33404 32452
rect 33460 32396 33470 32452
rect 34066 32396 34076 32452
rect 34132 32396 36092 32452
rect 36148 32396 36158 32452
rect 31948 32340 32004 32396
rect 8082 32284 8092 32340
rect 8148 32284 8932 32340
rect 8988 32284 11676 32340
rect 11732 32284 11742 32340
rect 14018 32284 14028 32340
rect 14084 32284 14094 32340
rect 14802 32284 14812 32340
rect 14868 32284 16492 32340
rect 16548 32284 18396 32340
rect 18452 32284 18462 32340
rect 19282 32284 19292 32340
rect 19348 32284 23100 32340
rect 23156 32284 23166 32340
rect 24994 32284 25004 32340
rect 25060 32284 25564 32340
rect 25620 32284 26572 32340
rect 26628 32284 29484 32340
rect 29540 32284 29550 32340
rect 30930 32284 30940 32340
rect 30996 32284 31948 32340
rect 32004 32284 32014 32340
rect 32274 32284 32284 32340
rect 32340 32284 35644 32340
rect 35700 32284 35710 32340
rect 36652 32228 36708 32732
rect 37650 32396 37660 32452
rect 37716 32396 37996 32452
rect 38052 32396 38062 32452
rect 9332 32172 9342 32228
rect 9398 32172 10332 32228
rect 10388 32172 10398 32228
rect 10658 32172 10668 32228
rect 10724 32172 10734 32228
rect 21746 32172 21756 32228
rect 21812 32172 22764 32228
rect 22820 32172 22830 32228
rect 36642 32172 36652 32228
rect 36708 32172 36718 32228
rect 5864 32116 5874 32172
rect 5930 32116 5978 32172
rect 6034 32116 6082 32172
rect 6138 32116 6148 32172
rect 10098 32060 10108 32116
rect 10164 32060 10444 32116
rect 10500 32060 10510 32116
rect 4274 31948 4284 32004
rect 4340 31948 8204 32004
rect 8260 31948 8270 32004
rect 10668 31892 10724 32172
rect 15188 32116 15198 32172
rect 15254 32116 15302 32172
rect 15358 32116 15406 32172
rect 15462 32116 15472 32172
rect 24512 32116 24522 32172
rect 24578 32116 24626 32172
rect 24682 32116 24730 32172
rect 24786 32116 24796 32172
rect 33836 32116 33846 32172
rect 33902 32116 33950 32172
rect 34006 32116 34054 32172
rect 34110 32116 34120 32172
rect 15586 32060 15596 32116
rect 15652 32060 17500 32116
rect 17556 32060 17566 32116
rect 18834 32060 18844 32116
rect 18900 32060 20076 32116
rect 20132 32060 20142 32116
rect 28130 32060 28140 32116
rect 28196 32060 30828 32116
rect 30884 32060 30894 32116
rect 35858 32060 35868 32116
rect 35924 32060 36204 32116
rect 36260 32060 36540 32116
rect 36596 32060 36606 32116
rect 17826 31948 17836 32004
rect 17892 31948 21532 32004
rect 21588 31948 21598 32004
rect 22362 31948 22372 32004
rect 22428 31948 23324 32004
rect 23380 31948 23390 32004
rect 23986 31948 23996 32004
rect 24052 31948 24108 32004
rect 24164 31948 24174 32004
rect 30370 31948 30380 32004
rect 30436 31948 31724 32004
rect 31780 31948 34300 32004
rect 34356 31948 34366 32004
rect 19964 31892 20020 31948
rect 2482 31836 2492 31892
rect 2548 31836 5180 31892
rect 5236 31836 5404 31892
rect 5460 31836 9100 31892
rect 9156 31836 9166 31892
rect 10668 31836 11956 31892
rect 12674 31836 12684 31892
rect 12740 31836 14028 31892
rect 14084 31836 14094 31892
rect 14998 31836 15036 31892
rect 15092 31836 15102 31892
rect 15810 31836 15820 31892
rect 15876 31836 16380 31892
rect 16436 31836 17500 31892
rect 17556 31836 19740 31892
rect 19796 31836 19806 31892
rect 19954 31836 19964 31892
rect 20020 31836 20030 31892
rect 35186 31836 35196 31892
rect 35252 31836 35924 31892
rect 35980 31836 35990 31892
rect 4610 31724 4620 31780
rect 4676 31724 5068 31780
rect 5124 31724 5134 31780
rect 7988 31724 7998 31780
rect 8054 31724 10556 31780
rect 10612 31724 10622 31780
rect 7074 31612 7084 31668
rect 7140 31612 8428 31668
rect 8484 31612 8494 31668
rect 11900 31556 11956 31836
rect 12114 31724 12124 31780
rect 12180 31724 13692 31780
rect 13748 31724 14924 31780
rect 14980 31724 14990 31780
rect 22642 31724 22652 31780
rect 22708 31724 23772 31780
rect 23828 31724 23838 31780
rect 31490 31724 31500 31780
rect 31556 31724 35420 31780
rect 35476 31724 35486 31780
rect 39200 31668 40000 31696
rect 12786 31612 12796 31668
rect 12852 31612 13804 31668
rect 13860 31612 13870 31668
rect 14476 31612 22092 31668
rect 22148 31612 22158 31668
rect 37426 31612 37436 31668
rect 37492 31612 40000 31668
rect 14476 31556 14532 31612
rect 39200 31584 40000 31612
rect 10042 31500 10052 31556
rect 10108 31500 11508 31556
rect 11564 31500 11574 31556
rect 11900 31500 12684 31556
rect 12740 31500 13468 31556
rect 13524 31500 14364 31556
rect 14420 31500 14532 31556
rect 14690 31500 14700 31556
rect 14756 31500 15708 31556
rect 15764 31500 15774 31556
rect 20626 31500 20636 31556
rect 20692 31500 22316 31556
rect 22372 31500 23436 31556
rect 23492 31500 23502 31556
rect 4274 31388 4284 31444
rect 4340 31388 6580 31444
rect 6636 31388 6646 31444
rect 14466 31388 14476 31444
rect 14532 31388 15204 31444
rect 15260 31388 15270 31444
rect 37090 31388 37100 31444
rect 37212 31388 37222 31444
rect 10526 31332 10536 31388
rect 10592 31332 10640 31388
rect 10696 31332 10744 31388
rect 10800 31332 10810 31388
rect 19850 31332 19860 31388
rect 19916 31332 19964 31388
rect 20020 31332 20068 31388
rect 20124 31332 20134 31388
rect 29174 31332 29184 31388
rect 29240 31332 29288 31388
rect 29344 31332 29392 31388
rect 29448 31332 29458 31388
rect 38498 31332 38508 31388
rect 38564 31332 38612 31388
rect 38668 31332 38716 31388
rect 38772 31332 38782 31388
rect 9650 31276 9660 31332
rect 9716 31276 10332 31332
rect 10388 31276 10398 31332
rect 10892 31276 14588 31332
rect 14644 31276 14654 31332
rect 10892 31220 10948 31276
rect 5058 31164 5068 31220
rect 5124 31164 6300 31220
rect 6356 31164 6366 31220
rect 10220 31164 10948 31220
rect 11648 31164 11658 31220
rect 11714 31164 13580 31220
rect 13636 31164 13646 31220
rect 13794 31164 13804 31220
rect 13860 31164 14476 31220
rect 14532 31164 14542 31220
rect 16930 31164 16940 31220
rect 16996 31164 17836 31220
rect 17892 31164 19516 31220
rect 19572 31164 19582 31220
rect 19842 31164 19852 31220
rect 19908 31164 20860 31220
rect 20916 31164 20926 31220
rect 26114 31164 26124 31220
rect 26180 31164 26796 31220
rect 26852 31164 26862 31220
rect 32162 31164 32172 31220
rect 32228 31164 33162 31220
rect 33218 31164 33228 31220
rect 35746 31164 35756 31220
rect 35812 31164 37212 31220
rect 37268 31164 37278 31220
rect 1978 31052 1988 31108
rect 2044 31052 5740 31108
rect 5796 31052 7756 31108
rect 7812 31052 7822 31108
rect 10220 30996 10276 31164
rect 13010 31052 13020 31108
rect 13076 31052 15540 31108
rect 15596 31052 15606 31108
rect 20066 31052 20076 31108
rect 20132 31052 20972 31108
rect 21028 31052 21038 31108
rect 23650 31052 23660 31108
rect 23716 31052 25452 31108
rect 25508 31052 27020 31108
rect 27076 31052 27086 31108
rect 27692 31052 30716 31108
rect 30772 31052 30782 31108
rect 32274 31052 32284 31108
rect 32340 31052 37324 31108
rect 37380 31052 37390 31108
rect 37622 31052 37660 31108
rect 37716 31052 37726 31108
rect 27692 30996 27748 31052
rect 3042 30940 3052 30996
rect 3108 30940 5628 30996
rect 5684 30940 5694 30996
rect 7298 30940 7308 30996
rect 7364 30940 8764 30996
rect 8820 30940 10276 30996
rect 14914 30940 14924 30996
rect 14980 30940 16940 30996
rect 16996 30940 17006 30996
rect 19506 30940 19516 30996
rect 19572 30940 20188 30996
rect 20244 30940 20254 30996
rect 22866 30940 22876 30996
rect 22932 30940 23772 30996
rect 23828 30940 23838 30996
rect 24098 30940 24108 30996
rect 24164 30940 26460 30996
rect 26516 30940 26526 30996
rect 26674 30940 26684 30996
rect 26740 30940 27748 30996
rect 27906 30940 27916 30996
rect 27972 30940 29036 30996
rect 29092 30940 29102 30996
rect 33394 30940 33404 30996
rect 33460 30940 36988 30996
rect 37044 30940 38220 30996
rect 38276 30940 38286 30996
rect 10220 30884 10276 30940
rect 2724 30828 2734 30884
rect 2790 30828 6076 30884
rect 6132 30828 6142 30884
rect 10210 30828 10220 30884
rect 10276 30828 10286 30884
rect 24714 30828 24724 30884
rect 24780 30828 25564 30884
rect 25620 30828 28028 30884
rect 28084 30828 28094 30884
rect 33898 30828 33908 30884
rect 33964 30828 34412 30884
rect 34468 30828 34478 30884
rect 35074 30828 35084 30884
rect 35140 30828 37660 30884
rect 37716 30828 37726 30884
rect 19954 30716 19964 30772
rect 20020 30716 21028 30772
rect 21084 30716 23996 30772
rect 24052 30716 26684 30772
rect 26740 30716 26750 30772
rect 28690 30716 28700 30772
rect 28756 30716 33404 30772
rect 33460 30716 33470 30772
rect 28700 30660 28756 30716
rect 13514 30604 13524 30660
rect 13580 30604 14364 30660
rect 14420 30604 15036 30660
rect 15092 30604 15102 30660
rect 16276 30604 16286 30660
rect 16342 30604 21420 30660
rect 21476 30604 21486 30660
rect 24210 30604 24220 30660
rect 24276 30604 24286 30660
rect 27066 30604 27076 30660
rect 27132 30604 28756 30660
rect 5864 30548 5874 30604
rect 5930 30548 5978 30604
rect 6034 30548 6082 30604
rect 6138 30548 6148 30604
rect 15188 30548 15198 30604
rect 15254 30548 15302 30604
rect 15358 30548 15406 30604
rect 15462 30548 15472 30604
rect 12198 30492 12236 30548
rect 12292 30492 12302 30548
rect 13346 30492 13356 30548
rect 13412 30492 14196 30548
rect 14252 30492 15036 30548
rect 15092 30492 15102 30548
rect 20178 30492 20188 30548
rect 20244 30492 20636 30548
rect 20692 30492 21532 30548
rect 21588 30492 21598 30548
rect 24220 30436 24276 30604
rect 24512 30548 24522 30604
rect 24578 30548 24626 30604
rect 24682 30548 24730 30604
rect 24786 30548 24796 30604
rect 33836 30548 33846 30604
rect 33902 30548 33950 30604
rect 34006 30548 34054 30604
rect 34110 30548 34120 30604
rect 24882 30492 24892 30548
rect 24948 30492 24958 30548
rect 15250 30380 15260 30436
rect 15316 30380 15932 30436
rect 15988 30380 16772 30436
rect 16828 30380 16838 30436
rect 20738 30380 20748 30436
rect 20804 30380 21700 30436
rect 21756 30380 22540 30436
rect 22596 30380 22606 30436
rect 24220 30380 24668 30436
rect 24724 30380 24734 30436
rect 2034 30268 2044 30324
rect 2100 30268 2380 30324
rect 2436 30268 2446 30324
rect 2612 30268 2622 30324
rect 2678 30268 4060 30324
rect 4116 30268 4126 30324
rect 9762 30268 9772 30324
rect 9828 30268 11900 30324
rect 11956 30268 11966 30324
rect 14932 30268 14942 30324
rect 14998 30268 16604 30324
rect 16660 30268 16670 30324
rect 17948 30268 22988 30324
rect 23044 30268 23054 30324
rect 1866 30156 1876 30212
rect 1932 30156 6748 30212
rect 6804 30156 7532 30212
rect 7588 30156 7598 30212
rect 7764 30156 7774 30212
rect 7830 30156 8988 30212
rect 9044 30156 9054 30212
rect 12226 30156 12236 30212
rect 12292 30156 13524 30212
rect 13580 30156 13590 30212
rect 15474 30156 15484 30212
rect 15540 30156 16772 30212
rect 16930 30156 16940 30212
rect 16996 30156 17612 30212
rect 17668 30156 17678 30212
rect 16716 30100 16772 30156
rect 17948 30100 18004 30268
rect 24892 30212 24948 30492
rect 26450 30268 26460 30324
rect 26516 30268 32620 30324
rect 32676 30268 32686 30324
rect 36026 30268 36036 30324
rect 36092 30268 36540 30324
rect 36596 30268 36606 30324
rect 19618 30156 19628 30212
rect 19684 30156 20188 30212
rect 20244 30156 20254 30212
rect 20402 30156 20412 30212
rect 20468 30156 21420 30212
rect 21476 30156 21486 30212
rect 23762 30156 23772 30212
rect 23828 30156 24332 30212
rect 24388 30156 26012 30212
rect 26068 30156 26078 30212
rect 29474 30156 29484 30212
rect 29540 30156 29596 30212
rect 29652 30156 29662 30212
rect 29866 30156 29876 30212
rect 29932 30156 37156 30212
rect 37212 30156 37222 30212
rect 7634 30044 7644 30100
rect 7700 30044 8540 30100
rect 8596 30044 8606 30100
rect 8754 30044 8764 30100
rect 8820 30044 9548 30100
rect 9604 30044 9614 30100
rect 10210 30044 10220 30100
rect 10276 30044 12572 30100
rect 12628 30044 12638 30100
rect 14018 30044 14028 30100
rect 14084 30044 14812 30100
rect 14868 30044 14878 30100
rect 16716 30044 18004 30100
rect 26114 30044 26124 30100
rect 26180 30044 32396 30100
rect 32452 30044 33236 30100
rect 33292 30044 33302 30100
rect 34738 30044 34748 30100
rect 34804 30044 37902 30100
rect 37958 30044 37968 30100
rect 14812 29988 14868 30044
rect 11218 29932 11228 29988
rect 11284 29932 11676 29988
rect 11732 29932 12124 29988
rect 12180 29932 13300 29988
rect 14812 29932 16156 29988
rect 16212 29932 23548 29988
rect 23604 29932 23614 29988
rect 32050 29932 32060 29988
rect 32116 29932 34188 29988
rect 34244 29932 34254 29988
rect 34402 29932 34412 29988
rect 34468 29932 37660 29988
rect 37716 29932 37726 29988
rect 13244 29876 13300 29932
rect 10994 29820 11004 29876
rect 11060 29820 12908 29876
rect 12964 29820 12974 29876
rect 13234 29820 13244 29876
rect 13300 29820 15372 29876
rect 15428 29820 15438 29876
rect 15558 29820 15596 29876
rect 15652 29820 16268 29876
rect 16324 29820 16334 29876
rect 21186 29820 21196 29876
rect 21252 29820 25004 29876
rect 25060 29820 25070 29876
rect 10526 29764 10536 29820
rect 10592 29764 10640 29820
rect 10696 29764 10744 29820
rect 10800 29764 10810 29820
rect 11004 29652 11060 29820
rect 19850 29764 19860 29820
rect 19916 29764 19964 29820
rect 20020 29764 20068 29820
rect 20124 29764 20134 29820
rect 29174 29764 29184 29820
rect 29240 29764 29288 29820
rect 29344 29764 29392 29820
rect 29448 29764 29458 29820
rect 38498 29764 38508 29820
rect 38564 29764 38612 29820
rect 38668 29764 38716 29820
rect 38772 29764 38782 29820
rect 11834 29708 11844 29764
rect 11900 29708 12404 29764
rect 12460 29708 14364 29764
rect 14420 29708 14430 29764
rect 32498 29708 32508 29764
rect 32564 29708 36316 29764
rect 36372 29708 36382 29764
rect 7970 29596 7980 29652
rect 8036 29596 9548 29652
rect 9604 29596 11060 29652
rect 12114 29596 12124 29652
rect 12180 29596 12684 29652
rect 12740 29596 12750 29652
rect 23762 29596 23772 29652
rect 23828 29596 24556 29652
rect 24612 29596 24622 29652
rect 28018 29596 28028 29652
rect 28084 29596 28364 29652
rect 28420 29596 29092 29652
rect 29148 29596 29158 29652
rect 30902 29596 30940 29652
rect 30996 29596 31006 29652
rect 32050 29596 32060 29652
rect 32116 29596 37100 29652
rect 37156 29596 37166 29652
rect 9874 29484 9884 29540
rect 9940 29484 12236 29540
rect 12292 29484 12302 29540
rect 18274 29484 18284 29540
rect 18340 29484 19908 29540
rect 19964 29484 19974 29540
rect 20850 29484 20860 29540
rect 20916 29484 21084 29540
rect 21140 29484 21150 29540
rect 25498 29484 25508 29540
rect 25564 29484 25676 29540
rect 25732 29484 26124 29540
rect 26180 29484 26190 29540
rect 29250 29484 29260 29540
rect 29316 29484 29596 29540
rect 29652 29484 29662 29540
rect 4946 29372 4956 29428
rect 5012 29372 9772 29428
rect 9828 29372 9838 29428
rect 10770 29372 10780 29428
rect 10836 29372 13356 29428
rect 13412 29372 13422 29428
rect 18386 29372 18396 29428
rect 18452 29372 19516 29428
rect 19572 29372 19582 29428
rect 21186 29372 21196 29428
rect 21252 29372 22708 29428
rect 22764 29372 22774 29428
rect 29362 29372 29372 29428
rect 29428 29372 30380 29428
rect 30436 29372 30446 29428
rect 38322 29372 38332 29428
rect 38388 29372 39284 29428
rect 7298 29260 7308 29316
rect 7364 29260 9660 29316
rect 9716 29260 10108 29316
rect 10164 29260 10174 29316
rect 19618 29260 19628 29316
rect 19684 29260 20860 29316
rect 20916 29260 20926 29316
rect 24714 29260 24724 29316
rect 24780 29260 27916 29316
rect 27972 29260 28140 29316
rect 28196 29260 28206 29316
rect 28466 29260 28476 29316
rect 28532 29260 29428 29316
rect 29372 29204 29428 29260
rect 3042 29148 3052 29204
rect 3108 29148 3612 29204
rect 3668 29148 3678 29204
rect 8530 29148 8540 29204
rect 8596 29148 9996 29204
rect 10052 29148 10444 29204
rect 10500 29148 10510 29204
rect 19394 29148 19404 29204
rect 19460 29148 19628 29204
rect 19684 29148 19694 29204
rect 25778 29148 25788 29204
rect 25844 29148 26012 29204
rect 26068 29148 26796 29204
rect 26852 29148 28756 29204
rect 28812 29148 29036 29204
rect 29092 29148 29102 29204
rect 29362 29148 29372 29204
rect 29428 29148 31612 29204
rect 31668 29148 34412 29204
rect 34468 29148 34478 29204
rect 34962 29148 34972 29204
rect 35028 29148 36764 29204
rect 36820 29148 36830 29204
rect 6570 29036 6580 29092
rect 6636 29036 10892 29092
rect 10948 29036 11452 29092
rect 11508 29036 11518 29092
rect 18666 29036 18676 29092
rect 18732 29036 19516 29092
rect 19572 29036 19582 29092
rect 28466 29036 28476 29092
rect 28532 29036 32844 29092
rect 32900 29036 32910 29092
rect 5864 28980 5874 29036
rect 5930 28980 5978 29036
rect 6034 28980 6082 29036
rect 6138 28980 6148 29036
rect 15188 28980 15198 29036
rect 15254 28980 15302 29036
rect 15358 28980 15406 29036
rect 15462 28980 15472 29036
rect 24512 28980 24522 29036
rect 24578 28980 24626 29036
rect 24682 28980 24730 29036
rect 24786 28980 24796 29036
rect 28812 28980 28868 29036
rect 33836 28980 33846 29036
rect 33902 28980 33950 29036
rect 34006 28980 34054 29036
rect 34110 28980 34120 29036
rect 39228 28980 39284 29372
rect 8754 28924 8764 28980
rect 8820 28924 9436 28980
rect 9492 28924 9502 28980
rect 15596 28924 23100 28980
rect 23156 28924 23166 28980
rect 28802 28924 28812 28980
rect 28868 28924 28878 28980
rect 30594 28924 30604 28980
rect 30660 28924 32060 28980
rect 32116 28924 32126 28980
rect 39004 28924 39284 28980
rect 15596 28868 15652 28924
rect 7970 28812 7980 28868
rect 8036 28812 8652 28868
rect 8708 28812 8718 28868
rect 9202 28812 9212 28868
rect 9268 28812 10892 28868
rect 10948 28812 10958 28868
rect 11666 28812 11676 28868
rect 11732 28812 12460 28868
rect 12516 28812 12740 28868
rect 12796 28812 13636 28868
rect 13692 28812 15652 28868
rect 15810 28812 15820 28868
rect 15876 28812 21532 28868
rect 21588 28812 21598 28868
rect 22250 28812 22260 28868
rect 22316 28812 23436 28868
rect 23492 28812 23502 28868
rect 24658 28812 24668 28868
rect 24724 28812 25900 28868
rect 25956 28812 25966 28868
rect 29586 28812 29596 28868
rect 29652 28812 32844 28868
rect 32900 28812 32910 28868
rect 39004 28756 39060 28924
rect 39200 28756 40000 28784
rect 7634 28700 7644 28756
rect 7700 28700 9156 28756
rect 21074 28700 21084 28756
rect 21140 28700 22764 28756
rect 22820 28700 22830 28756
rect 23650 28700 23660 28756
rect 23716 28700 24500 28756
rect 24556 28700 24566 28756
rect 24770 28700 24780 28756
rect 24836 28700 26964 28756
rect 32722 28700 32732 28756
rect 32788 28700 36988 28756
rect 37044 28700 37054 28756
rect 39004 28700 40000 28756
rect 9100 28644 9156 28700
rect 24780 28644 24836 28700
rect 8194 28588 8204 28644
rect 8260 28588 8876 28644
rect 8932 28588 8942 28644
rect 9100 28588 9716 28644
rect 9772 28588 10444 28644
rect 10500 28588 10510 28644
rect 16594 28588 16604 28644
rect 16660 28588 17388 28644
rect 17444 28588 17454 28644
rect 19114 28588 19124 28644
rect 19180 28588 20412 28644
rect 20468 28588 20478 28644
rect 23538 28588 23548 28644
rect 23604 28588 24836 28644
rect 17154 28476 17164 28532
rect 17220 28476 18396 28532
rect 18452 28476 18462 28532
rect 21858 28476 21868 28532
rect 21924 28476 21934 28532
rect 18396 28420 18452 28476
rect 21868 28420 21924 28476
rect 10770 28364 10780 28420
rect 10836 28364 11900 28420
rect 11956 28364 11966 28420
rect 16482 28364 16492 28420
rect 16548 28364 17052 28420
rect 17108 28364 17388 28420
rect 17444 28364 17454 28420
rect 18396 28364 22148 28420
rect 22204 28364 22214 28420
rect 23090 28364 23100 28420
rect 23156 28364 23492 28420
rect 23548 28364 25116 28420
rect 25172 28364 25182 28420
rect 26908 28364 26964 28700
rect 39200 28672 40000 28700
rect 29586 28588 29596 28644
rect 29652 28588 32060 28644
rect 32116 28588 32900 28644
rect 33058 28588 33068 28644
rect 33124 28588 37436 28644
rect 37492 28588 37502 28644
rect 32844 28532 32900 28588
rect 30370 28476 30380 28532
rect 30436 28476 32302 28532
rect 32358 28476 32368 28532
rect 32844 28476 33740 28532
rect 33796 28476 33806 28532
rect 27020 28364 27030 28420
rect 32162 28364 32172 28420
rect 32228 28364 37660 28420
rect 37716 28364 37726 28420
rect 10526 28196 10536 28252
rect 10592 28196 10640 28252
rect 10696 28196 10744 28252
rect 10800 28196 10810 28252
rect 19850 28196 19860 28252
rect 19916 28196 19964 28252
rect 20020 28196 20068 28252
rect 20124 28196 20134 28252
rect 29174 28196 29184 28252
rect 29240 28196 29288 28252
rect 29344 28196 29392 28252
rect 29448 28196 29458 28252
rect 38498 28196 38508 28252
rect 38564 28196 38612 28252
rect 38668 28196 38716 28252
rect 38772 28196 38782 28252
rect 13346 28140 13356 28196
rect 13412 28140 14588 28196
rect 14644 28140 17388 28196
rect 17444 28140 17454 28196
rect 18050 28140 18060 28196
rect 18116 28140 18732 28196
rect 18788 28140 18956 28196
rect 19012 28140 19022 28196
rect 18274 28028 18284 28084
rect 18340 28028 19404 28084
rect 19460 28028 20972 28084
rect 21028 28028 21038 28084
rect 21718 28028 21756 28084
rect 21812 28028 21822 28084
rect 26562 28028 26572 28084
rect 26628 28028 28140 28084
rect 28196 28028 28206 28084
rect 28578 28028 28588 28084
rect 28644 28028 34860 28084
rect 34916 28028 34926 28084
rect 10780 27916 12124 27972
rect 12180 27916 12190 27972
rect 20066 27916 20076 27972
rect 20132 27916 21308 27972
rect 21364 27916 21374 27972
rect 24658 27916 24668 27972
rect 24724 27916 25583 27972
rect 25639 27916 25649 27972
rect 26124 27916 27132 27972
rect 27188 27916 27198 27972
rect 34178 27916 34188 27972
rect 34244 27916 34468 27972
rect 3266 27804 3276 27860
rect 3332 27804 4844 27860
rect 4900 27804 4910 27860
rect 9818 27804 9828 27860
rect 9884 27804 10724 27860
rect 10780 27804 10836 27916
rect 26124 27860 26180 27916
rect 11498 27804 11508 27860
rect 11564 27804 16604 27860
rect 16660 27804 17500 27860
rect 17556 27804 17566 27860
rect 17938 27804 17948 27860
rect 18004 27804 19010 27860
rect 19066 27804 19076 27860
rect 19730 27804 19740 27860
rect 19796 27804 20188 27860
rect 20244 27804 20636 27860
rect 20692 27804 20702 27860
rect 24546 27804 24556 27860
rect 24612 27804 25004 27860
rect 25060 27804 25070 27860
rect 25330 27804 25340 27860
rect 25396 27804 26180 27860
rect 26450 27804 26460 27860
rect 26516 27804 28644 27860
rect 28700 27804 28710 27860
rect 29586 27804 29596 27860
rect 29652 27804 30492 27860
rect 30548 27804 30558 27860
rect 31602 27804 31612 27860
rect 31724 27804 31734 27860
rect 26460 27748 26516 27804
rect 20738 27692 20748 27748
rect 20804 27692 21532 27748
rect 21588 27692 21598 27748
rect 25666 27692 25676 27748
rect 25732 27692 26516 27748
rect 29642 27692 29652 27748
rect 29708 27692 30156 27748
rect 30212 27692 30222 27748
rect 34412 27636 34468 27916
rect 3602 27580 3612 27636
rect 3668 27580 4228 27636
rect 4284 27580 14476 27636
rect 14532 27580 14542 27636
rect 18946 27580 18956 27636
rect 19012 27580 19628 27636
rect 19684 27580 19694 27636
rect 21644 27580 27356 27636
rect 27412 27580 27422 27636
rect 30706 27580 30716 27636
rect 30772 27580 30940 27636
rect 30996 27580 31006 27636
rect 34402 27580 34412 27636
rect 34468 27580 34478 27636
rect 21644 27524 21700 27580
rect 17490 27468 17500 27524
rect 17556 27468 19572 27524
rect 21634 27468 21644 27524
rect 21700 27468 21710 27524
rect 5864 27412 5874 27468
rect 5930 27412 5978 27468
rect 6034 27412 6082 27468
rect 6138 27412 6148 27468
rect 15188 27412 15198 27468
rect 15254 27412 15302 27468
rect 15358 27412 15406 27468
rect 15462 27412 15472 27468
rect 19516 27412 19572 27468
rect 24512 27412 24522 27468
rect 24578 27412 24626 27468
rect 24682 27412 24730 27468
rect 24786 27412 24796 27468
rect 33836 27412 33846 27468
rect 33902 27412 33950 27468
rect 34006 27412 34054 27468
rect 34110 27412 34120 27468
rect 10882 27356 10892 27412
rect 10948 27356 11564 27412
rect 11620 27356 11630 27412
rect 16594 27356 16604 27412
rect 16660 27356 18396 27412
rect 18452 27356 19292 27412
rect 19348 27356 19358 27412
rect 19516 27356 24050 27412
rect 24106 27356 24116 27412
rect 25106 27356 25116 27412
rect 25172 27356 26348 27412
rect 26404 27356 27860 27412
rect 27916 27356 27926 27412
rect 14000 27244 14010 27300
rect 14066 27244 16716 27300
rect 16772 27244 16782 27300
rect 24994 27244 25004 27300
rect 25060 27244 26012 27300
rect 26068 27244 26078 27300
rect 31154 27244 31164 27300
rect 31220 27244 32396 27300
rect 32452 27244 32462 27300
rect 9090 27132 9100 27188
rect 9156 27132 9996 27188
rect 10052 27132 12124 27188
rect 12180 27132 12852 27188
rect 12908 27132 13356 27188
rect 13412 27132 13636 27188
rect 13692 27132 17276 27188
rect 17332 27132 17342 27188
rect 21074 27132 21084 27188
rect 21140 27132 21420 27188
rect 21476 27132 21486 27188
rect 25554 27132 25564 27188
rect 25620 27132 26236 27188
rect 26292 27132 26302 27188
rect 31266 27132 31276 27188
rect 31332 27132 32508 27188
rect 32564 27132 32574 27188
rect 8866 27020 8876 27076
rect 8932 27020 9716 27076
rect 9772 27020 9782 27076
rect 15092 27020 15260 27076
rect 15316 27020 15326 27076
rect 15418 27020 15428 27076
rect 15484 27020 15820 27076
rect 15876 27020 15886 27076
rect 16164 27020 16174 27076
rect 16230 27020 18844 27076
rect 18900 27020 18910 27076
rect 19394 27020 19404 27076
rect 19460 27020 19516 27076
rect 19572 27020 19582 27076
rect 20794 27020 20804 27076
rect 20860 27020 21644 27076
rect 21700 27020 21710 27076
rect 23874 27020 23884 27076
rect 23940 27020 26516 27076
rect 26572 27020 26582 27076
rect 27346 27020 27356 27076
rect 27412 27020 28252 27076
rect 28308 27020 28318 27076
rect 30818 27020 30828 27076
rect 30884 27020 31500 27076
rect 31556 27020 31566 27076
rect 36474 27020 36484 27076
rect 36540 27020 38332 27076
rect 38388 27020 38398 27076
rect 15092 26964 15148 27020
rect 8754 26908 8764 26964
rect 8820 26908 13804 26964
rect 13860 26908 14924 26964
rect 14980 26908 15148 26964
rect 17378 26908 17388 26964
rect 17444 26908 17948 26964
rect 18004 26908 18014 26964
rect 19058 26908 19068 26964
rect 19124 26908 24220 26964
rect 24276 26908 25004 26964
rect 25060 26908 25070 26964
rect 25228 26908 25564 26964
rect 25620 26908 25630 26964
rect 25890 26908 25900 26964
rect 25956 26908 27244 26964
rect 27300 26908 27310 26964
rect 31042 26908 31052 26964
rect 31108 26908 32060 26964
rect 32116 26908 32126 26964
rect 36866 26908 36876 26964
rect 36932 26908 37996 26964
rect 38052 26908 38062 26964
rect 25228 26852 25284 26908
rect 10882 26796 10892 26852
rect 10948 26796 11788 26852
rect 11844 26796 11854 26852
rect 19170 26796 19180 26852
rect 19236 26796 20524 26852
rect 20580 26796 20590 26852
rect 24882 26796 24892 26852
rect 24948 26796 25284 26852
rect 31266 26796 31276 26852
rect 31332 26796 31500 26852
rect 31556 26796 31566 26852
rect 30594 26684 30604 26740
rect 30660 26684 31612 26740
rect 31668 26684 31678 26740
rect 10526 26628 10536 26684
rect 10592 26628 10640 26684
rect 10696 26628 10744 26684
rect 10800 26628 10810 26684
rect 19850 26628 19860 26684
rect 19916 26628 19964 26684
rect 20020 26628 20068 26684
rect 20124 26628 20134 26684
rect 29174 26628 29184 26684
rect 29240 26628 29288 26684
rect 29344 26628 29392 26684
rect 29448 26628 29458 26684
rect 38498 26628 38508 26684
rect 38564 26628 38612 26684
rect 38668 26628 38716 26684
rect 38772 26628 38782 26684
rect 19562 26572 19572 26628
rect 19684 26572 19694 26628
rect 20262 26572 20300 26628
rect 20356 26572 20366 26628
rect 23202 26572 23212 26628
rect 23268 26572 25676 26628
rect 25732 26572 25742 26628
rect 11274 26460 11284 26516
rect 11340 26460 11564 26516
rect 11620 26460 21028 26516
rect 24994 26460 25004 26516
rect 25060 26460 25340 26516
rect 25396 26460 27188 26516
rect 27244 26460 28140 26516
rect 28196 26460 28206 26516
rect 20972 26404 21028 26460
rect 3098 26348 3108 26404
rect 3164 26348 4956 26404
rect 5012 26348 5022 26404
rect 10434 26348 10444 26404
rect 10500 26348 11452 26404
rect 11508 26348 15820 26404
rect 15876 26348 15886 26404
rect 16818 26348 16828 26404
rect 16884 26348 19852 26404
rect 19908 26348 20356 26404
rect 20514 26348 20524 26404
rect 20580 26348 20748 26404
rect 20804 26348 20814 26404
rect 20972 26348 26908 26404
rect 30314 26348 30324 26404
rect 30380 26348 30940 26404
rect 30996 26348 31006 26404
rect 20300 26292 20356 26348
rect 26852 26292 26908 26348
rect 1698 26236 1708 26292
rect 1764 26236 2940 26292
rect 2996 26236 4060 26292
rect 4116 26236 5516 26292
rect 5572 26236 5582 26292
rect 16370 26236 16380 26292
rect 16436 26236 17276 26292
rect 17332 26236 17342 26292
rect 18722 26236 18732 26292
rect 18788 26236 20076 26292
rect 20132 26236 20142 26292
rect 20300 26236 24612 26292
rect 26852 26236 28196 26292
rect 28252 26236 28476 26292
rect 28532 26236 28542 26292
rect 24556 26180 24612 26236
rect 15922 26124 15932 26180
rect 15988 26124 23772 26180
rect 23828 26124 23838 26180
rect 24546 26124 24556 26180
rect 24612 26124 27020 26180
rect 27076 26124 27086 26180
rect 28354 26124 28364 26180
rect 28420 26124 31724 26180
rect 31780 26124 32396 26180
rect 32452 26124 32462 26180
rect 9650 26012 9660 26068
rect 9716 26012 10164 26068
rect 10220 26012 12348 26068
rect 12404 26012 14980 26068
rect 15036 26012 22204 26068
rect 22260 26012 25788 26068
rect 25844 26012 25854 26068
rect 31490 26012 31500 26068
rect 31556 26012 33628 26068
rect 33684 26012 33694 26068
rect 17612 25900 19180 25956
rect 19236 25900 19516 25956
rect 19572 25900 19582 25956
rect 31154 25900 31164 25956
rect 31220 25900 31836 25956
rect 31892 25900 31902 25956
rect 5864 25844 5874 25900
rect 5930 25844 5978 25900
rect 6034 25844 6082 25900
rect 6138 25844 6148 25900
rect 15188 25844 15198 25900
rect 15254 25844 15302 25900
rect 15358 25844 15406 25900
rect 15462 25844 15472 25900
rect 17612 25844 17668 25900
rect 24512 25844 24522 25900
rect 24578 25844 24626 25900
rect 24682 25844 24730 25900
rect 24786 25844 24796 25900
rect 33836 25844 33846 25900
rect 33902 25844 33950 25900
rect 34006 25844 34054 25900
rect 34110 25844 34120 25900
rect 39200 25844 40000 25872
rect 17602 25788 17612 25844
rect 17668 25788 17678 25844
rect 19366 25788 19404 25844
rect 19460 25788 19470 25844
rect 38322 25788 38332 25844
rect 38388 25788 40000 25844
rect 39200 25760 40000 25788
rect 19282 25676 19292 25732
rect 19348 25676 20692 25732
rect 20748 25676 20758 25732
rect 24770 25676 24780 25732
rect 24836 25676 25340 25732
rect 25396 25676 25406 25732
rect 31826 25676 31836 25732
rect 31892 25676 34412 25732
rect 34468 25676 34478 25732
rect 6178 25564 6188 25620
rect 6244 25564 6972 25620
rect 7028 25564 7038 25620
rect 15810 25564 15820 25620
rect 15876 25564 20300 25620
rect 20356 25564 20366 25620
rect 23538 25564 23548 25620
rect 23604 25564 23772 25620
rect 23828 25564 23838 25620
rect 27906 25564 27916 25620
rect 27972 25564 28588 25620
rect 28644 25564 28654 25620
rect 6682 25452 6692 25508
rect 6748 25452 7196 25508
rect 7252 25452 8316 25508
rect 8372 25452 8382 25508
rect 10994 25452 11004 25508
rect 11060 25452 11788 25508
rect 11844 25452 11854 25508
rect 12450 25452 12460 25508
rect 12516 25452 14140 25508
rect 14196 25452 15260 25508
rect 15316 25452 16380 25508
rect 16436 25452 16446 25508
rect 18610 25452 18620 25508
rect 18676 25452 20076 25508
rect 20132 25452 20142 25508
rect 24210 25452 24220 25508
rect 24276 25452 25004 25508
rect 25060 25452 26068 25508
rect 26124 25452 26134 25508
rect 29418 25452 29428 25508
rect 29484 25452 29932 25508
rect 29988 25452 33516 25508
rect 33572 25452 33582 25508
rect 35410 25452 35420 25508
rect 35476 25452 35756 25508
rect 35812 25452 35822 25508
rect 19292 25340 20524 25396
rect 20580 25340 20590 25396
rect 23538 25340 23548 25396
rect 23604 25340 24780 25396
rect 24836 25340 24846 25396
rect 31490 25340 31500 25396
rect 31556 25340 33852 25396
rect 33908 25340 34692 25396
rect 34748 25340 35364 25396
rect 35420 25340 35430 25396
rect 35522 25340 35532 25396
rect 35588 25340 35644 25396
rect 35700 25340 35710 25396
rect 19292 25284 19348 25340
rect 2034 25228 2044 25284
rect 2100 25228 2268 25284
rect 2324 25228 4340 25284
rect 4396 25228 4406 25284
rect 4946 25228 4956 25284
rect 5012 25228 5740 25284
rect 5796 25228 5806 25284
rect 11778 25228 11788 25284
rect 11844 25228 13076 25284
rect 13132 25228 13142 25284
rect 18442 25228 18452 25284
rect 18508 25228 18956 25284
rect 19012 25228 19022 25284
rect 19282 25228 19292 25284
rect 19348 25228 19358 25284
rect 19516 25228 19852 25284
rect 19908 25228 19918 25284
rect 20402 25228 20412 25284
rect 20468 25228 21476 25284
rect 21532 25228 21756 25284
rect 21812 25228 23884 25284
rect 23940 25228 23950 25284
rect 28018 25228 28028 25284
rect 28084 25228 30380 25284
rect 30436 25228 31276 25284
rect 31332 25228 31342 25284
rect 31500 25228 31724 25284
rect 31780 25228 32284 25284
rect 32340 25228 34188 25284
rect 34244 25228 34254 25284
rect 10526 25060 10536 25116
rect 10592 25060 10640 25116
rect 10696 25060 10744 25116
rect 10800 25060 10810 25116
rect 3602 25004 3612 25060
rect 3668 25004 4732 25060
rect 4788 25004 4798 25060
rect 3826 24892 3836 24948
rect 3892 24892 5068 24948
rect 5124 24892 5134 24948
rect 19516 24836 19572 25228
rect 31500 25172 31556 25228
rect 25778 25116 25788 25172
rect 25844 25116 26516 25172
rect 26572 25116 26582 25172
rect 30818 25116 30828 25172
rect 30884 25116 31556 25172
rect 19850 25060 19860 25116
rect 19916 25060 19964 25116
rect 20020 25060 20068 25116
rect 20124 25060 20134 25116
rect 29174 25060 29184 25116
rect 29240 25060 29288 25116
rect 29344 25060 29392 25116
rect 29448 25060 29458 25116
rect 38498 25060 38508 25116
rect 38564 25060 38612 25116
rect 38668 25060 38716 25116
rect 38772 25060 38782 25116
rect 29810 25004 29820 25060
rect 29876 25004 32508 25060
rect 32564 25004 35980 25060
rect 36036 25004 36046 25060
rect 24098 24892 24108 24948
rect 24164 24892 29036 24948
rect 29092 24892 29102 24948
rect 31378 24892 31388 24948
rect 31444 24892 31454 24948
rect 31388 24836 31444 24892
rect 3938 24780 3948 24836
rect 4004 24780 5572 24836
rect 5628 24780 5638 24836
rect 18274 24780 18284 24836
rect 18340 24780 19516 24836
rect 19572 24780 19582 24836
rect 30146 24780 30156 24836
rect 30212 24780 33404 24836
rect 33460 24780 33470 24836
rect 35186 24780 35196 24836
rect 35252 24780 36876 24836
rect 36932 24780 36942 24836
rect 37874 24780 37884 24836
rect 37940 24780 38220 24836
rect 38276 24780 38286 24836
rect 37884 24724 37940 24780
rect 4946 24668 4956 24724
rect 5012 24668 7756 24724
rect 7812 24668 12908 24724
rect 12964 24668 12974 24724
rect 17826 24668 17836 24724
rect 17892 24668 18116 24724
rect 18172 24668 18182 24724
rect 19730 24668 19740 24724
rect 19796 24668 20300 24724
rect 20356 24668 20366 24724
rect 21298 24668 21308 24724
rect 21364 24668 24332 24724
rect 24388 24668 24398 24724
rect 26506 24668 26516 24724
rect 26572 24668 29820 24724
rect 29876 24668 30268 24724
rect 30324 24668 30334 24724
rect 31378 24668 31388 24724
rect 31444 24668 32060 24724
rect 32116 24668 32126 24724
rect 34962 24668 34972 24724
rect 35028 24668 37212 24724
rect 37268 24668 37278 24724
rect 37426 24668 37436 24724
rect 37492 24668 37940 24724
rect 6626 24556 6636 24612
rect 6692 24556 8988 24612
rect 9044 24556 9054 24612
rect 20962 24556 20972 24612
rect 21028 24556 22092 24612
rect 22148 24556 22158 24612
rect 31714 24556 31724 24612
rect 31780 24556 32732 24612
rect 32788 24556 32798 24612
rect 36194 24556 36204 24612
rect 36260 24556 37548 24612
rect 37604 24556 37996 24612
rect 38052 24556 38062 24612
rect 38266 24556 38276 24612
rect 38332 24556 39004 24612
rect 39060 24556 39070 24612
rect 7074 24444 7084 24500
rect 7140 24444 8074 24500
rect 8130 24444 8140 24500
rect 13626 24444 13636 24500
rect 13692 24444 14252 24500
rect 14308 24444 15484 24500
rect 15540 24444 15550 24500
rect 19114 24444 19124 24500
rect 19180 24444 20524 24500
rect 20580 24444 20590 24500
rect 31686 24332 31724 24388
rect 31780 24332 31790 24388
rect 5864 24276 5874 24332
rect 5930 24276 5978 24332
rect 6034 24276 6082 24332
rect 6138 24276 6148 24332
rect 15188 24276 15198 24332
rect 15254 24276 15302 24332
rect 15358 24276 15406 24332
rect 15462 24276 15472 24332
rect 24512 24276 24522 24332
rect 24578 24276 24626 24332
rect 24682 24276 24730 24332
rect 24786 24276 24796 24332
rect 33836 24276 33846 24332
rect 33902 24276 33950 24332
rect 34006 24276 34054 24332
rect 34110 24276 34120 24332
rect 18162 24220 18172 24276
rect 18228 24220 24108 24276
rect 24164 24220 24174 24276
rect 12730 24108 12740 24164
rect 12796 24108 13916 24164
rect 13972 24108 15036 24164
rect 15092 24108 15102 24164
rect 23650 24108 23660 24164
rect 23716 24108 23884 24164
rect 23940 24108 23950 24164
rect 29026 24108 29036 24164
rect 29092 24108 29652 24164
rect 29708 24108 34580 24164
rect 34636 24108 35308 24164
rect 35364 24108 37996 24164
rect 38052 24108 38276 24164
rect 38332 24108 38342 24164
rect 14130 23996 14140 24052
rect 14196 23996 24108 24052
rect 24164 23996 24174 24052
rect 29810 23996 29820 24052
rect 29876 23996 30716 24052
rect 30772 23996 31892 24052
rect 35382 23996 35420 24052
rect 35476 23996 35486 24052
rect 35634 23996 35644 24052
rect 35700 23996 35738 24052
rect 31836 23940 31892 23996
rect 12226 23884 12236 23940
rect 12292 23884 13636 23940
rect 13692 23884 13702 23940
rect 17490 23884 17500 23940
rect 17556 23884 19180 23940
rect 19236 23884 19404 23940
rect 19460 23884 19470 23940
rect 20738 23884 20748 23940
rect 20804 23884 21980 23940
rect 22036 23884 22046 23940
rect 27570 23884 27580 23940
rect 27636 23884 28252 23940
rect 28308 23884 29036 23940
rect 29092 23884 29372 23940
rect 29428 23884 29438 23940
rect 30930 23884 30940 23940
rect 30996 23884 31006 23940
rect 31826 23884 31836 23940
rect 31892 23884 35980 23940
rect 36036 23884 36046 23940
rect 36362 23884 36372 23940
rect 36428 23884 37324 23940
rect 37380 23884 37390 23940
rect 9314 23772 9324 23828
rect 9380 23772 10332 23828
rect 10388 23772 13636 23828
rect 18918 23772 18956 23828
rect 19012 23772 19022 23828
rect 13580 23716 13636 23772
rect 4722 23660 4732 23716
rect 4788 23660 5740 23716
rect 5796 23660 5806 23716
rect 11778 23660 11788 23716
rect 11844 23660 12236 23716
rect 12292 23660 12302 23716
rect 13570 23660 13580 23716
rect 13636 23660 13646 23716
rect 17826 23660 17836 23716
rect 17892 23660 19292 23716
rect 19348 23660 23660 23716
rect 23716 23660 23726 23716
rect 10882 23548 10892 23604
rect 10948 23548 18172 23604
rect 18228 23548 18238 23604
rect 18330 23548 18340 23604
rect 18396 23548 18844 23604
rect 18900 23548 18910 23604
rect 10526 23492 10536 23548
rect 10592 23492 10640 23548
rect 10696 23492 10744 23548
rect 10800 23492 10810 23548
rect 19850 23492 19860 23548
rect 19916 23492 19964 23548
rect 20020 23492 20068 23548
rect 20124 23492 20134 23548
rect 29174 23492 29184 23548
rect 29240 23492 29288 23548
rect 29344 23492 29392 23548
rect 29448 23492 29458 23548
rect 28018 23436 28028 23492
rect 28084 23436 28644 23492
rect 28700 23436 28924 23492
rect 28980 23436 28990 23492
rect 2930 23324 2940 23380
rect 2996 23324 4284 23380
rect 4340 23324 4844 23380
rect 4900 23324 5292 23380
rect 5348 23324 5358 23380
rect 9426 23324 9436 23380
rect 9492 23324 11116 23380
rect 11172 23324 11182 23380
rect 11554 23324 11564 23380
rect 11620 23324 12012 23380
rect 12068 23324 13356 23380
rect 13412 23324 15652 23380
rect 15708 23324 15932 23380
rect 15988 23324 15998 23380
rect 16594 23324 16604 23380
rect 16660 23324 17164 23380
rect 17220 23324 17230 23380
rect 17938 23324 17948 23380
rect 18004 23324 22316 23380
rect 22372 23324 22382 23380
rect 27794 23324 27804 23380
rect 27860 23324 30380 23380
rect 30436 23324 30446 23380
rect 6234 23212 6244 23268
rect 6300 23212 6860 23268
rect 6916 23212 7980 23268
rect 8036 23212 8046 23268
rect 10770 23212 10780 23268
rect 10836 23212 11452 23268
rect 11508 23212 11518 23268
rect 18050 23212 18060 23268
rect 18116 23212 20076 23268
rect 20132 23212 23212 23268
rect 23268 23212 23278 23268
rect 6570 23100 6580 23156
rect 6636 23100 7196 23156
rect 7252 23100 7262 23156
rect 9202 23100 9212 23156
rect 9268 23100 9884 23156
rect 9940 23100 11004 23156
rect 11060 23100 11070 23156
rect 16930 23100 16940 23156
rect 16996 23100 19068 23156
rect 19124 23100 20300 23156
rect 20356 23100 20366 23156
rect 22418 23100 22428 23156
rect 22484 23100 23436 23156
rect 23492 23100 23502 23156
rect 26450 23100 26460 23156
rect 26516 23100 27132 23156
rect 27188 23100 27198 23156
rect 4610 22988 4620 23044
rect 4676 22988 5012 23044
rect 5068 22988 6076 23044
rect 6132 22988 8652 23044
rect 8708 22988 8718 23044
rect 10378 22988 10388 23044
rect 10444 22988 10892 23044
rect 10948 22988 10958 23044
rect 14802 22988 14812 23044
rect 14868 22988 16100 23044
rect 16156 22988 16166 23044
rect 27804 22932 27860 23324
rect 30940 23268 30996 23884
rect 34962 23772 34972 23828
rect 35028 23772 37436 23828
rect 37492 23772 37502 23828
rect 31938 23548 31948 23604
rect 32004 23548 32844 23604
rect 32900 23548 32910 23604
rect 35186 23548 35196 23604
rect 35252 23548 35868 23604
rect 35924 23548 37996 23604
rect 38052 23548 38062 23604
rect 38498 23492 38508 23548
rect 38564 23492 38612 23548
rect 38668 23492 38716 23548
rect 38772 23492 38782 23548
rect 32946 23436 32956 23492
rect 33012 23436 37156 23492
rect 37212 23436 37222 23492
rect 31378 23324 31388 23380
rect 31444 23324 34860 23380
rect 34916 23324 34926 23380
rect 30146 23212 30156 23268
rect 30212 23212 30492 23268
rect 30548 23212 34580 23268
rect 34524 23156 34580 23212
rect 31042 23100 31052 23156
rect 31108 23100 31612 23156
rect 31668 23100 31678 23156
rect 34514 23100 34524 23156
rect 34580 23100 35420 23156
rect 35476 23100 35486 23156
rect 39200 22932 40000 22960
rect 8194 22876 8204 22932
rect 8260 22876 9642 22932
rect 9698 22876 9708 22932
rect 14018 22876 14028 22932
rect 14084 22876 15092 22932
rect 15148 22876 15158 22932
rect 25666 22876 25676 22932
rect 25732 22876 27860 22932
rect 31266 22876 31276 22932
rect 31332 22876 32060 22932
rect 32116 22876 32126 22932
rect 32274 22876 32284 22932
rect 32340 22876 34860 22932
rect 34916 22876 35644 22932
rect 35700 22876 35710 22932
rect 38322 22876 38332 22932
rect 38388 22876 40000 22932
rect 39200 22848 40000 22876
rect 32386 22764 32396 22820
rect 32452 22764 32732 22820
rect 32788 22764 32798 22820
rect 5864 22708 5874 22764
rect 5930 22708 5978 22764
rect 6034 22708 6082 22764
rect 6138 22708 6148 22764
rect 15188 22708 15198 22764
rect 15254 22708 15302 22764
rect 15358 22708 15406 22764
rect 15462 22708 15472 22764
rect 24512 22708 24522 22764
rect 24578 22708 24626 22764
rect 24682 22708 24730 22764
rect 24786 22708 24796 22764
rect 33836 22708 33846 22764
rect 33902 22708 33950 22764
rect 34006 22708 34054 22764
rect 34110 22708 34120 22764
rect 7970 22652 7980 22708
rect 8036 22652 14812 22708
rect 14868 22652 14878 22708
rect 26338 22652 26348 22708
rect 26404 22652 29148 22708
rect 29204 22652 29214 22708
rect 32498 22540 32508 22596
rect 32564 22540 33516 22596
rect 33572 22540 33582 22596
rect 18722 22428 18732 22484
rect 18788 22428 23548 22484
rect 23604 22428 23614 22484
rect 25554 22428 25564 22484
rect 25620 22428 26012 22484
rect 26068 22428 27580 22484
rect 27636 22428 27646 22484
rect 32162 22428 32172 22484
rect 32228 22428 33404 22484
rect 33460 22428 33470 22484
rect 11106 22316 11116 22372
rect 11172 22316 11900 22372
rect 11956 22316 11966 22372
rect 15474 22316 15484 22372
rect 15540 22316 16828 22372
rect 16884 22316 16894 22372
rect 23706 22316 23716 22372
rect 23772 22316 25676 22372
rect 25732 22316 25742 22372
rect 30482 22316 30492 22372
rect 30548 22316 31388 22372
rect 31444 22316 32396 22372
rect 32452 22316 32462 22372
rect 33730 22316 33740 22372
rect 33796 22316 34636 22372
rect 34692 22316 34702 22372
rect 23426 22204 23436 22260
rect 23492 22204 26012 22260
rect 26068 22204 30044 22260
rect 30100 22204 30110 22260
rect 33954 22204 33964 22260
rect 34020 22204 34318 22260
rect 34374 22204 34384 22260
rect 2034 22092 2044 22148
rect 2100 22092 5796 22148
rect 5852 22092 7364 22148
rect 7420 22092 8316 22148
rect 8372 22092 8382 22148
rect 30706 22092 30716 22148
rect 30772 22092 31052 22148
rect 31108 22092 32172 22148
rect 32228 22092 32238 22148
rect 30482 21980 30492 22036
rect 30548 21980 31836 22036
rect 31892 21980 32284 22036
rect 32340 21980 32350 22036
rect 10526 21924 10536 21980
rect 10592 21924 10640 21980
rect 10696 21924 10744 21980
rect 10800 21924 10810 21980
rect 19850 21924 19860 21980
rect 19916 21924 19964 21980
rect 20020 21924 20068 21980
rect 20124 21924 20134 21980
rect 29174 21924 29184 21980
rect 29240 21924 29288 21980
rect 29344 21924 29392 21980
rect 29448 21924 29458 21980
rect 38498 21924 38508 21980
rect 38564 21924 38612 21980
rect 38668 21924 38716 21980
rect 38772 21924 38782 21980
rect 14802 21868 14812 21924
rect 14868 21868 16604 21924
rect 16660 21868 16670 21924
rect 3154 21756 3164 21812
rect 3220 21756 5274 21812
rect 5330 21756 5340 21812
rect 10210 21756 10220 21812
rect 10276 21756 10892 21812
rect 10948 21756 10958 21812
rect 15092 21756 25340 21812
rect 25396 21756 25406 21812
rect 28700 21756 32732 21812
rect 32788 21756 32798 21812
rect 15092 21700 15148 21756
rect 28700 21700 28756 21756
rect 4050 21644 4060 21700
rect 4116 21644 6188 21700
rect 6244 21644 6524 21700
rect 6580 21644 6590 21700
rect 13794 21644 13804 21700
rect 13860 21644 14476 21700
rect 14532 21644 15148 21700
rect 21420 21644 25788 21700
rect 25844 21644 25854 21700
rect 26786 21644 26796 21700
rect 26852 21644 28700 21700
rect 28756 21644 28766 21700
rect 28914 21644 28924 21700
rect 28980 21644 32340 21700
rect 21420 21588 21476 21644
rect 32284 21588 32340 21644
rect 19394 21532 19404 21588
rect 19460 21532 19796 21588
rect 19852 21532 21476 21588
rect 21634 21532 21644 21588
rect 21700 21532 22652 21588
rect 22708 21532 23212 21588
rect 23268 21532 23278 21588
rect 27122 21532 27132 21588
rect 27188 21532 28588 21588
rect 28644 21532 29036 21588
rect 29092 21532 30156 21588
rect 30212 21532 30222 21588
rect 31322 21532 31332 21588
rect 31388 21532 31612 21588
rect 31668 21532 31678 21588
rect 32274 21532 32284 21588
rect 32340 21532 32620 21588
rect 32676 21532 32686 21588
rect 4722 21420 4732 21476
rect 4788 21420 5516 21476
rect 5572 21420 5582 21476
rect 8362 21420 8372 21476
rect 8428 21420 8876 21476
rect 8932 21420 8942 21476
rect 28074 21420 28084 21476
rect 28140 21420 31164 21476
rect 31220 21420 31230 21476
rect 21970 21308 21980 21364
rect 22036 21308 22316 21364
rect 22372 21308 22764 21364
rect 22820 21308 25228 21364
rect 25284 21308 25294 21364
rect 33506 21308 33516 21364
rect 33572 21308 34972 21364
rect 35028 21308 35038 21364
rect 30594 21196 30604 21252
rect 30660 21196 31164 21252
rect 31220 21196 31230 21252
rect 5864 21140 5874 21196
rect 5930 21140 5978 21196
rect 6034 21140 6082 21196
rect 6138 21140 6148 21196
rect 15188 21140 15198 21196
rect 15254 21140 15302 21196
rect 15358 21140 15406 21196
rect 15462 21140 15472 21196
rect 24512 21140 24522 21196
rect 24578 21140 24626 21196
rect 24682 21140 24730 21196
rect 24786 21140 24796 21196
rect 33836 21140 33846 21196
rect 33902 21140 33950 21196
rect 34006 21140 34054 21196
rect 34110 21140 34120 21196
rect 8372 21084 13692 21140
rect 13748 21084 13758 21140
rect 34850 21084 34860 21140
rect 34916 21084 35644 21140
rect 35700 21084 37660 21140
rect 37716 21084 37726 21140
rect 8372 21028 8428 21084
rect 5506 20972 5516 21028
rect 5572 20972 5582 21028
rect 6458 20972 6468 21028
rect 6524 20972 6860 21028
rect 6916 20972 7308 21028
rect 7364 20972 8428 21028
rect 11554 20972 11564 21028
rect 11620 20972 13562 21028
rect 13618 20972 13628 21028
rect 19394 20972 19404 21028
rect 19460 20972 21532 21028
rect 21588 20972 25788 21028
rect 25844 20972 25854 21028
rect 26450 20972 26460 21028
rect 26516 20972 26908 21028
rect 26964 20972 27468 21028
rect 27524 20972 27534 21028
rect 5516 20916 5572 20972
rect 25788 20916 25844 20972
rect 31276 20916 31332 21028
rect 31388 20972 31398 21028
rect 5516 20860 7700 20916
rect 12226 20860 12236 20916
rect 12292 20860 20188 20916
rect 20244 20860 20254 20916
rect 25788 20860 31332 20916
rect 36978 20860 36988 20916
rect 37044 20860 38892 20916
rect 38948 20860 38958 20916
rect 7644 20804 7700 20860
rect 37996 20804 38052 20860
rect 2034 20748 2044 20804
rect 2100 20748 2492 20804
rect 2548 20748 2558 20804
rect 5954 20748 5964 20804
rect 6020 20748 7420 20804
rect 7476 20748 7486 20804
rect 7644 20748 7812 20804
rect 7868 20748 13356 20804
rect 13412 20748 13422 20804
rect 13906 20748 13916 20804
rect 13972 20748 14700 20804
rect 14756 20748 14766 20804
rect 21746 20748 21756 20804
rect 21812 20748 26124 20804
rect 26180 20748 26190 20804
rect 33842 20748 33852 20804
rect 33908 20748 37156 20804
rect 37212 20748 37222 20804
rect 37986 20748 37996 20804
rect 38052 20748 38062 20804
rect 4050 20636 4060 20692
rect 4116 20636 7066 20692
rect 7122 20636 7132 20692
rect 20178 20636 20188 20692
rect 20244 20636 26236 20692
rect 26292 20636 26302 20692
rect 6626 20524 6636 20580
rect 6692 20524 7196 20580
rect 7252 20524 7980 20580
rect 8036 20524 8046 20580
rect 20290 20524 20300 20580
rect 20356 20524 21420 20580
rect 21476 20524 21486 20580
rect 24098 20524 24108 20580
rect 24164 20524 27076 20580
rect 27132 20524 27142 20580
rect 10526 20356 10536 20412
rect 10592 20356 10640 20412
rect 10696 20356 10744 20412
rect 10800 20356 10810 20412
rect 19850 20356 19860 20412
rect 19916 20356 19964 20412
rect 20020 20356 20068 20412
rect 20124 20356 20134 20412
rect 29174 20356 29184 20412
rect 29240 20356 29288 20412
rect 29344 20356 29392 20412
rect 29448 20356 29458 20412
rect 38498 20356 38508 20412
rect 38564 20356 38612 20412
rect 38668 20356 38716 20412
rect 38772 20356 38782 20412
rect 7410 20300 7420 20356
rect 7476 20300 8484 20356
rect 30930 20300 30940 20356
rect 30996 20300 32564 20356
rect 32620 20300 32630 20356
rect 34196 20300 34206 20356
rect 34262 20300 35980 20356
rect 36036 20300 36046 20356
rect 8428 20244 8484 20300
rect 8418 20188 8428 20244
rect 8484 20188 9436 20244
rect 9492 20188 9502 20244
rect 28802 20188 28812 20244
rect 28868 20188 31052 20244
rect 31108 20188 31118 20244
rect 32060 20188 35308 20244
rect 35364 20188 35374 20244
rect 9594 20076 9604 20132
rect 9660 20076 18956 20132
rect 19012 20076 19022 20132
rect 19898 20076 19908 20132
rect 19964 20076 23436 20132
rect 23492 20076 23502 20132
rect 23986 20076 23996 20132
rect 24052 20076 24556 20132
rect 24612 20076 24622 20132
rect 29036 20076 30268 20132
rect 30324 20076 30334 20132
rect 29036 20020 29092 20076
rect 2146 19964 2156 20020
rect 2212 19964 4172 20020
rect 4228 19964 4238 20020
rect 14354 19964 14364 20020
rect 14420 19964 20188 20020
rect 20244 19964 20254 20020
rect 22866 19964 22876 20020
rect 22932 19964 24444 20020
rect 24500 19964 29036 20020
rect 29092 19964 29102 20020
rect 29530 19964 29540 20020
rect 29596 19964 31276 20020
rect 31332 19964 31612 20020
rect 31668 19964 31678 20020
rect 32060 19908 32116 20188
rect 39200 20020 40000 20048
rect 38434 19964 38444 20020
rect 38500 19964 40000 20020
rect 39200 19936 40000 19964
rect 10658 19852 10668 19908
rect 10724 19852 12236 19908
rect 12292 19852 15596 19908
rect 15652 19852 15662 19908
rect 17948 19852 26908 19908
rect 17948 19796 18004 19852
rect 13906 19740 13916 19796
rect 13972 19740 15764 19796
rect 15820 19740 18004 19796
rect 21130 19740 21140 19796
rect 21196 19740 21756 19796
rect 21812 19740 21822 19796
rect 23426 19740 23436 19796
rect 23492 19740 23772 19796
rect 23828 19740 24108 19796
rect 24164 19740 24174 19796
rect 26852 19684 26908 19852
rect 29484 19852 29932 19908
rect 29988 19852 31388 19908
rect 31444 19852 31454 19908
rect 32050 19852 32060 19908
rect 32116 19852 32126 19908
rect 34626 19852 34636 19908
rect 34692 19852 35252 19908
rect 35308 19852 36428 19908
rect 36484 19852 36494 19908
rect 29484 19796 29540 19852
rect 29474 19740 29484 19796
rect 29540 19740 29550 19796
rect 29810 19740 29820 19796
rect 29876 19740 30604 19796
rect 30660 19740 30670 19796
rect 12562 19628 12572 19684
rect 12628 19628 14252 19684
rect 14308 19628 14318 19684
rect 26852 19628 31892 19684
rect 31948 19628 32340 19684
rect 32396 19628 32406 19684
rect 5864 19572 5874 19628
rect 5930 19572 5978 19628
rect 6034 19572 6082 19628
rect 6138 19572 6148 19628
rect 15188 19572 15198 19628
rect 15254 19572 15302 19628
rect 15358 19572 15406 19628
rect 15462 19572 15472 19628
rect 24512 19572 24522 19628
rect 24578 19572 24626 19628
rect 24682 19572 24730 19628
rect 24786 19572 24796 19628
rect 33836 19572 33846 19628
rect 33902 19572 33950 19628
rect 34006 19572 34054 19628
rect 34110 19572 34120 19628
rect 20514 19516 20524 19572
rect 20580 19516 22988 19572
rect 23044 19516 23054 19572
rect 23762 19516 23772 19572
rect 23828 19516 24332 19572
rect 24388 19516 24398 19572
rect 29250 19516 29260 19572
rect 29316 19516 29820 19572
rect 29876 19516 29886 19572
rect 30482 19516 30492 19572
rect 30548 19516 31164 19572
rect 31220 19516 31230 19572
rect 7970 19404 7980 19460
rect 8036 19404 10668 19460
rect 10724 19404 10734 19460
rect 13402 19404 13412 19460
rect 13468 19404 13916 19460
rect 13972 19404 13982 19460
rect 20290 19404 20300 19460
rect 20356 19404 21812 19460
rect 21868 19404 21878 19460
rect 22418 19404 22428 19460
rect 22484 19404 25284 19460
rect 25340 19404 25350 19460
rect 36418 19404 36428 19460
rect 36484 19404 37156 19460
rect 37212 19404 38332 19460
rect 38388 19404 38398 19460
rect 11890 19292 11900 19348
rect 11956 19292 12460 19348
rect 12516 19292 14028 19348
rect 14084 19292 14094 19348
rect 14242 19292 14252 19348
rect 14308 19292 17164 19348
rect 17220 19292 18172 19348
rect 18228 19292 18238 19348
rect 4610 19180 4620 19236
rect 4676 19180 5516 19236
rect 5572 19180 5582 19236
rect 7970 19180 7980 19236
rect 8036 19180 8428 19236
rect 13682 19180 13692 19236
rect 13748 19180 14476 19236
rect 14532 19180 17500 19236
rect 17556 19180 17780 19236
rect 17836 19180 17846 19236
rect 19506 19180 19516 19236
rect 19572 19180 19582 19236
rect 22978 19180 22988 19236
rect 23044 19180 23996 19236
rect 24052 19180 24062 19236
rect 25442 19180 25452 19236
rect 25508 19180 26572 19236
rect 26628 19180 26638 19236
rect 29138 19180 29148 19236
rect 29204 19180 30548 19236
rect 30604 19180 30614 19236
rect 31042 19180 31052 19236
rect 31108 19180 31892 19236
rect 37594 19180 37604 19236
rect 37660 19180 38332 19236
rect 38388 19180 38398 19236
rect 8372 19012 8428 19180
rect 19516 19124 19572 19180
rect 31836 19124 31892 19180
rect 13570 19068 13580 19124
rect 13636 19068 14028 19124
rect 14084 19068 14094 19124
rect 19516 19068 19740 19124
rect 19796 19068 19964 19124
rect 20020 19068 25900 19124
rect 25956 19068 25966 19124
rect 31826 19068 31836 19124
rect 31892 19068 31902 19124
rect 8372 18956 9044 19012
rect 9100 18956 11284 19012
rect 11340 18956 11350 19012
rect 15092 18956 23100 19012
rect 23156 18956 23166 19012
rect 4162 18844 4172 18900
rect 4228 18844 5740 18900
rect 5796 18844 7812 18900
rect 7868 18844 7878 18900
rect 10526 18788 10536 18844
rect 10592 18788 10640 18844
rect 10696 18788 10744 18844
rect 10800 18788 10810 18844
rect 15092 18788 15148 18956
rect 20626 18844 20636 18900
rect 20692 18844 29036 18900
rect 29092 18844 29102 18900
rect 19850 18788 19860 18844
rect 19916 18788 19964 18844
rect 20020 18788 20068 18844
rect 20124 18788 20134 18844
rect 29174 18788 29184 18844
rect 29240 18788 29288 18844
rect 29344 18788 29392 18844
rect 29448 18788 29458 18844
rect 38498 18788 38508 18844
rect 38564 18788 38612 18844
rect 38668 18788 38716 18844
rect 38772 18788 38782 18844
rect 13794 18732 13804 18788
rect 13860 18732 14364 18788
rect 14420 18732 14924 18788
rect 14980 18732 15148 18788
rect 30258 18732 30268 18788
rect 30324 18732 31164 18788
rect 31220 18732 31230 18788
rect 18834 18620 18844 18676
rect 18900 18620 18910 18676
rect 19058 18620 19068 18676
rect 19124 18620 19404 18676
rect 19460 18620 19470 18676
rect 23548 18620 25004 18676
rect 25060 18620 25564 18676
rect 25620 18620 25630 18676
rect 18844 18452 18900 18620
rect 23548 18564 23604 18620
rect 21308 18508 22092 18564
rect 22148 18508 22158 18564
rect 22754 18508 22764 18564
rect 22820 18508 23380 18564
rect 23436 18508 23604 18564
rect 23762 18508 23772 18564
rect 23828 18508 24108 18564
rect 24164 18508 24174 18564
rect 29474 18508 29484 18564
rect 29540 18508 30268 18564
rect 30324 18508 30334 18564
rect 21308 18452 21364 18508
rect 8194 18396 8204 18452
rect 8260 18396 9436 18452
rect 9492 18396 9502 18452
rect 9650 18396 9660 18452
rect 9716 18396 10892 18452
rect 10948 18396 11116 18452
rect 11172 18396 12908 18452
rect 12964 18396 13244 18452
rect 13300 18396 13310 18452
rect 13402 18396 13412 18452
rect 13468 18396 13804 18452
rect 13860 18396 13870 18452
rect 14130 18396 14140 18452
rect 14196 18396 15148 18452
rect 18844 18396 20300 18452
rect 20356 18396 20366 18452
rect 20748 18396 21364 18452
rect 21522 18396 21532 18452
rect 21588 18396 22540 18452
rect 22596 18396 22606 18452
rect 24602 18396 24612 18452
rect 24668 18396 28028 18452
rect 28084 18396 29820 18452
rect 29876 18396 29886 18452
rect 34458 18396 34468 18452
rect 34524 18396 34748 18452
rect 34804 18396 34814 18452
rect 15092 18340 15148 18396
rect 20748 18340 20804 18396
rect 15092 18284 19180 18340
rect 19236 18284 19246 18340
rect 20178 18284 20188 18340
rect 20244 18284 20748 18340
rect 20804 18284 20814 18340
rect 25218 18284 25228 18340
rect 25284 18284 25788 18340
rect 25844 18284 26908 18340
rect 26964 18284 27692 18340
rect 27748 18284 27758 18340
rect 26460 18228 26516 18284
rect 20514 18172 20524 18228
rect 20580 18172 21084 18228
rect 21140 18172 22316 18228
rect 22372 18172 22382 18228
rect 24770 18172 24780 18228
rect 24836 18172 25564 18228
rect 25620 18172 25630 18228
rect 26450 18172 26460 18228
rect 26516 18172 26526 18228
rect 29362 18172 29372 18228
rect 29428 18172 30268 18228
rect 30324 18172 31164 18228
rect 31220 18172 31230 18228
rect 34402 18172 34412 18228
rect 34468 18172 35084 18228
rect 35140 18172 35150 18228
rect 8530 18060 8540 18116
rect 8596 18060 8988 18116
rect 9044 18060 9054 18116
rect 20402 18060 20412 18116
rect 20468 18060 21868 18116
rect 21924 18060 21934 18116
rect 22866 18060 22876 18116
rect 22932 18060 24332 18116
rect 24388 18060 24398 18116
rect 5864 18004 5874 18060
rect 5930 18004 5978 18060
rect 6034 18004 6082 18060
rect 6138 18004 6148 18060
rect 15188 18004 15198 18060
rect 15254 18004 15302 18060
rect 15358 18004 15406 18060
rect 15462 18004 15472 18060
rect 8530 17836 8540 17892
rect 8596 17836 8764 17892
rect 8820 17836 8830 17892
rect 9874 17836 9884 17892
rect 9940 17836 10724 17892
rect 10780 17836 10790 17892
rect 15092 17836 18172 17892
rect 18228 17836 18238 17892
rect 15092 17780 15148 17836
rect 11890 17724 11900 17780
rect 11956 17724 12684 17780
rect 12740 17724 15148 17780
rect 24108 17780 24164 18060
rect 24512 18004 24522 18060
rect 24578 18004 24626 18060
rect 24682 18004 24730 18060
rect 24786 18004 24796 18060
rect 33836 18004 33846 18060
rect 33902 18004 33950 18060
rect 34006 18004 34054 18060
rect 34110 18004 34120 18060
rect 24322 17836 24332 17892
rect 24388 17836 26684 17892
rect 26740 17836 27076 17892
rect 27132 17836 27142 17892
rect 24108 17724 26012 17780
rect 26068 17724 26572 17780
rect 26628 17724 26638 17780
rect 26852 17724 27188 17780
rect 27244 17724 27254 17780
rect 28634 17724 28644 17780
rect 28700 17724 29372 17780
rect 29428 17724 29596 17780
rect 29652 17724 31108 17780
rect 31164 17724 32060 17780
rect 32116 17724 32126 17780
rect 26852 17668 26908 17724
rect 18162 17612 18172 17668
rect 18228 17612 25172 17668
rect 25228 17612 25238 17668
rect 25442 17612 25452 17668
rect 25508 17612 26908 17668
rect 29810 17612 29820 17668
rect 29876 17612 29886 17668
rect 29820 17556 29876 17612
rect 19282 17500 19292 17556
rect 19348 17500 20020 17556
rect 20076 17500 21756 17556
rect 21812 17500 21822 17556
rect 22642 17500 22652 17556
rect 22708 17500 23660 17556
rect 23716 17500 24220 17556
rect 24276 17500 24286 17556
rect 26674 17500 26684 17556
rect 26740 17500 28140 17556
rect 28196 17500 29876 17556
rect 20402 17388 20412 17444
rect 20468 17388 21532 17444
rect 21588 17388 21598 17444
rect 25890 17388 25900 17444
rect 25956 17388 30098 17444
rect 30154 17388 30164 17444
rect 20290 17276 20300 17332
rect 20356 17276 22316 17332
rect 22372 17276 22382 17332
rect 34178 17276 34188 17332
rect 34244 17276 35084 17332
rect 35140 17276 35150 17332
rect 10526 17220 10536 17276
rect 10592 17220 10640 17276
rect 10696 17220 10744 17276
rect 10800 17220 10810 17276
rect 19850 17220 19860 17276
rect 19916 17220 19964 17276
rect 20020 17220 20068 17276
rect 20124 17220 20134 17276
rect 29174 17220 29184 17276
rect 29240 17220 29288 17276
rect 29344 17220 29392 17276
rect 29448 17220 29458 17276
rect 38498 17220 38508 17276
rect 38564 17220 38612 17276
rect 38668 17220 38716 17276
rect 38772 17220 38782 17276
rect 13356 17164 14476 17220
rect 14532 17164 15596 17220
rect 15652 17164 15662 17220
rect 25442 17164 25452 17220
rect 25508 17164 25732 17220
rect 25788 17164 26684 17220
rect 26740 17164 26750 17220
rect 27794 17164 27804 17220
rect 27860 17164 29036 17220
rect 29092 17164 29102 17220
rect 32396 17164 37996 17220
rect 38052 17164 38062 17220
rect 13356 17108 13412 17164
rect 32396 17108 32452 17164
rect 39200 17108 40000 17136
rect 8978 17052 8988 17108
rect 9044 17052 9716 17108
rect 9772 17052 13412 17108
rect 13570 17052 13580 17108
rect 13636 17052 13860 17108
rect 13916 17052 13926 17108
rect 18386 17052 18396 17108
rect 18452 17052 20524 17108
rect 20580 17052 20972 17108
rect 21028 17052 21038 17108
rect 21746 17052 21756 17108
rect 21812 17052 23044 17108
rect 23100 17052 23772 17108
rect 23828 17052 32452 17108
rect 37594 17052 37604 17108
rect 37660 17052 38332 17108
rect 38388 17052 40000 17108
rect 39200 17024 40000 17052
rect 12114 16940 12124 16996
rect 12180 16940 13020 16996
rect 13076 16940 16380 16996
rect 16436 16940 17724 16996
rect 17780 16940 17790 16996
rect 19394 16940 19404 16996
rect 19460 16940 23660 16996
rect 23716 16940 23726 16996
rect 24322 16940 24332 16996
rect 24388 16940 25564 16996
rect 25620 16940 25630 16996
rect 25722 16940 25732 16996
rect 25788 16940 27804 16996
rect 27860 16940 27870 16996
rect 30482 16940 30492 16996
rect 30548 16940 31108 16996
rect 31164 16940 31556 16996
rect 19618 16828 19628 16884
rect 19684 16828 20524 16884
rect 20580 16828 20590 16884
rect 20748 16772 20804 16940
rect 21242 16828 21252 16884
rect 21308 16828 26012 16884
rect 26068 16828 26078 16884
rect 26282 16828 26292 16884
rect 26348 16828 28588 16884
rect 28644 16828 28654 16884
rect 29362 16828 29372 16884
rect 29428 16828 30380 16884
rect 30436 16828 30446 16884
rect 20738 16716 20748 16772
rect 20804 16716 20814 16772
rect 21858 16716 21868 16772
rect 21924 16716 22764 16772
rect 22820 16716 22830 16772
rect 31500 16660 31556 16940
rect 31714 16828 31724 16884
rect 31780 16828 32172 16884
rect 32228 16828 32844 16884
rect 32900 16828 32910 16884
rect 34066 16716 34076 16772
rect 34132 16716 35308 16772
rect 35364 16716 35374 16772
rect 36978 16716 36988 16772
rect 37044 16716 37212 16772
rect 37268 16716 37278 16772
rect 18050 16604 18060 16660
rect 18116 16604 18788 16660
rect 18844 16604 21980 16660
rect 22036 16604 22046 16660
rect 22212 16604 22222 16660
rect 22278 16604 30156 16660
rect 30212 16604 30222 16660
rect 31500 16604 31724 16660
rect 31780 16604 31790 16660
rect 31994 16604 32004 16660
rect 32060 16604 37324 16660
rect 37380 16604 37390 16660
rect 20850 16492 20860 16548
rect 20916 16492 21756 16548
rect 21812 16492 21822 16548
rect 28578 16492 28588 16548
rect 28644 16492 29820 16548
rect 29876 16492 30716 16548
rect 30772 16492 30782 16548
rect 5864 16436 5874 16492
rect 5930 16436 5978 16492
rect 6034 16436 6082 16492
rect 6138 16436 6148 16492
rect 15188 16436 15198 16492
rect 15254 16436 15302 16492
rect 15358 16436 15406 16492
rect 15462 16436 15472 16492
rect 24512 16436 24522 16492
rect 24578 16436 24626 16492
rect 24682 16436 24730 16492
rect 24786 16436 24796 16492
rect 33836 16436 33846 16492
rect 33902 16436 33950 16492
rect 34006 16436 34054 16492
rect 34110 16436 34120 16492
rect 16706 16380 16716 16436
rect 16772 16380 17276 16436
rect 17332 16380 22484 16436
rect 22540 16380 22550 16436
rect 27402 16380 27412 16436
rect 27468 16380 28252 16436
rect 28308 16380 30828 16436
rect 30884 16380 32004 16436
rect 32060 16380 32070 16436
rect 8642 16268 8652 16324
rect 8708 16268 33516 16324
rect 33572 16268 33582 16324
rect 34402 16268 34412 16324
rect 34468 16268 37380 16324
rect 37436 16268 37446 16324
rect 18834 16156 18844 16212
rect 18900 16156 21868 16212
rect 21924 16156 21934 16212
rect 28354 16156 28364 16212
rect 28420 16156 29932 16212
rect 29988 16156 29998 16212
rect 30370 16156 30380 16212
rect 30436 16156 31388 16212
rect 31444 16156 31454 16212
rect 36474 16156 36484 16212
rect 36540 16156 36876 16212
rect 36932 16156 36942 16212
rect 10322 16044 10332 16100
rect 10388 16044 10892 16100
rect 10948 16044 11340 16100
rect 11396 16044 11406 16100
rect 19954 16044 19964 16100
rect 20020 16044 21308 16100
rect 21364 16044 21756 16100
rect 21812 16044 23100 16100
rect 23156 16044 23166 16100
rect 23930 16044 23940 16100
rect 23996 16044 24575 16100
rect 24631 16044 24641 16100
rect 25414 16044 25452 16100
rect 25508 16044 25518 16100
rect 29026 16044 29036 16100
rect 29092 16044 30994 16100
rect 31050 16044 31060 16100
rect 36306 16044 36316 16100
rect 36372 16044 37100 16100
rect 37156 16044 37166 16100
rect 22306 15932 22316 15988
rect 22372 15932 22876 15988
rect 22932 15932 22942 15988
rect 19618 15820 19628 15876
rect 19684 15820 20524 15876
rect 20580 15820 21476 15876
rect 21532 15820 21542 15876
rect 21970 15820 21980 15876
rect 22036 15820 22204 15876
rect 22260 15820 23492 15876
rect 23548 15820 23558 15876
rect 33170 15820 33180 15876
rect 33236 15820 33852 15876
rect 33908 15820 35980 15876
rect 36036 15820 36046 15876
rect 10526 15652 10536 15708
rect 10592 15652 10640 15708
rect 10696 15652 10744 15708
rect 10800 15652 10810 15708
rect 19850 15652 19860 15708
rect 19916 15652 19964 15708
rect 20020 15652 20068 15708
rect 20124 15652 20134 15708
rect 29174 15652 29184 15708
rect 29240 15652 29288 15708
rect 29344 15652 29392 15708
rect 29448 15652 29458 15708
rect 38498 15652 38508 15708
rect 38564 15652 38612 15708
rect 38668 15652 38716 15708
rect 38772 15652 38782 15708
rect 20794 15484 20804 15540
rect 20860 15484 21122 15540
rect 21178 15484 21188 15540
rect 31378 15484 31388 15540
rect 31444 15484 31836 15540
rect 31892 15484 31902 15540
rect 31490 15372 31500 15428
rect 31556 15372 31724 15428
rect 31780 15372 31790 15428
rect 36194 15372 36204 15428
rect 36260 15372 36876 15428
rect 36932 15372 36942 15428
rect 12450 15260 12460 15316
rect 12516 15260 13468 15316
rect 13524 15260 14252 15316
rect 14308 15260 14318 15316
rect 18050 15260 18060 15316
rect 18116 15260 19292 15316
rect 19348 15260 19358 15316
rect 20738 15260 20748 15316
rect 20804 15260 21644 15316
rect 21700 15260 21710 15316
rect 22418 15260 22428 15316
rect 22484 15260 23436 15316
rect 23492 15260 24388 15316
rect 24444 15260 24454 15316
rect 28130 15260 28140 15316
rect 28196 15260 28588 15316
rect 28644 15260 28654 15316
rect 35522 15260 35532 15316
rect 35588 15260 36988 15316
rect 37044 15260 37054 15316
rect 33842 15148 33852 15204
rect 33908 15148 35308 15204
rect 35364 15148 35374 15204
rect 36204 15092 36260 15260
rect 20402 15036 20412 15092
rect 20468 15036 21308 15092
rect 21364 15036 21644 15092
rect 21700 15036 21710 15092
rect 32946 15036 32956 15092
rect 33012 15036 33628 15092
rect 33684 15036 33694 15092
rect 34010 15036 34020 15092
rect 34076 15036 34300 15092
rect 34356 15036 34366 15092
rect 36194 15036 36204 15092
rect 36260 15036 36270 15092
rect 21132 14924 21142 14980
rect 21198 14924 22764 14980
rect 22820 14924 22830 14980
rect 5864 14868 5874 14924
rect 5930 14868 5978 14924
rect 6034 14868 6082 14924
rect 6138 14868 6148 14924
rect 15188 14868 15198 14924
rect 15254 14868 15302 14924
rect 15358 14868 15406 14924
rect 15462 14868 15472 14924
rect 24512 14868 24522 14924
rect 24578 14868 24626 14924
rect 24682 14868 24730 14924
rect 24786 14868 24796 14924
rect 33836 14868 33846 14924
rect 33902 14868 33950 14924
rect 34006 14868 34054 14924
rect 34110 14868 34120 14924
rect 10210 14700 10220 14756
rect 10276 14700 13580 14756
rect 13636 14700 13646 14756
rect 22194 14700 22204 14756
rect 22260 14700 38052 14756
rect 25890 14588 25900 14644
rect 25956 14588 27076 14644
rect 27132 14588 29316 14644
rect 29372 14588 29382 14644
rect 16930 14476 16940 14532
rect 16996 14476 19404 14532
rect 19460 14476 19470 14532
rect 20066 14476 20076 14532
rect 20132 14476 21308 14532
rect 21364 14476 22652 14532
rect 22708 14476 22718 14532
rect 25330 14476 25340 14532
rect 25396 14476 26404 14532
rect 26460 14476 26470 14532
rect 37996 14420 38052 14700
rect 21970 14364 21980 14420
rect 22036 14364 23100 14420
rect 23156 14364 23166 14420
rect 24826 14364 24836 14420
rect 24892 14364 25788 14420
rect 25844 14364 25854 14420
rect 33842 14364 33852 14420
rect 33908 14364 34300 14420
rect 34356 14364 34366 14420
rect 37986 14364 37996 14420
rect 38052 14364 38062 14420
rect 13906 14252 13916 14308
rect 13972 14252 14308 14308
rect 14364 14252 14374 14308
rect 37594 14252 37604 14308
rect 37660 14252 38332 14308
rect 38388 14252 38948 14308
rect 38892 14196 38948 14252
rect 39200 14196 40000 14224
rect 14466 14140 14476 14196
rect 14532 14140 14700 14196
rect 14756 14140 14766 14196
rect 26852 14140 27244 14196
rect 27300 14140 28812 14196
rect 28868 14140 28878 14196
rect 35578 14140 35588 14196
rect 35644 14140 36298 14196
rect 36354 14140 36364 14196
rect 38892 14140 40000 14196
rect 10526 14084 10536 14140
rect 10592 14084 10640 14140
rect 10696 14084 10744 14140
rect 10800 14084 10810 14140
rect 19850 14084 19860 14140
rect 19916 14084 19964 14140
rect 20020 14084 20068 14140
rect 20124 14084 20134 14140
rect 26852 14084 26908 14140
rect 29174 14084 29184 14140
rect 29240 14084 29288 14140
rect 29344 14084 29392 14140
rect 29448 14084 29458 14140
rect 38498 14084 38508 14140
rect 38564 14084 38612 14140
rect 38668 14084 38716 14140
rect 38772 14084 38782 14140
rect 39200 14112 40000 14140
rect 20850 14028 20860 14084
rect 20916 14028 21308 14084
rect 21364 14028 23548 14084
rect 23604 14028 26908 14084
rect 34514 14028 34524 14084
rect 34580 14028 35308 14084
rect 35364 14028 35812 14084
rect 19394 13916 19404 13972
rect 19460 13916 22876 13972
rect 22932 13916 22942 13972
rect 23930 13916 23940 13972
rect 23996 13916 29708 13972
rect 29764 13916 29774 13972
rect 34402 13916 34412 13972
rect 34468 13916 34478 13972
rect 13570 13804 13580 13860
rect 13636 13804 14924 13860
rect 14980 13804 14990 13860
rect 15698 13804 15708 13860
rect 15764 13804 26908 13860
rect 23220 13692 23230 13748
rect 23286 13692 23772 13748
rect 23828 13692 23838 13748
rect 26852 13636 26908 13804
rect 31574 13692 31612 13748
rect 31668 13692 31678 13748
rect 33058 13692 33068 13748
rect 33124 13692 33628 13748
rect 33684 13692 33694 13748
rect 26852 13580 30660 13636
rect 30716 13580 31388 13636
rect 31444 13580 33628 13636
rect 33684 13580 33694 13636
rect 9212 13468 10332 13524
rect 10388 13468 10398 13524
rect 21634 13468 21644 13524
rect 21700 13468 22876 13524
rect 22932 13468 22942 13524
rect 24322 13468 24332 13524
rect 24388 13468 25340 13524
rect 25396 13468 25406 13524
rect 29922 13468 29932 13524
rect 29988 13468 30996 13524
rect 31052 13468 31062 13524
rect 31154 13468 31164 13524
rect 31220 13468 31612 13524
rect 31668 13468 31678 13524
rect 5864 13300 5874 13356
rect 5930 13300 5978 13356
rect 6034 13300 6082 13356
rect 6138 13300 6148 13356
rect 9212 13300 9268 13468
rect 34412 13412 34468 13916
rect 35756 13748 35812 14028
rect 35746 13692 35756 13748
rect 35812 13692 35822 13748
rect 36362 13468 36372 13524
rect 36428 13468 37436 13524
rect 37492 13468 37502 13524
rect 13682 13356 13692 13412
rect 13748 13356 14140 13412
rect 14196 13356 14532 13412
rect 14588 13356 15036 13412
rect 15092 13356 15102 13412
rect 17266 13356 17276 13412
rect 17332 13356 18172 13412
rect 18228 13356 18238 13412
rect 21522 13356 21532 13412
rect 21588 13356 21598 13412
rect 21970 13356 21980 13412
rect 22036 13356 22316 13412
rect 22372 13356 22988 13412
rect 23044 13356 23054 13412
rect 30146 13356 30156 13412
rect 30212 13356 31500 13412
rect 31556 13356 31566 13412
rect 34290 13356 34300 13412
rect 34356 13356 34468 13412
rect 35410 13356 35420 13412
rect 35476 13356 36988 13412
rect 37044 13356 37054 13412
rect 37202 13356 37212 13412
rect 37268 13356 37278 13412
rect 15188 13300 15198 13356
rect 15254 13300 15302 13356
rect 15358 13300 15406 13356
rect 15462 13300 15472 13356
rect 21532 13300 21588 13356
rect 24512 13300 24522 13356
rect 24578 13300 24626 13356
rect 24682 13300 24730 13356
rect 24786 13300 24796 13356
rect 33836 13300 33846 13356
rect 33902 13300 33950 13356
rect 34006 13300 34054 13356
rect 34110 13300 34120 13356
rect 37212 13300 37268 13356
rect 9202 13244 9212 13300
rect 9268 13244 9278 13300
rect 21532 13244 23212 13300
rect 23268 13244 23278 13300
rect 24882 13244 24892 13300
rect 24948 13244 24958 13300
rect 31266 13244 31276 13300
rect 31332 13244 32060 13300
rect 32116 13244 32126 13300
rect 34636 13244 36876 13300
rect 36932 13244 37268 13300
rect 24892 13188 24948 13244
rect 34636 13188 34692 13244
rect 13626 13132 13636 13188
rect 13692 13132 14028 13188
rect 14084 13132 14094 13188
rect 23090 13132 23100 13188
rect 23156 13132 23324 13188
rect 23380 13132 24108 13188
rect 24164 13132 34468 13188
rect 34626 13132 34636 13188
rect 34692 13132 34702 13188
rect 34412 13076 34468 13132
rect 13906 13020 13916 13076
rect 13972 13020 14196 13076
rect 14252 13020 27804 13076
rect 27860 13020 27870 13076
rect 31938 13020 31948 13076
rect 32004 13020 33180 13076
rect 33236 13020 34356 13076
rect 34412 13020 38108 13076
rect 38164 13020 38174 13076
rect 10994 12908 11004 12964
rect 11060 12908 11452 12964
rect 11508 12908 11518 12964
rect 10210 12796 10220 12852
rect 10276 12796 13804 12852
rect 13860 12796 13870 12852
rect 14588 12740 14644 13020
rect 34300 12964 34356 13020
rect 17714 12908 17724 12964
rect 17780 12908 20188 12964
rect 20244 12908 20254 12964
rect 20514 12908 20524 12964
rect 20580 12908 21308 12964
rect 21364 12908 23100 12964
rect 23156 12908 23166 12964
rect 29586 12908 29596 12964
rect 29652 12908 30828 12964
rect 30884 12908 30894 12964
rect 32722 12908 32732 12964
rect 32788 12908 33852 12964
rect 33908 12908 33918 12964
rect 34300 12908 34636 12964
rect 34692 12908 34702 12964
rect 35540 12908 35550 12964
rect 35606 12908 37156 12964
rect 37212 12908 37222 12964
rect 15026 12796 15036 12852
rect 15092 12796 17276 12852
rect 17332 12796 18340 12852
rect 18396 12796 18406 12852
rect 20402 12796 20412 12852
rect 20468 12796 22184 12852
rect 22240 12796 22764 12852
rect 22820 12796 23436 12852
rect 23492 12796 23502 12852
rect 34084 12796 34094 12852
rect 34150 12796 34300 12852
rect 34356 12796 34366 12852
rect 35420 12796 35868 12852
rect 35924 12796 35934 12852
rect 36082 12796 36092 12852
rect 36148 12796 37902 12852
rect 37958 12796 37968 12852
rect 35420 12740 35476 12796
rect 9538 12684 9548 12740
rect 9604 12684 10668 12740
rect 10724 12684 11900 12740
rect 11956 12684 11966 12740
rect 14578 12684 14588 12740
rect 14644 12684 14654 12740
rect 31574 12684 31612 12740
rect 31668 12684 31678 12740
rect 33618 12684 33628 12740
rect 33684 12684 33908 12740
rect 33964 12684 34636 12740
rect 34692 12684 35252 12740
rect 35308 12684 35476 12740
rect 35634 12684 35644 12740
rect 35700 12684 36540 12740
rect 36596 12684 37660 12740
rect 37716 12684 37726 12740
rect 10526 12516 10536 12572
rect 10592 12516 10640 12572
rect 10696 12516 10744 12572
rect 10800 12516 10810 12572
rect 19850 12516 19860 12572
rect 19916 12516 19964 12572
rect 20020 12516 20068 12572
rect 20124 12516 20134 12572
rect 29174 12516 29184 12572
rect 29240 12516 29288 12572
rect 29344 12516 29392 12572
rect 29448 12516 29458 12572
rect 38498 12516 38508 12572
rect 38564 12516 38612 12572
rect 38668 12516 38716 12572
rect 38772 12516 38782 12572
rect 7298 12348 7308 12404
rect 7364 12348 8652 12404
rect 8708 12348 9884 12404
rect 9940 12348 9950 12404
rect 10994 12348 11004 12404
rect 11060 12348 13636 12404
rect 13692 12348 13702 12404
rect 14690 12348 14700 12404
rect 14756 12348 30492 12404
rect 30548 12348 30558 12404
rect 7634 12236 7644 12292
rect 7700 12236 9940 12292
rect 10098 12236 10108 12292
rect 10164 12236 10668 12292
rect 10724 12236 10892 12292
rect 10948 12236 14364 12292
rect 14420 12236 14430 12292
rect 28578 12236 28588 12292
rect 28644 12236 32620 12292
rect 32676 12236 32686 12292
rect 9884 12180 9940 12236
rect 8026 12124 8036 12180
rect 8092 12124 9604 12180
rect 9660 12124 9670 12180
rect 9884 12124 11004 12180
rect 11060 12124 11070 12180
rect 12058 12124 12068 12180
rect 12124 12124 14084 12180
rect 14140 12124 14150 12180
rect 18050 12124 18060 12180
rect 18116 12124 19628 12180
rect 19684 12124 19694 12180
rect 20178 12124 20188 12180
rect 20244 12124 25116 12180
rect 25172 12124 25182 12180
rect 31826 12124 31836 12180
rect 31892 12124 32732 12180
rect 32788 12124 32798 12180
rect 7858 12012 7868 12068
rect 7924 12012 13132 12068
rect 13188 12012 13198 12068
rect 14130 11788 14140 11844
rect 14196 11788 14700 11844
rect 14756 11788 14766 11844
rect 21074 11788 21084 11844
rect 21140 11788 23212 11844
rect 23268 11788 23278 11844
rect 5864 11732 5874 11788
rect 5930 11732 5978 11788
rect 6034 11732 6082 11788
rect 6138 11732 6148 11788
rect 15188 11732 15198 11788
rect 15254 11732 15302 11788
rect 15358 11732 15406 11788
rect 15462 11732 15472 11788
rect 24512 11732 24522 11788
rect 24578 11732 24626 11788
rect 24682 11732 24730 11788
rect 24786 11732 24796 11788
rect 33836 11732 33846 11788
rect 33902 11732 33950 11788
rect 34006 11732 34054 11788
rect 34110 11732 34120 11788
rect 7074 11676 7084 11732
rect 7140 11676 7150 11732
rect 25106 11676 25116 11732
rect 25172 11676 28700 11732
rect 28756 11676 29372 11732
rect 29428 11676 29438 11732
rect 7084 11620 7140 11676
rect 5842 11564 5852 11620
rect 5908 11564 10668 11620
rect 10724 11564 12236 11620
rect 12292 11564 12302 11620
rect 12562 11452 12572 11508
rect 12628 11452 14588 11508
rect 14644 11452 14654 11508
rect 17042 11452 17052 11508
rect 17108 11452 17668 11508
rect 17724 11452 17734 11508
rect 21970 11452 21980 11508
rect 22036 11452 28084 11508
rect 28140 11452 28588 11508
rect 28644 11452 28654 11508
rect 8772 11340 8782 11396
rect 8838 11340 9324 11396
rect 9380 11340 9390 11396
rect 10378 11340 10388 11396
rect 10444 11340 12068 11396
rect 12124 11340 12134 11396
rect 12804 11340 12814 11396
rect 12870 11340 14028 11396
rect 14084 11340 14094 11396
rect 18722 11340 18732 11396
rect 18788 11340 20524 11396
rect 20580 11340 20590 11396
rect 39200 11284 40000 11312
rect 7970 11228 7980 11284
rect 8036 11228 9044 11284
rect 9100 11228 9110 11284
rect 13738 11228 13748 11284
rect 13804 11228 14364 11284
rect 14420 11228 14430 11284
rect 37594 11228 37604 11284
rect 37660 11228 38332 11284
rect 38388 11228 40000 11284
rect 39200 11200 40000 11228
rect 25890 11116 25900 11172
rect 25956 11116 26908 11172
rect 26964 11116 26974 11172
rect 30482 11116 30492 11172
rect 30548 11116 31164 11172
rect 31220 11116 31230 11172
rect 10526 10948 10536 11004
rect 10592 10948 10640 11004
rect 10696 10948 10744 11004
rect 10800 10948 10810 11004
rect 19850 10948 19860 11004
rect 19916 10948 19964 11004
rect 20020 10948 20068 11004
rect 20124 10948 20134 11004
rect 29174 10948 29184 11004
rect 29240 10948 29288 11004
rect 29344 10948 29392 11004
rect 29448 10948 29458 11004
rect 38498 10948 38508 11004
rect 38564 10948 38612 11004
rect 38668 10948 38716 11004
rect 38772 10948 38782 11004
rect 10098 10780 10108 10836
rect 10164 10780 10174 10836
rect 20514 10780 20524 10836
rect 20580 10780 21028 10836
rect 21084 10780 21094 10836
rect 26002 10780 26012 10836
rect 26068 10780 26348 10836
rect 26404 10780 26414 10836
rect 37258 10780 37268 10836
rect 37324 10780 38220 10836
rect 38276 10780 38286 10836
rect 8306 10668 8316 10724
rect 8372 10668 9436 10724
rect 9492 10668 9502 10724
rect 10108 10612 10164 10780
rect 36642 10668 36652 10724
rect 36708 10668 37660 10724
rect 37716 10668 37726 10724
rect 8642 10556 8652 10612
rect 8708 10556 10164 10612
rect 13458 10556 13468 10612
rect 13524 10556 19292 10612
rect 19348 10556 19740 10612
rect 19796 10556 19806 10612
rect 9874 10444 9884 10500
rect 9940 10444 10220 10500
rect 10276 10444 10286 10500
rect 29250 10332 29260 10388
rect 29316 10332 29708 10388
rect 29764 10332 30604 10388
rect 30660 10332 30670 10388
rect 8418 10220 8428 10276
rect 8484 10220 10164 10276
rect 10220 10220 12572 10276
rect 12628 10220 12638 10276
rect 5864 10164 5874 10220
rect 5930 10164 5978 10220
rect 6034 10164 6082 10220
rect 6138 10164 6148 10220
rect 15188 10164 15198 10220
rect 15254 10164 15302 10220
rect 15358 10164 15406 10220
rect 15462 10164 15472 10220
rect 24512 10164 24522 10220
rect 24578 10164 24626 10220
rect 24682 10164 24730 10220
rect 24786 10164 24796 10220
rect 33836 10164 33846 10220
rect 33902 10164 33950 10220
rect 34006 10164 34054 10220
rect 34110 10164 34120 10220
rect 11218 10108 11228 10164
rect 11284 10108 12964 10164
rect 13020 10108 13030 10164
rect 23874 10108 23884 10164
rect 23940 10108 23950 10164
rect 26002 10108 26012 10164
rect 26068 10108 29036 10164
rect 29092 10108 29932 10164
rect 29988 10108 29998 10164
rect 23884 10052 23940 10108
rect 10452 9996 10462 10052
rect 10518 9996 11788 10052
rect 11844 9996 11854 10052
rect 23884 9996 25676 10052
rect 25732 9996 25742 10052
rect 26852 9996 27916 10052
rect 27972 9996 27982 10052
rect 26852 9940 26908 9996
rect 7858 9884 7868 9940
rect 7924 9884 9660 9940
rect 9716 9884 9726 9940
rect 12954 9884 12964 9940
rect 13020 9884 15484 9940
rect 15540 9884 15550 9940
rect 20458 9884 20468 9940
rect 20524 9884 26908 9940
rect 8194 9772 8204 9828
rect 8260 9772 8988 9828
rect 9044 9772 9054 9828
rect 21858 9772 21868 9828
rect 21924 9772 22428 9828
rect 22484 9772 22494 9828
rect 25106 9772 25116 9828
rect 25172 9772 26124 9828
rect 26180 9772 26190 9828
rect 28354 9772 28364 9828
rect 28420 9772 29148 9828
rect 29204 9772 32620 9828
rect 32676 9772 32686 9828
rect 32834 9772 32844 9828
rect 32900 9772 37902 9828
rect 37958 9772 37968 9828
rect 8082 9660 8092 9716
rect 8148 9660 8746 9716
rect 8802 9660 8812 9716
rect 12786 9660 12796 9716
rect 12852 9660 13524 9716
rect 13580 9660 13590 9716
rect 26786 9660 26796 9716
rect 26852 9604 26908 9716
rect 16930 9548 16940 9604
rect 16996 9548 17556 9604
rect 17612 9548 20076 9604
rect 20132 9548 20468 9604
rect 20524 9548 20534 9604
rect 26852 9548 27132 9604
rect 27188 9548 30380 9604
rect 30436 9548 30446 9604
rect 31938 9548 31948 9604
rect 32004 9548 32340 9604
rect 32396 9548 32956 9604
rect 33012 9548 33628 9604
rect 33684 9548 34972 9604
rect 35028 9548 35252 9604
rect 35308 9548 35318 9604
rect 10526 9380 10536 9436
rect 10592 9380 10640 9436
rect 10696 9380 10744 9436
rect 10800 9380 10810 9436
rect 19850 9380 19860 9436
rect 19916 9380 19964 9436
rect 20020 9380 20068 9436
rect 20124 9380 20134 9436
rect 29174 9380 29184 9436
rect 29240 9380 29288 9436
rect 29344 9380 29392 9436
rect 29448 9380 29458 9436
rect 38498 9380 38508 9436
rect 38564 9380 38612 9436
rect 38668 9380 38716 9436
rect 38772 9380 38782 9436
rect 26852 9324 29092 9380
rect 26852 9268 26908 9324
rect 29036 9268 29092 9324
rect 15474 9212 15484 9268
rect 15540 9212 18228 9268
rect 18284 9212 21980 9268
rect 22036 9212 22046 9268
rect 22754 9212 22764 9268
rect 22820 9212 26908 9268
rect 27804 9212 28364 9268
rect 28420 9212 28430 9268
rect 29036 9212 35812 9268
rect 35970 9212 35980 9268
rect 36036 9212 37156 9268
rect 37212 9212 37222 9268
rect 27804 9156 27860 9212
rect 35756 9156 35812 9212
rect 9538 9100 9548 9156
rect 9604 9100 9996 9156
rect 10052 9100 10062 9156
rect 26450 9100 26460 9156
rect 26516 9100 27804 9156
rect 27860 9100 27870 9156
rect 30370 9100 30380 9156
rect 30436 9100 31500 9156
rect 31556 9100 31566 9156
rect 35756 9100 38108 9156
rect 38164 9100 38174 9156
rect 28112 8988 28122 9044
rect 28178 8988 30212 9044
rect 30268 8988 30278 9044
rect 30706 8988 30716 9044
rect 30772 8988 31612 9044
rect 31668 8988 32060 9044
rect 32116 8988 32126 9044
rect 7074 8764 7084 8820
rect 7140 8764 8204 8820
rect 8260 8764 8270 8820
rect 18722 8764 18732 8820
rect 18788 8764 19180 8820
rect 19236 8764 19246 8820
rect 25984 8764 25994 8820
rect 26050 8764 27020 8820
rect 27076 8764 27086 8820
rect 32162 8764 32172 8820
rect 32228 8764 33292 8820
rect 33348 8764 37324 8820
rect 37380 8764 37390 8820
rect 36988 8708 37044 8764
rect 36978 8652 36988 8708
rect 37044 8652 37054 8708
rect 5864 8596 5874 8652
rect 5930 8596 5978 8652
rect 6034 8596 6082 8652
rect 6138 8596 6148 8652
rect 15188 8596 15198 8652
rect 15254 8596 15302 8652
rect 15358 8596 15406 8652
rect 15462 8596 15472 8652
rect 24512 8596 24522 8652
rect 24578 8596 24626 8652
rect 24682 8596 24730 8652
rect 24786 8596 24796 8652
rect 33836 8596 33846 8652
rect 33902 8596 33950 8652
rect 34006 8596 34054 8652
rect 34110 8596 34120 8652
rect 8642 8540 8652 8596
rect 8708 8540 8718 8596
rect 8652 8372 8708 8540
rect 21858 8428 21868 8484
rect 21924 8428 24892 8484
rect 24948 8428 24958 8484
rect 36642 8428 36652 8484
rect 36708 8428 37548 8484
rect 37604 8428 37614 8484
rect 39200 8372 40000 8400
rect 7298 8316 7308 8372
rect 7364 8316 9660 8372
rect 9716 8316 9726 8372
rect 26898 8316 26908 8372
rect 26964 8316 27468 8372
rect 27524 8316 27534 8372
rect 34402 8316 34412 8372
rect 34468 8316 37902 8372
rect 37958 8316 37968 8372
rect 38322 8316 38332 8372
rect 38388 8316 40000 8372
rect 39200 8288 40000 8316
rect 12450 8204 12460 8260
rect 12516 8204 13804 8260
rect 13860 8204 13870 8260
rect 20066 8204 20076 8260
rect 20132 8204 21756 8260
rect 21812 8204 22204 8260
rect 22260 8204 28588 8260
rect 28644 8204 29036 8260
rect 29092 8204 29102 8260
rect 30930 8204 30940 8260
rect 30996 8204 32172 8260
rect 32228 8204 32238 8260
rect 35746 8204 35756 8260
rect 35812 8204 37660 8260
rect 37716 8204 37726 8260
rect 8306 8092 8316 8148
rect 8372 8092 8540 8148
rect 8596 8092 8606 8148
rect 34682 8092 34692 8148
rect 34748 8092 35532 8148
rect 35588 8092 35598 8148
rect 9426 7980 9436 8036
rect 9492 7980 9940 8036
rect 9996 7980 11060 8036
rect 11116 7980 11126 8036
rect 17154 7980 17164 8036
rect 17220 7980 17780 8036
rect 17836 7980 17846 8036
rect 35242 7980 35252 8036
rect 35308 7980 36204 8036
rect 36260 7980 37324 8036
rect 37380 7980 37390 8036
rect 10526 7812 10536 7868
rect 10592 7812 10640 7868
rect 10696 7812 10744 7868
rect 10800 7812 10810 7868
rect 19850 7812 19860 7868
rect 19916 7812 19964 7868
rect 20020 7812 20068 7868
rect 20124 7812 20134 7868
rect 29174 7812 29184 7868
rect 29240 7812 29288 7868
rect 29344 7812 29392 7868
rect 29448 7812 29458 7868
rect 38498 7812 38508 7868
rect 38564 7812 38612 7868
rect 38668 7812 38716 7868
rect 38772 7812 38782 7868
rect 11050 7756 11060 7812
rect 11116 7756 16604 7812
rect 16660 7756 16670 7812
rect 13906 7644 13916 7700
rect 13972 7644 13982 7700
rect 23314 7644 23324 7700
rect 23380 7644 25434 7700
rect 25490 7644 25500 7700
rect 35204 7644 35214 7700
rect 35270 7644 37156 7700
rect 37212 7644 37222 7700
rect 8306 7532 8316 7588
rect 8372 7532 9044 7588
rect 9100 7532 9110 7588
rect 13916 7476 13972 7644
rect 26338 7532 26348 7588
rect 26404 7532 28588 7588
rect 28644 7532 29036 7588
rect 29092 7532 30268 7588
rect 30324 7532 30604 7588
rect 30660 7532 30670 7588
rect 8138 7420 8148 7476
rect 8204 7420 9940 7476
rect 9996 7420 10006 7476
rect 10882 7420 10892 7476
rect 10948 7420 11900 7476
rect 11956 7420 11966 7476
rect 12114 7420 12124 7476
rect 12180 7420 14588 7476
rect 14644 7420 14654 7476
rect 15138 7420 15148 7476
rect 15204 7420 15540 7476
rect 15596 7420 17108 7476
rect 17164 7420 17276 7476
rect 17332 7420 17342 7476
rect 24546 7420 24556 7476
rect 24612 7420 25676 7476
rect 25732 7420 27356 7476
rect 27412 7420 27422 7476
rect 32498 7420 32508 7476
rect 32564 7420 34300 7476
rect 34356 7420 35084 7476
rect 35140 7420 35150 7476
rect 37762 7420 37772 7476
rect 37828 7420 38332 7476
rect 38388 7420 38398 7476
rect 8530 7308 8540 7364
rect 8596 7308 9436 7364
rect 9492 7308 9502 7364
rect 26842 7308 26852 7364
rect 26908 7308 27468 7364
rect 27524 7308 27534 7364
rect 34458 7308 34468 7364
rect 34524 7308 37436 7364
rect 37492 7308 37502 7364
rect 7970 7196 7980 7252
rect 8036 7196 8428 7252
rect 8484 7196 8494 7252
rect 5864 7028 5874 7084
rect 5930 7028 5978 7084
rect 6034 7028 6082 7084
rect 6138 7028 6148 7084
rect 15188 7028 15198 7084
rect 15254 7028 15302 7084
rect 15358 7028 15406 7084
rect 15462 7028 15472 7084
rect 24512 7028 24522 7084
rect 24578 7028 24626 7084
rect 24682 7028 24730 7084
rect 24786 7028 24796 7084
rect 33836 7028 33846 7084
rect 33902 7028 33950 7084
rect 34006 7028 34054 7084
rect 34110 7028 34120 7084
rect 15344 6860 15354 6916
rect 15410 6860 16716 6916
rect 16772 6860 16782 6916
rect 27010 6860 27020 6916
rect 27076 6860 29484 6916
rect 29540 6860 30044 6916
rect 30100 6860 30604 6916
rect 30660 6860 30670 6916
rect 6514 6748 6524 6804
rect 6580 6748 8540 6804
rect 8596 6748 8606 6804
rect 10892 6748 12460 6804
rect 12516 6748 12526 6804
rect 19002 6748 19012 6804
rect 19068 6748 19964 6804
rect 20020 6748 20030 6804
rect 8884 6636 8894 6692
rect 8950 6636 10668 6692
rect 10724 6636 10734 6692
rect 8642 6524 8652 6580
rect 8708 6524 9548 6580
rect 9604 6524 9614 6580
rect 10892 6468 10948 6748
rect 15586 6636 15596 6692
rect 15652 6636 15662 6692
rect 16258 6636 16268 6692
rect 16324 6636 18844 6692
rect 18900 6636 19180 6692
rect 19236 6636 19246 6692
rect 19748 6636 19758 6692
rect 19814 6636 20300 6692
rect 20356 6636 20366 6692
rect 22866 6636 22876 6692
rect 22932 6636 23996 6692
rect 24052 6636 24062 6692
rect 28354 6636 28364 6692
rect 28420 6636 30156 6692
rect 30212 6636 30222 6692
rect 33954 6636 33964 6692
rect 34020 6636 35644 6692
rect 35700 6636 35710 6692
rect 15596 6580 15652 6636
rect 15596 6524 18060 6580
rect 18116 6524 19012 6580
rect 19068 6524 19078 6580
rect 19506 6524 19516 6580
rect 19572 6524 21084 6580
rect 21140 6524 21150 6580
rect 29596 6468 29652 6636
rect 29810 6524 29820 6580
rect 29876 6524 30716 6580
rect 30772 6524 31948 6580
rect 32004 6524 32014 6580
rect 32162 6524 32172 6580
rect 32228 6524 34206 6580
rect 34262 6524 34272 6580
rect 35186 6524 35196 6580
rect 35252 6524 37660 6580
rect 37716 6524 38108 6580
rect 38164 6524 38174 6580
rect 31948 6468 32004 6524
rect 10098 6412 10108 6468
rect 10164 6412 10948 6468
rect 16930 6412 16940 6468
rect 16996 6412 17948 6468
rect 18004 6412 20076 6468
rect 20132 6412 20142 6468
rect 20290 6412 20300 6468
rect 20356 6412 21420 6468
rect 21476 6412 21486 6468
rect 29586 6412 29596 6468
rect 29652 6412 29662 6468
rect 31948 6412 34076 6468
rect 34132 6412 34142 6468
rect 29698 6300 29708 6356
rect 29764 6300 29932 6356
rect 29988 6300 32284 6356
rect 32340 6300 32350 6356
rect 10526 6244 10536 6300
rect 10592 6244 10640 6300
rect 10696 6244 10744 6300
rect 10800 6244 10810 6300
rect 19850 6244 19860 6300
rect 19916 6244 19964 6300
rect 20020 6244 20068 6300
rect 20124 6244 20134 6300
rect 29174 6244 29184 6300
rect 29240 6244 29288 6300
rect 29344 6244 29392 6300
rect 29448 6244 29458 6300
rect 38498 6244 38508 6300
rect 38564 6244 38612 6300
rect 38668 6244 38716 6300
rect 38772 6244 38782 6300
rect 9986 6076 9996 6132
rect 10052 6076 14476 6132
rect 14532 6076 15820 6132
rect 15876 6076 15886 6132
rect 16090 6076 16100 6132
rect 16156 6076 16492 6132
rect 16548 6076 17500 6132
rect 17556 6076 18172 6132
rect 18228 6076 18238 6132
rect 28690 6076 28700 6132
rect 28756 6076 30212 6132
rect 30268 6076 30278 6132
rect 35970 6076 35980 6132
rect 36036 6076 37156 6132
rect 37212 6076 37222 6132
rect 10434 5964 10444 6020
rect 10500 5964 13692 6020
rect 13748 5964 14140 6020
rect 14196 5964 14206 6020
rect 19170 5964 19180 6020
rect 19236 5964 21420 6020
rect 21476 5964 21486 6020
rect 21746 5964 21756 6020
rect 21812 5964 22092 6020
rect 22148 5964 25228 6020
rect 25284 5964 25294 6020
rect 27570 5964 27580 6020
rect 27636 5964 28868 6020
rect 28924 5964 28934 6020
rect 34850 5964 34860 6020
rect 34916 5964 37902 6020
rect 37958 5964 37968 6020
rect 5842 5852 5852 5908
rect 5908 5852 11004 5908
rect 11060 5852 11070 5908
rect 22754 5852 22764 5908
rect 22820 5852 22830 5908
rect 24322 5852 24332 5908
rect 24388 5852 28122 5908
rect 28178 5852 28188 5908
rect 28354 5852 28364 5908
rect 28420 5852 29708 5908
rect 29764 5852 29774 5908
rect 34178 5852 34188 5908
rect 34244 5852 34636 5908
rect 34692 5852 34702 5908
rect 22764 5796 22820 5852
rect 22764 5740 23772 5796
rect 23828 5740 24108 5796
rect 24164 5740 25788 5796
rect 25844 5740 25854 5796
rect 13570 5628 13580 5684
rect 13636 5628 15148 5684
rect 15204 5628 15214 5684
rect 17378 5628 17388 5684
rect 17444 5628 18508 5684
rect 18564 5628 18574 5684
rect 24322 5628 24332 5684
rect 24388 5628 26236 5684
rect 26292 5628 26302 5684
rect 5864 5460 5874 5516
rect 5930 5460 5978 5516
rect 6034 5460 6082 5516
rect 6138 5460 6148 5516
rect 15188 5460 15198 5516
rect 15254 5460 15302 5516
rect 15358 5460 15406 5516
rect 15462 5460 15472 5516
rect 24512 5460 24522 5516
rect 24578 5460 24626 5516
rect 24682 5460 24730 5516
rect 24786 5460 24796 5516
rect 33836 5460 33846 5516
rect 33902 5460 33950 5516
rect 34006 5460 34054 5516
rect 34110 5460 34120 5516
rect 39200 5460 40000 5488
rect 31378 5404 31388 5460
rect 31444 5404 32620 5460
rect 32676 5404 33404 5460
rect 33460 5404 33470 5460
rect 38322 5404 38332 5460
rect 38388 5404 40000 5460
rect 39200 5376 40000 5404
rect 26852 5292 37996 5348
rect 38052 5292 38062 5348
rect 26852 5236 26908 5292
rect 6178 5180 6188 5236
rect 6244 5180 8316 5236
rect 8372 5180 8382 5236
rect 8978 5180 8988 5236
rect 9044 5180 10220 5236
rect 10276 5180 10286 5236
rect 14242 5180 14252 5236
rect 14308 5180 16268 5236
rect 16324 5180 16334 5236
rect 19618 5180 19628 5236
rect 19684 5180 26908 5236
rect 27458 5180 27468 5236
rect 27524 5180 28364 5236
rect 28420 5180 28430 5236
rect 35410 5180 35420 5236
rect 35476 5180 36260 5236
rect 36316 5180 37156 5236
rect 37212 5180 38220 5236
rect 38276 5180 38286 5236
rect 4162 5068 4172 5124
rect 4228 5068 9100 5124
rect 9156 5068 9166 5124
rect 10994 5068 11004 5124
rect 11060 5068 12572 5124
rect 12628 5068 12638 5124
rect 15474 5068 15484 5124
rect 15540 5068 16884 5124
rect 23146 5068 23156 5124
rect 23212 5068 23660 5124
rect 23716 5068 23726 5124
rect 26236 5068 27916 5124
rect 27972 5068 27982 5124
rect 16828 5012 16884 5068
rect 3490 4956 3500 5012
rect 3556 4956 10332 5012
rect 10388 4956 10398 5012
rect 16828 4956 18788 5012
rect 18844 4956 18854 5012
rect 26236 4900 26292 5068
rect 7634 4844 7644 4900
rect 7700 4844 8428 4900
rect 26226 4844 26236 4900
rect 26292 4844 26302 4900
rect 8372 4788 8428 4844
rect 8372 4732 10108 4788
rect 10164 4732 10174 4788
rect 10526 4676 10536 4732
rect 10592 4676 10640 4732
rect 10696 4676 10744 4732
rect 10800 4676 10810 4732
rect 19850 4676 19860 4732
rect 19916 4676 19964 4732
rect 20020 4676 20068 4732
rect 20124 4676 20134 4732
rect 29174 4676 29184 4732
rect 29240 4676 29288 4732
rect 29344 4676 29392 4732
rect 29448 4676 29458 4732
rect 38498 4676 38508 4732
rect 38564 4676 38612 4732
rect 38668 4676 38716 4732
rect 38772 4676 38782 4732
rect 2762 4508 2772 4564
rect 2828 4508 3500 4564
rect 3556 4508 3566 4564
rect 13794 4508 13804 4564
rect 13860 4508 13972 4564
rect 13916 4340 13972 4508
rect 15362 4396 15372 4452
rect 15428 4396 17444 4452
rect 17500 4396 17510 4452
rect 11890 4284 11900 4340
rect 11956 4284 13356 4340
rect 13412 4284 13422 4340
rect 13916 4284 15260 4340
rect 15316 4284 15988 4340
rect 16044 4284 16054 4340
rect 16724 4284 16734 4340
rect 16790 4284 17724 4340
rect 17780 4284 17790 4340
rect 22530 4284 22540 4340
rect 22596 4284 23660 4340
rect 23716 4284 23726 4340
rect 24434 4284 24444 4340
rect 24500 4284 26908 4340
rect 26964 4284 29932 4340
rect 29988 4284 29998 4340
rect 6514 4060 6524 4116
rect 6580 4060 7532 4116
rect 7588 4060 7598 4116
rect 13916 4004 13972 4284
rect 13906 3948 13916 4004
rect 13972 3948 13982 4004
rect 5864 3892 5874 3948
rect 5930 3892 5978 3948
rect 6034 3892 6082 3948
rect 6138 3892 6148 3948
rect 15188 3892 15198 3948
rect 15254 3892 15302 3948
rect 15358 3892 15406 3948
rect 15462 3892 15472 3948
rect 24512 3892 24522 3948
rect 24578 3892 24626 3948
rect 24682 3892 24730 3948
rect 24786 3892 24796 3948
rect 33836 3892 33846 3948
rect 33902 3892 33950 3948
rect 34006 3892 34054 3948
rect 34110 3892 34120 3948
rect 20962 3724 20972 3780
rect 21028 3724 21196 3780
rect 21252 3724 24556 3780
rect 24612 3724 24622 3780
rect 35242 3724 35252 3780
rect 35308 3724 36204 3780
rect 36260 3724 36270 3780
rect 20850 3612 20860 3668
rect 20916 3612 22092 3668
rect 22148 3612 22158 3668
rect 22642 3612 22652 3668
rect 22708 3612 25564 3668
rect 25620 3612 25630 3668
rect 13570 3500 13580 3556
rect 13636 3500 14588 3556
rect 14644 3500 14654 3556
rect 26226 3500 26236 3556
rect 26292 3500 27804 3556
rect 27860 3500 27870 3556
rect 28018 3500 28028 3556
rect 28084 3500 28812 3556
rect 28868 3500 29652 3556
rect 29708 3500 29718 3556
rect 29810 3500 29820 3556
rect 29876 3500 30492 3556
rect 30548 3500 30884 3556
rect 30940 3500 30950 3556
rect 27804 3444 27860 3500
rect 1138 3388 1148 3444
rect 1204 3388 1932 3444
rect 1988 3388 1998 3444
rect 2930 3388 2940 3444
rect 2996 3388 3500 3444
rect 3556 3388 3566 3444
rect 27804 3388 29204 3444
rect 29260 3388 29270 3444
rect 10526 3108 10536 3164
rect 10592 3108 10640 3164
rect 10696 3108 10744 3164
rect 10800 3108 10810 3164
rect 19850 3108 19860 3164
rect 19916 3108 19964 3164
rect 20020 3108 20068 3164
rect 20124 3108 20134 3164
rect 29174 3108 29184 3164
rect 29240 3108 29288 3164
rect 29344 3108 29392 3164
rect 29448 3108 29458 3164
rect 38498 3108 38508 3164
rect 38564 3108 38612 3164
rect 38668 3108 38716 3164
rect 38772 3108 38782 3164
rect 39200 2548 40000 2576
rect 24210 2492 24220 2548
rect 24276 2492 40000 2548
rect 39200 2464 40000 2492
rect 10098 812 10108 868
rect 10164 812 10892 868
rect 10948 812 10958 868
<< via3 >>
rect 5874 36820 5930 36876
rect 5978 36820 6034 36876
rect 6082 36820 6138 36876
rect 15198 36820 15254 36876
rect 15302 36820 15358 36876
rect 15406 36820 15462 36876
rect 24522 36820 24578 36876
rect 24626 36820 24682 36876
rect 24730 36820 24786 36876
rect 33846 36820 33902 36876
rect 33950 36820 34006 36876
rect 34054 36820 34110 36876
rect 10536 36036 10592 36092
rect 10640 36036 10696 36092
rect 10744 36036 10800 36092
rect 19860 36036 19916 36092
rect 19964 36036 20020 36092
rect 20068 36036 20124 36092
rect 29184 36036 29240 36092
rect 29288 36036 29344 36092
rect 29392 36036 29448 36092
rect 38508 36036 38564 36092
rect 38612 36036 38668 36092
rect 38716 36036 38772 36092
rect 26908 35308 26964 35364
rect 5874 35252 5930 35308
rect 5978 35252 6034 35308
rect 6082 35252 6138 35308
rect 15198 35252 15254 35308
rect 15302 35252 15358 35308
rect 15406 35252 15462 35308
rect 24522 35252 24578 35308
rect 24626 35252 24682 35308
rect 24730 35252 24786 35308
rect 33846 35252 33902 35308
rect 33950 35252 34006 35308
rect 34054 35252 34110 35308
rect 26908 34972 26964 35028
rect 35644 34972 35700 35028
rect 35308 34748 35364 34804
rect 10536 34468 10592 34524
rect 10640 34468 10696 34524
rect 10744 34468 10800 34524
rect 19860 34468 19916 34524
rect 19964 34468 20020 34524
rect 20068 34468 20124 34524
rect 29184 34468 29240 34524
rect 29288 34468 29344 34524
rect 29392 34468 29448 34524
rect 38508 34468 38564 34524
rect 38612 34468 38668 34524
rect 38716 34468 38772 34524
rect 35420 34412 35476 34468
rect 35644 33852 35700 33908
rect 5874 33684 5930 33740
rect 5978 33684 6034 33740
rect 6082 33684 6138 33740
rect 15198 33684 15254 33740
rect 15302 33684 15358 33740
rect 15406 33684 15462 33740
rect 24522 33684 24578 33740
rect 24626 33684 24682 33740
rect 24730 33684 24786 33740
rect 33846 33684 33902 33740
rect 33950 33684 34006 33740
rect 34054 33684 34110 33740
rect 35644 32956 35700 33012
rect 10536 32900 10592 32956
rect 10640 32900 10696 32956
rect 10744 32900 10800 32956
rect 19860 32900 19916 32956
rect 19964 32900 20020 32956
rect 20068 32900 20124 32956
rect 29184 32900 29240 32956
rect 29288 32900 29344 32956
rect 29392 32900 29448 32956
rect 38508 32900 38564 32956
rect 38612 32900 38668 32956
rect 38716 32900 38772 32956
rect 31724 32844 31780 32900
rect 21756 32732 21812 32788
rect 5874 32116 5930 32172
rect 5978 32116 6034 32172
rect 6082 32116 6138 32172
rect 15198 32116 15254 32172
rect 15302 32116 15358 32172
rect 15406 32116 15462 32172
rect 24522 32116 24578 32172
rect 24626 32116 24682 32172
rect 24730 32116 24786 32172
rect 33846 32116 33902 32172
rect 33950 32116 34006 32172
rect 34054 32116 34110 32172
rect 15596 32060 15652 32116
rect 24108 31948 24164 32004
rect 15036 31836 15092 31892
rect 35420 31724 35476 31780
rect 37100 31388 37156 31444
rect 10536 31332 10592 31388
rect 10640 31332 10696 31388
rect 10744 31332 10800 31388
rect 19860 31332 19916 31388
rect 19964 31332 20020 31388
rect 20068 31332 20124 31388
rect 29184 31332 29240 31388
rect 29288 31332 29344 31388
rect 29392 31332 29448 31388
rect 38508 31332 38564 31388
rect 38612 31332 38668 31388
rect 38716 31332 38772 31388
rect 37660 31052 37716 31108
rect 26684 30940 26740 30996
rect 26684 30716 26740 30772
rect 15036 30604 15092 30660
rect 5874 30548 5930 30604
rect 5978 30548 6034 30604
rect 6082 30548 6138 30604
rect 15198 30548 15254 30604
rect 15302 30548 15358 30604
rect 15406 30548 15462 30604
rect 12236 30492 12292 30548
rect 24522 30548 24578 30604
rect 24626 30548 24682 30604
rect 24730 30548 24786 30604
rect 33846 30548 33902 30604
rect 33950 30548 34006 30604
rect 34054 30548 34110 30604
rect 29596 30156 29652 30212
rect 15596 29820 15652 29876
rect 10536 29764 10592 29820
rect 10640 29764 10696 29820
rect 10744 29764 10800 29820
rect 19860 29764 19916 29820
rect 19964 29764 20020 29820
rect 20068 29764 20124 29820
rect 29184 29764 29240 29820
rect 29288 29764 29344 29820
rect 29392 29764 29448 29820
rect 38508 29764 38564 29820
rect 38612 29764 38668 29820
rect 38716 29764 38772 29820
rect 30940 29596 30996 29652
rect 37100 29596 37156 29652
rect 12236 29484 12292 29540
rect 29596 29484 29652 29540
rect 19628 29260 19684 29316
rect 31612 29148 31668 29204
rect 10892 29036 10948 29092
rect 5874 28980 5930 29036
rect 5978 28980 6034 29036
rect 6082 28980 6138 29036
rect 15198 28980 15254 29036
rect 15302 28980 15358 29036
rect 15406 28980 15462 29036
rect 24522 28980 24578 29036
rect 24626 28980 24682 29036
rect 24730 28980 24786 29036
rect 33846 28980 33902 29036
rect 33950 28980 34006 29036
rect 34054 28980 34110 29036
rect 29596 28812 29652 28868
rect 37660 28364 37716 28420
rect 10536 28196 10592 28252
rect 10640 28196 10696 28252
rect 10744 28196 10800 28252
rect 19860 28196 19916 28252
rect 19964 28196 20020 28252
rect 20068 28196 20124 28252
rect 29184 28196 29240 28252
rect 29288 28196 29344 28252
rect 29392 28196 29448 28252
rect 38508 28196 38564 28252
rect 38612 28196 38668 28252
rect 38716 28196 38772 28252
rect 19404 28028 19460 28084
rect 21756 28028 21812 28084
rect 29596 27804 29652 27860
rect 31612 27804 31668 27860
rect 18956 27580 19012 27636
rect 30940 27580 30996 27636
rect 5874 27412 5930 27468
rect 5978 27412 6034 27468
rect 6082 27412 6138 27468
rect 15198 27412 15254 27468
rect 15302 27412 15358 27468
rect 15406 27412 15462 27468
rect 24522 27412 24578 27468
rect 24626 27412 24682 27468
rect 24730 27412 24786 27468
rect 33846 27412 33902 27468
rect 33950 27412 34006 27468
rect 34054 27412 34110 27468
rect 19404 27020 19460 27076
rect 10892 26796 10948 26852
rect 10536 26628 10592 26684
rect 10640 26628 10696 26684
rect 10744 26628 10800 26684
rect 19860 26628 19916 26684
rect 19964 26628 20020 26684
rect 20068 26628 20124 26684
rect 29184 26628 29240 26684
rect 29288 26628 29344 26684
rect 29392 26628 29448 26684
rect 38508 26628 38564 26684
rect 38612 26628 38668 26684
rect 38716 26628 38772 26684
rect 19628 26572 19684 26628
rect 20300 26572 20356 26628
rect 5874 25844 5930 25900
rect 5978 25844 6034 25900
rect 6082 25844 6138 25900
rect 15198 25844 15254 25900
rect 15302 25844 15358 25900
rect 15406 25844 15462 25900
rect 24522 25844 24578 25900
rect 24626 25844 24682 25900
rect 24730 25844 24786 25900
rect 33846 25844 33902 25900
rect 33950 25844 34006 25900
rect 34054 25844 34110 25900
rect 19404 25788 19460 25844
rect 20300 25564 20356 25620
rect 35420 25452 35476 25508
rect 35644 25340 35700 25396
rect 10536 25060 10592 25116
rect 10640 25060 10696 25116
rect 10744 25060 10800 25116
rect 19860 25060 19916 25116
rect 19964 25060 20020 25116
rect 20068 25060 20124 25116
rect 29184 25060 29240 25116
rect 29288 25060 29344 25116
rect 29392 25060 29448 25116
rect 38508 25060 38564 25116
rect 38612 25060 38668 25116
rect 38716 25060 38772 25116
rect 24108 24892 24164 24948
rect 20300 24668 20356 24724
rect 31724 24332 31780 24388
rect 5874 24276 5930 24332
rect 5978 24276 6034 24332
rect 6082 24276 6138 24332
rect 15198 24276 15254 24332
rect 15302 24276 15358 24332
rect 15406 24276 15462 24332
rect 24522 24276 24578 24332
rect 24626 24276 24682 24332
rect 24730 24276 24786 24332
rect 33846 24276 33902 24332
rect 33950 24276 34006 24332
rect 34054 24276 34110 24332
rect 18172 24220 18228 24276
rect 24108 24220 24164 24276
rect 35420 23996 35476 24052
rect 35644 23996 35700 24052
rect 18956 23772 19012 23828
rect 18172 23548 18228 23604
rect 10536 23492 10592 23548
rect 10640 23492 10696 23548
rect 10744 23492 10800 23548
rect 19860 23492 19916 23548
rect 19964 23492 20020 23548
rect 20068 23492 20124 23548
rect 29184 23492 29240 23548
rect 29288 23492 29344 23548
rect 29392 23492 29448 23548
rect 38508 23492 38564 23548
rect 38612 23492 38668 23548
rect 38716 23492 38772 23548
rect 5874 22708 5930 22764
rect 5978 22708 6034 22764
rect 6082 22708 6138 22764
rect 15198 22708 15254 22764
rect 15302 22708 15358 22764
rect 15406 22708 15462 22764
rect 24522 22708 24578 22764
rect 24626 22708 24682 22764
rect 24730 22708 24786 22764
rect 33846 22708 33902 22764
rect 33950 22708 34006 22764
rect 34054 22708 34110 22764
rect 10536 21924 10592 21980
rect 10640 21924 10696 21980
rect 10744 21924 10800 21980
rect 19860 21924 19916 21980
rect 19964 21924 20020 21980
rect 20068 21924 20124 21980
rect 29184 21924 29240 21980
rect 29288 21924 29344 21980
rect 29392 21924 29448 21980
rect 38508 21924 38564 21980
rect 38612 21924 38668 21980
rect 38716 21924 38772 21980
rect 5874 21140 5930 21196
rect 5978 21140 6034 21196
rect 6082 21140 6138 21196
rect 15198 21140 15254 21196
rect 15302 21140 15358 21196
rect 15406 21140 15462 21196
rect 24522 21140 24578 21196
rect 24626 21140 24682 21196
rect 24730 21140 24786 21196
rect 33846 21140 33902 21196
rect 33950 21140 34006 21196
rect 34054 21140 34110 21196
rect 10536 20356 10592 20412
rect 10640 20356 10696 20412
rect 10744 20356 10800 20412
rect 19860 20356 19916 20412
rect 19964 20356 20020 20412
rect 20068 20356 20124 20412
rect 29184 20356 29240 20412
rect 29288 20356 29344 20412
rect 29392 20356 29448 20412
rect 38508 20356 38564 20412
rect 38612 20356 38668 20412
rect 38716 20356 38772 20412
rect 35308 20188 35364 20244
rect 5874 19572 5930 19628
rect 5978 19572 6034 19628
rect 6082 19572 6138 19628
rect 15198 19572 15254 19628
rect 15302 19572 15358 19628
rect 15406 19572 15462 19628
rect 24522 19572 24578 19628
rect 24626 19572 24682 19628
rect 24730 19572 24786 19628
rect 33846 19572 33902 19628
rect 33950 19572 34006 19628
rect 34054 19572 34110 19628
rect 10536 18788 10592 18844
rect 10640 18788 10696 18844
rect 10744 18788 10800 18844
rect 19860 18788 19916 18844
rect 19964 18788 20020 18844
rect 20068 18788 20124 18844
rect 29184 18788 29240 18844
rect 29288 18788 29344 18844
rect 29392 18788 29448 18844
rect 38508 18788 38564 18844
rect 38612 18788 38668 18844
rect 38716 18788 38772 18844
rect 5874 18004 5930 18060
rect 5978 18004 6034 18060
rect 6082 18004 6138 18060
rect 15198 18004 15254 18060
rect 15302 18004 15358 18060
rect 15406 18004 15462 18060
rect 24522 18004 24578 18060
rect 24626 18004 24682 18060
rect 24730 18004 24786 18060
rect 33846 18004 33902 18060
rect 33950 18004 34006 18060
rect 34054 18004 34110 18060
rect 10536 17220 10592 17276
rect 10640 17220 10696 17276
rect 10744 17220 10800 17276
rect 19860 17220 19916 17276
rect 19964 17220 20020 17276
rect 20068 17220 20124 17276
rect 29184 17220 29240 17276
rect 29288 17220 29344 17276
rect 29392 17220 29448 17276
rect 38508 17220 38564 17276
rect 38612 17220 38668 17276
rect 38716 17220 38772 17276
rect 25452 17164 25508 17220
rect 5874 16436 5930 16492
rect 5978 16436 6034 16492
rect 6082 16436 6138 16492
rect 15198 16436 15254 16492
rect 15302 16436 15358 16492
rect 15406 16436 15462 16492
rect 24522 16436 24578 16492
rect 24626 16436 24682 16492
rect 24730 16436 24786 16492
rect 33846 16436 33902 16492
rect 33950 16436 34006 16492
rect 34054 16436 34110 16492
rect 25452 16044 25508 16100
rect 10536 15652 10592 15708
rect 10640 15652 10696 15708
rect 10744 15652 10800 15708
rect 19860 15652 19916 15708
rect 19964 15652 20020 15708
rect 20068 15652 20124 15708
rect 29184 15652 29240 15708
rect 29288 15652 29344 15708
rect 29392 15652 29448 15708
rect 38508 15652 38564 15708
rect 38612 15652 38668 15708
rect 38716 15652 38772 15708
rect 34300 15036 34356 15092
rect 5874 14868 5930 14924
rect 5978 14868 6034 14924
rect 6082 14868 6138 14924
rect 15198 14868 15254 14924
rect 15302 14868 15358 14924
rect 15406 14868 15462 14924
rect 24522 14868 24578 14924
rect 24626 14868 24682 14924
rect 24730 14868 24786 14924
rect 33846 14868 33902 14924
rect 33950 14868 34006 14924
rect 34054 14868 34110 14924
rect 10536 14084 10592 14140
rect 10640 14084 10696 14140
rect 10744 14084 10800 14140
rect 19860 14084 19916 14140
rect 19964 14084 20020 14140
rect 20068 14084 20124 14140
rect 29184 14084 29240 14140
rect 29288 14084 29344 14140
rect 29392 14084 29448 14140
rect 38508 14084 38564 14140
rect 38612 14084 38668 14140
rect 38716 14084 38772 14140
rect 31612 13692 31668 13748
rect 33628 13580 33684 13636
rect 5874 13300 5930 13356
rect 5978 13300 6034 13356
rect 6082 13300 6138 13356
rect 15198 13300 15254 13356
rect 15302 13300 15358 13356
rect 15406 13300 15462 13356
rect 24522 13300 24578 13356
rect 24626 13300 24682 13356
rect 24730 13300 24786 13356
rect 33846 13300 33902 13356
rect 33950 13300 34006 13356
rect 34054 13300 34110 13356
rect 34300 12796 34356 12852
rect 31612 12684 31668 12740
rect 33628 12684 33684 12740
rect 10536 12516 10592 12572
rect 10640 12516 10696 12572
rect 10744 12516 10800 12572
rect 19860 12516 19916 12572
rect 19964 12516 20020 12572
rect 20068 12516 20124 12572
rect 29184 12516 29240 12572
rect 29288 12516 29344 12572
rect 29392 12516 29448 12572
rect 38508 12516 38564 12572
rect 38612 12516 38668 12572
rect 38716 12516 38772 12572
rect 5874 11732 5930 11788
rect 5978 11732 6034 11788
rect 6082 11732 6138 11788
rect 15198 11732 15254 11788
rect 15302 11732 15358 11788
rect 15406 11732 15462 11788
rect 24522 11732 24578 11788
rect 24626 11732 24682 11788
rect 24730 11732 24786 11788
rect 33846 11732 33902 11788
rect 33950 11732 34006 11788
rect 34054 11732 34110 11788
rect 10536 10948 10592 11004
rect 10640 10948 10696 11004
rect 10744 10948 10800 11004
rect 19860 10948 19916 11004
rect 19964 10948 20020 11004
rect 20068 10948 20124 11004
rect 29184 10948 29240 11004
rect 29288 10948 29344 11004
rect 29392 10948 29448 11004
rect 38508 10948 38564 11004
rect 38612 10948 38668 11004
rect 38716 10948 38772 11004
rect 5874 10164 5930 10220
rect 5978 10164 6034 10220
rect 6082 10164 6138 10220
rect 15198 10164 15254 10220
rect 15302 10164 15358 10220
rect 15406 10164 15462 10220
rect 24522 10164 24578 10220
rect 24626 10164 24682 10220
rect 24730 10164 24786 10220
rect 33846 10164 33902 10220
rect 33950 10164 34006 10220
rect 34054 10164 34110 10220
rect 10536 9380 10592 9436
rect 10640 9380 10696 9436
rect 10744 9380 10800 9436
rect 19860 9380 19916 9436
rect 19964 9380 20020 9436
rect 20068 9380 20124 9436
rect 29184 9380 29240 9436
rect 29288 9380 29344 9436
rect 29392 9380 29448 9436
rect 38508 9380 38564 9436
rect 38612 9380 38668 9436
rect 38716 9380 38772 9436
rect 5874 8596 5930 8652
rect 5978 8596 6034 8652
rect 6082 8596 6138 8652
rect 15198 8596 15254 8652
rect 15302 8596 15358 8652
rect 15406 8596 15462 8652
rect 24522 8596 24578 8652
rect 24626 8596 24682 8652
rect 24730 8596 24786 8652
rect 33846 8596 33902 8652
rect 33950 8596 34006 8652
rect 34054 8596 34110 8652
rect 10536 7812 10592 7868
rect 10640 7812 10696 7868
rect 10744 7812 10800 7868
rect 19860 7812 19916 7868
rect 19964 7812 20020 7868
rect 20068 7812 20124 7868
rect 29184 7812 29240 7868
rect 29288 7812 29344 7868
rect 29392 7812 29448 7868
rect 38508 7812 38564 7868
rect 38612 7812 38668 7868
rect 38716 7812 38772 7868
rect 5874 7028 5930 7084
rect 5978 7028 6034 7084
rect 6082 7028 6138 7084
rect 15198 7028 15254 7084
rect 15302 7028 15358 7084
rect 15406 7028 15462 7084
rect 24522 7028 24578 7084
rect 24626 7028 24682 7084
rect 24730 7028 24786 7084
rect 33846 7028 33902 7084
rect 33950 7028 34006 7084
rect 34054 7028 34110 7084
rect 10536 6244 10592 6300
rect 10640 6244 10696 6300
rect 10744 6244 10800 6300
rect 19860 6244 19916 6300
rect 19964 6244 20020 6300
rect 20068 6244 20124 6300
rect 29184 6244 29240 6300
rect 29288 6244 29344 6300
rect 29392 6244 29448 6300
rect 38508 6244 38564 6300
rect 38612 6244 38668 6300
rect 38716 6244 38772 6300
rect 5874 5460 5930 5516
rect 5978 5460 6034 5516
rect 6082 5460 6138 5516
rect 15198 5460 15254 5516
rect 15302 5460 15358 5516
rect 15406 5460 15462 5516
rect 24522 5460 24578 5516
rect 24626 5460 24682 5516
rect 24730 5460 24786 5516
rect 33846 5460 33902 5516
rect 33950 5460 34006 5516
rect 34054 5460 34110 5516
rect 10536 4676 10592 4732
rect 10640 4676 10696 4732
rect 10744 4676 10800 4732
rect 19860 4676 19916 4732
rect 19964 4676 20020 4732
rect 20068 4676 20124 4732
rect 29184 4676 29240 4732
rect 29288 4676 29344 4732
rect 29392 4676 29448 4732
rect 38508 4676 38564 4732
rect 38612 4676 38668 4732
rect 38716 4676 38772 4732
rect 5874 3892 5930 3948
rect 5978 3892 6034 3948
rect 6082 3892 6138 3948
rect 15198 3892 15254 3948
rect 15302 3892 15358 3948
rect 15406 3892 15462 3948
rect 24522 3892 24578 3948
rect 24626 3892 24682 3948
rect 24730 3892 24786 3948
rect 33846 3892 33902 3948
rect 33950 3892 34006 3948
rect 34054 3892 34110 3948
rect 10536 3108 10592 3164
rect 10640 3108 10696 3164
rect 10744 3108 10800 3164
rect 19860 3108 19916 3164
rect 19964 3108 20020 3164
rect 20068 3108 20124 3164
rect 29184 3108 29240 3164
rect 29288 3108 29344 3164
rect 29392 3108 29448 3164
rect 38508 3108 38564 3164
rect 38612 3108 38668 3164
rect 38716 3108 38772 3164
<< metal4 >>
rect 5846 36876 6166 36908
rect 5846 36820 5874 36876
rect 5930 36820 5978 36876
rect 6034 36820 6082 36876
rect 6138 36820 6166 36876
rect 5846 35308 6166 36820
rect 5846 35252 5874 35308
rect 5930 35252 5978 35308
rect 6034 35252 6082 35308
rect 6138 35252 6166 35308
rect 5846 33740 6166 35252
rect 5846 33684 5874 33740
rect 5930 33684 5978 33740
rect 6034 33684 6082 33740
rect 6138 33684 6166 33740
rect 5846 32172 6166 33684
rect 5846 32116 5874 32172
rect 5930 32116 5978 32172
rect 6034 32116 6082 32172
rect 6138 32116 6166 32172
rect 5846 30604 6166 32116
rect 5846 30548 5874 30604
rect 5930 30548 5978 30604
rect 6034 30548 6082 30604
rect 6138 30548 6166 30604
rect 5846 29036 6166 30548
rect 5846 28980 5874 29036
rect 5930 28980 5978 29036
rect 6034 28980 6082 29036
rect 6138 28980 6166 29036
rect 5846 27468 6166 28980
rect 5846 27412 5874 27468
rect 5930 27412 5978 27468
rect 6034 27412 6082 27468
rect 6138 27412 6166 27468
rect 5846 25900 6166 27412
rect 5846 25844 5874 25900
rect 5930 25844 5978 25900
rect 6034 25844 6082 25900
rect 6138 25844 6166 25900
rect 5846 24332 6166 25844
rect 5846 24276 5874 24332
rect 5930 24276 5978 24332
rect 6034 24276 6082 24332
rect 6138 24276 6166 24332
rect 5846 22764 6166 24276
rect 5846 22708 5874 22764
rect 5930 22708 5978 22764
rect 6034 22708 6082 22764
rect 6138 22708 6166 22764
rect 5846 21196 6166 22708
rect 5846 21140 5874 21196
rect 5930 21140 5978 21196
rect 6034 21140 6082 21196
rect 6138 21140 6166 21196
rect 5846 19628 6166 21140
rect 5846 19572 5874 19628
rect 5930 19572 5978 19628
rect 6034 19572 6082 19628
rect 6138 19572 6166 19628
rect 5846 18060 6166 19572
rect 5846 18004 5874 18060
rect 5930 18004 5978 18060
rect 6034 18004 6082 18060
rect 6138 18004 6166 18060
rect 5846 16492 6166 18004
rect 5846 16436 5874 16492
rect 5930 16436 5978 16492
rect 6034 16436 6082 16492
rect 6138 16436 6166 16492
rect 5846 14924 6166 16436
rect 5846 14868 5874 14924
rect 5930 14868 5978 14924
rect 6034 14868 6082 14924
rect 6138 14868 6166 14924
rect 5846 13356 6166 14868
rect 5846 13300 5874 13356
rect 5930 13300 5978 13356
rect 6034 13300 6082 13356
rect 6138 13300 6166 13356
rect 5846 11788 6166 13300
rect 5846 11732 5874 11788
rect 5930 11732 5978 11788
rect 6034 11732 6082 11788
rect 6138 11732 6166 11788
rect 5846 10220 6166 11732
rect 5846 10164 5874 10220
rect 5930 10164 5978 10220
rect 6034 10164 6082 10220
rect 6138 10164 6166 10220
rect 5846 8652 6166 10164
rect 5846 8596 5874 8652
rect 5930 8596 5978 8652
rect 6034 8596 6082 8652
rect 6138 8596 6166 8652
rect 5846 7084 6166 8596
rect 5846 7028 5874 7084
rect 5930 7028 5978 7084
rect 6034 7028 6082 7084
rect 6138 7028 6166 7084
rect 5846 5516 6166 7028
rect 5846 5460 5874 5516
rect 5930 5460 5978 5516
rect 6034 5460 6082 5516
rect 6138 5460 6166 5516
rect 5846 3948 6166 5460
rect 5846 3892 5874 3948
rect 5930 3892 5978 3948
rect 6034 3892 6082 3948
rect 6138 3892 6166 3948
rect 5846 3076 6166 3892
rect 10508 36092 10828 36908
rect 10508 36036 10536 36092
rect 10592 36036 10640 36092
rect 10696 36036 10744 36092
rect 10800 36036 10828 36092
rect 10508 34524 10828 36036
rect 10508 34468 10536 34524
rect 10592 34468 10640 34524
rect 10696 34468 10744 34524
rect 10800 34468 10828 34524
rect 10508 32956 10828 34468
rect 10508 32900 10536 32956
rect 10592 32900 10640 32956
rect 10696 32900 10744 32956
rect 10800 32900 10828 32956
rect 10508 31388 10828 32900
rect 15170 36876 15490 36908
rect 15170 36820 15198 36876
rect 15254 36820 15302 36876
rect 15358 36820 15406 36876
rect 15462 36820 15490 36876
rect 15170 35308 15490 36820
rect 15170 35252 15198 35308
rect 15254 35252 15302 35308
rect 15358 35252 15406 35308
rect 15462 35252 15490 35308
rect 15170 33740 15490 35252
rect 15170 33684 15198 33740
rect 15254 33684 15302 33740
rect 15358 33684 15406 33740
rect 15462 33684 15490 33740
rect 15170 32172 15490 33684
rect 15170 32116 15198 32172
rect 15254 32116 15302 32172
rect 15358 32116 15406 32172
rect 15462 32116 15490 32172
rect 19832 36092 20152 36908
rect 19832 36036 19860 36092
rect 19916 36036 19964 36092
rect 20020 36036 20068 36092
rect 20124 36036 20152 36092
rect 19832 34524 20152 36036
rect 19832 34468 19860 34524
rect 19916 34468 19964 34524
rect 20020 34468 20068 34524
rect 20124 34468 20152 34524
rect 19832 32956 20152 34468
rect 19832 32900 19860 32956
rect 19916 32900 19964 32956
rect 20020 32900 20068 32956
rect 20124 32900 20152 32956
rect 10508 31332 10536 31388
rect 10592 31332 10640 31388
rect 10696 31332 10744 31388
rect 10800 31332 10828 31388
rect 10508 29820 10828 31332
rect 15036 31892 15092 31902
rect 15036 30660 15092 31836
rect 15036 30594 15092 30604
rect 15170 30604 15490 32116
rect 10508 29764 10536 29820
rect 10592 29764 10640 29820
rect 10696 29764 10744 29820
rect 10800 29764 10828 29820
rect 10508 28252 10828 29764
rect 12236 30548 12292 30558
rect 12236 29540 12292 30492
rect 12236 29474 12292 29484
rect 15170 30548 15198 30604
rect 15254 30548 15302 30604
rect 15358 30548 15406 30604
rect 15462 30548 15490 30604
rect 10508 28196 10536 28252
rect 10592 28196 10640 28252
rect 10696 28196 10744 28252
rect 10800 28196 10828 28252
rect 10508 26684 10828 28196
rect 10892 29092 10948 29102
rect 10892 26852 10948 29036
rect 10892 26786 10948 26796
rect 15170 29036 15490 30548
rect 15596 32116 15652 32126
rect 15596 29876 15652 32060
rect 15596 29810 15652 29820
rect 19832 31388 20152 32900
rect 24494 36876 24814 36908
rect 24494 36820 24522 36876
rect 24578 36820 24626 36876
rect 24682 36820 24730 36876
rect 24786 36820 24814 36876
rect 24494 35308 24814 36820
rect 29156 36092 29476 36908
rect 29156 36036 29184 36092
rect 29240 36036 29288 36092
rect 29344 36036 29392 36092
rect 29448 36036 29476 36092
rect 24494 35252 24522 35308
rect 24578 35252 24626 35308
rect 24682 35252 24730 35308
rect 24786 35252 24814 35308
rect 24494 33740 24814 35252
rect 26908 35364 26964 35374
rect 26908 35028 26964 35308
rect 26908 34962 26964 34972
rect 24494 33684 24522 33740
rect 24578 33684 24626 33740
rect 24682 33684 24730 33740
rect 24786 33684 24814 33740
rect 19832 31332 19860 31388
rect 19916 31332 19964 31388
rect 20020 31332 20068 31388
rect 20124 31332 20152 31388
rect 19832 29820 20152 31332
rect 19832 29764 19860 29820
rect 19916 29764 19964 29820
rect 20020 29764 20068 29820
rect 20124 29764 20152 29820
rect 15170 28980 15198 29036
rect 15254 28980 15302 29036
rect 15358 28980 15406 29036
rect 15462 28980 15490 29036
rect 15170 27468 15490 28980
rect 19628 29316 19684 29326
rect 19404 28084 19460 28094
rect 15170 27412 15198 27468
rect 15254 27412 15302 27468
rect 15358 27412 15406 27468
rect 15462 27412 15490 27468
rect 10508 26628 10536 26684
rect 10592 26628 10640 26684
rect 10696 26628 10744 26684
rect 10800 26628 10828 26684
rect 10508 25116 10828 26628
rect 10508 25060 10536 25116
rect 10592 25060 10640 25116
rect 10696 25060 10744 25116
rect 10800 25060 10828 25116
rect 10508 23548 10828 25060
rect 10508 23492 10536 23548
rect 10592 23492 10640 23548
rect 10696 23492 10744 23548
rect 10800 23492 10828 23548
rect 10508 21980 10828 23492
rect 10508 21924 10536 21980
rect 10592 21924 10640 21980
rect 10696 21924 10744 21980
rect 10800 21924 10828 21980
rect 10508 20412 10828 21924
rect 10508 20356 10536 20412
rect 10592 20356 10640 20412
rect 10696 20356 10744 20412
rect 10800 20356 10828 20412
rect 10508 18844 10828 20356
rect 10508 18788 10536 18844
rect 10592 18788 10640 18844
rect 10696 18788 10744 18844
rect 10800 18788 10828 18844
rect 10508 17276 10828 18788
rect 10508 17220 10536 17276
rect 10592 17220 10640 17276
rect 10696 17220 10744 17276
rect 10800 17220 10828 17276
rect 10508 15708 10828 17220
rect 10508 15652 10536 15708
rect 10592 15652 10640 15708
rect 10696 15652 10744 15708
rect 10800 15652 10828 15708
rect 10508 14140 10828 15652
rect 10508 14084 10536 14140
rect 10592 14084 10640 14140
rect 10696 14084 10744 14140
rect 10800 14084 10828 14140
rect 10508 12572 10828 14084
rect 10508 12516 10536 12572
rect 10592 12516 10640 12572
rect 10696 12516 10744 12572
rect 10800 12516 10828 12572
rect 10508 11004 10828 12516
rect 10508 10948 10536 11004
rect 10592 10948 10640 11004
rect 10696 10948 10744 11004
rect 10800 10948 10828 11004
rect 10508 9436 10828 10948
rect 10508 9380 10536 9436
rect 10592 9380 10640 9436
rect 10696 9380 10744 9436
rect 10800 9380 10828 9436
rect 10508 7868 10828 9380
rect 10508 7812 10536 7868
rect 10592 7812 10640 7868
rect 10696 7812 10744 7868
rect 10800 7812 10828 7868
rect 10508 6300 10828 7812
rect 10508 6244 10536 6300
rect 10592 6244 10640 6300
rect 10696 6244 10744 6300
rect 10800 6244 10828 6300
rect 10508 4732 10828 6244
rect 10508 4676 10536 4732
rect 10592 4676 10640 4732
rect 10696 4676 10744 4732
rect 10800 4676 10828 4732
rect 10508 3164 10828 4676
rect 10508 3108 10536 3164
rect 10592 3108 10640 3164
rect 10696 3108 10744 3164
rect 10800 3108 10828 3164
rect 10508 3076 10828 3108
rect 15170 25900 15490 27412
rect 15170 25844 15198 25900
rect 15254 25844 15302 25900
rect 15358 25844 15406 25900
rect 15462 25844 15490 25900
rect 15170 24332 15490 25844
rect 15170 24276 15198 24332
rect 15254 24276 15302 24332
rect 15358 24276 15406 24332
rect 15462 24276 15490 24332
rect 18956 27636 19012 27646
rect 15170 22764 15490 24276
rect 18172 24276 18228 24286
rect 18172 23604 18228 24220
rect 18956 23828 19012 27580
rect 19404 27076 19460 28028
rect 19404 25844 19460 27020
rect 19628 26628 19684 29260
rect 19628 26562 19684 26572
rect 19832 28252 20152 29764
rect 19832 28196 19860 28252
rect 19916 28196 19964 28252
rect 20020 28196 20068 28252
rect 20124 28196 20152 28252
rect 19832 26684 20152 28196
rect 21756 32788 21812 32798
rect 21756 28084 21812 32732
rect 24494 32172 24814 33684
rect 24494 32116 24522 32172
rect 24578 32116 24626 32172
rect 24682 32116 24730 32172
rect 24786 32116 24814 32172
rect 21756 28018 21812 28028
rect 24108 32004 24164 32014
rect 19832 26628 19860 26684
rect 19916 26628 19964 26684
rect 20020 26628 20068 26684
rect 20124 26628 20152 26684
rect 19404 25778 19460 25788
rect 18956 23762 19012 23772
rect 19832 25116 20152 26628
rect 19832 25060 19860 25116
rect 19916 25060 19964 25116
rect 20020 25060 20068 25116
rect 20124 25060 20152 25116
rect 18172 23538 18228 23548
rect 19832 23548 20152 25060
rect 20300 26628 20356 26638
rect 20300 25620 20356 26572
rect 20300 24724 20356 25564
rect 20300 24658 20356 24668
rect 24108 24948 24164 31948
rect 24108 24276 24164 24892
rect 24108 24210 24164 24220
rect 24494 30604 24814 32116
rect 29156 34524 29476 36036
rect 29156 34468 29184 34524
rect 29240 34468 29288 34524
rect 29344 34468 29392 34524
rect 29448 34468 29476 34524
rect 29156 32956 29476 34468
rect 29156 32900 29184 32956
rect 29240 32900 29288 32956
rect 29344 32900 29392 32956
rect 29448 32900 29476 32956
rect 33818 36876 34138 36908
rect 33818 36820 33846 36876
rect 33902 36820 33950 36876
rect 34006 36820 34054 36876
rect 34110 36820 34138 36876
rect 33818 35308 34138 36820
rect 33818 35252 33846 35308
rect 33902 35252 33950 35308
rect 34006 35252 34054 35308
rect 34110 35252 34138 35308
rect 33818 33740 34138 35252
rect 38480 36092 38800 36908
rect 38480 36036 38508 36092
rect 38564 36036 38612 36092
rect 38668 36036 38716 36092
rect 38772 36036 38800 36092
rect 35644 35028 35700 35038
rect 33818 33684 33846 33740
rect 33902 33684 33950 33740
rect 34006 33684 34054 33740
rect 34110 33684 34138 33740
rect 29156 31388 29476 32900
rect 29156 31332 29184 31388
rect 29240 31332 29288 31388
rect 29344 31332 29392 31388
rect 29448 31332 29476 31388
rect 26684 30996 26740 31006
rect 26684 30772 26740 30940
rect 26684 30706 26740 30716
rect 24494 30548 24522 30604
rect 24578 30548 24626 30604
rect 24682 30548 24730 30604
rect 24786 30548 24814 30604
rect 24494 29036 24814 30548
rect 24494 28980 24522 29036
rect 24578 28980 24626 29036
rect 24682 28980 24730 29036
rect 24786 28980 24814 29036
rect 24494 27468 24814 28980
rect 24494 27412 24522 27468
rect 24578 27412 24626 27468
rect 24682 27412 24730 27468
rect 24786 27412 24814 27468
rect 24494 25900 24814 27412
rect 24494 25844 24522 25900
rect 24578 25844 24626 25900
rect 24682 25844 24730 25900
rect 24786 25844 24814 25900
rect 24494 24332 24814 25844
rect 24494 24276 24522 24332
rect 24578 24276 24626 24332
rect 24682 24276 24730 24332
rect 24786 24276 24814 24332
rect 15170 22708 15198 22764
rect 15254 22708 15302 22764
rect 15358 22708 15406 22764
rect 15462 22708 15490 22764
rect 15170 21196 15490 22708
rect 15170 21140 15198 21196
rect 15254 21140 15302 21196
rect 15358 21140 15406 21196
rect 15462 21140 15490 21196
rect 15170 19628 15490 21140
rect 15170 19572 15198 19628
rect 15254 19572 15302 19628
rect 15358 19572 15406 19628
rect 15462 19572 15490 19628
rect 15170 18060 15490 19572
rect 15170 18004 15198 18060
rect 15254 18004 15302 18060
rect 15358 18004 15406 18060
rect 15462 18004 15490 18060
rect 15170 16492 15490 18004
rect 15170 16436 15198 16492
rect 15254 16436 15302 16492
rect 15358 16436 15406 16492
rect 15462 16436 15490 16492
rect 15170 14924 15490 16436
rect 15170 14868 15198 14924
rect 15254 14868 15302 14924
rect 15358 14868 15406 14924
rect 15462 14868 15490 14924
rect 15170 13356 15490 14868
rect 15170 13300 15198 13356
rect 15254 13300 15302 13356
rect 15358 13300 15406 13356
rect 15462 13300 15490 13356
rect 15170 11788 15490 13300
rect 15170 11732 15198 11788
rect 15254 11732 15302 11788
rect 15358 11732 15406 11788
rect 15462 11732 15490 11788
rect 15170 10220 15490 11732
rect 15170 10164 15198 10220
rect 15254 10164 15302 10220
rect 15358 10164 15406 10220
rect 15462 10164 15490 10220
rect 15170 8652 15490 10164
rect 15170 8596 15198 8652
rect 15254 8596 15302 8652
rect 15358 8596 15406 8652
rect 15462 8596 15490 8652
rect 15170 7084 15490 8596
rect 15170 7028 15198 7084
rect 15254 7028 15302 7084
rect 15358 7028 15406 7084
rect 15462 7028 15490 7084
rect 15170 5516 15490 7028
rect 15170 5460 15198 5516
rect 15254 5460 15302 5516
rect 15358 5460 15406 5516
rect 15462 5460 15490 5516
rect 15170 3948 15490 5460
rect 15170 3892 15198 3948
rect 15254 3892 15302 3948
rect 15358 3892 15406 3948
rect 15462 3892 15490 3948
rect 15170 3076 15490 3892
rect 19832 23492 19860 23548
rect 19916 23492 19964 23548
rect 20020 23492 20068 23548
rect 20124 23492 20152 23548
rect 19832 21980 20152 23492
rect 19832 21924 19860 21980
rect 19916 21924 19964 21980
rect 20020 21924 20068 21980
rect 20124 21924 20152 21980
rect 19832 20412 20152 21924
rect 19832 20356 19860 20412
rect 19916 20356 19964 20412
rect 20020 20356 20068 20412
rect 20124 20356 20152 20412
rect 19832 18844 20152 20356
rect 19832 18788 19860 18844
rect 19916 18788 19964 18844
rect 20020 18788 20068 18844
rect 20124 18788 20152 18844
rect 19832 17276 20152 18788
rect 19832 17220 19860 17276
rect 19916 17220 19964 17276
rect 20020 17220 20068 17276
rect 20124 17220 20152 17276
rect 19832 15708 20152 17220
rect 19832 15652 19860 15708
rect 19916 15652 19964 15708
rect 20020 15652 20068 15708
rect 20124 15652 20152 15708
rect 19832 14140 20152 15652
rect 19832 14084 19860 14140
rect 19916 14084 19964 14140
rect 20020 14084 20068 14140
rect 20124 14084 20152 14140
rect 19832 12572 20152 14084
rect 19832 12516 19860 12572
rect 19916 12516 19964 12572
rect 20020 12516 20068 12572
rect 20124 12516 20152 12572
rect 19832 11004 20152 12516
rect 19832 10948 19860 11004
rect 19916 10948 19964 11004
rect 20020 10948 20068 11004
rect 20124 10948 20152 11004
rect 19832 9436 20152 10948
rect 19832 9380 19860 9436
rect 19916 9380 19964 9436
rect 20020 9380 20068 9436
rect 20124 9380 20152 9436
rect 19832 7868 20152 9380
rect 19832 7812 19860 7868
rect 19916 7812 19964 7868
rect 20020 7812 20068 7868
rect 20124 7812 20152 7868
rect 19832 6300 20152 7812
rect 19832 6244 19860 6300
rect 19916 6244 19964 6300
rect 20020 6244 20068 6300
rect 20124 6244 20152 6300
rect 19832 4732 20152 6244
rect 19832 4676 19860 4732
rect 19916 4676 19964 4732
rect 20020 4676 20068 4732
rect 20124 4676 20152 4732
rect 19832 3164 20152 4676
rect 19832 3108 19860 3164
rect 19916 3108 19964 3164
rect 20020 3108 20068 3164
rect 20124 3108 20152 3164
rect 19832 3076 20152 3108
rect 24494 22764 24814 24276
rect 24494 22708 24522 22764
rect 24578 22708 24626 22764
rect 24682 22708 24730 22764
rect 24786 22708 24814 22764
rect 24494 21196 24814 22708
rect 24494 21140 24522 21196
rect 24578 21140 24626 21196
rect 24682 21140 24730 21196
rect 24786 21140 24814 21196
rect 24494 19628 24814 21140
rect 24494 19572 24522 19628
rect 24578 19572 24626 19628
rect 24682 19572 24730 19628
rect 24786 19572 24814 19628
rect 24494 18060 24814 19572
rect 24494 18004 24522 18060
rect 24578 18004 24626 18060
rect 24682 18004 24730 18060
rect 24786 18004 24814 18060
rect 24494 16492 24814 18004
rect 29156 29820 29476 31332
rect 31724 32900 31780 32910
rect 29156 29764 29184 29820
rect 29240 29764 29288 29820
rect 29344 29764 29392 29820
rect 29448 29764 29476 29820
rect 29156 28252 29476 29764
rect 29156 28196 29184 28252
rect 29240 28196 29288 28252
rect 29344 28196 29392 28252
rect 29448 28196 29476 28252
rect 29156 26684 29476 28196
rect 29596 30212 29652 30222
rect 29596 29540 29652 30156
rect 29596 28868 29652 29484
rect 29596 27860 29652 28812
rect 29596 27794 29652 27804
rect 30940 29652 30996 29662
rect 30940 27636 30996 29596
rect 31612 29204 31668 29214
rect 31612 27860 31668 29148
rect 31612 27794 31668 27804
rect 30940 27570 30996 27580
rect 29156 26628 29184 26684
rect 29240 26628 29288 26684
rect 29344 26628 29392 26684
rect 29448 26628 29476 26684
rect 29156 25116 29476 26628
rect 29156 25060 29184 25116
rect 29240 25060 29288 25116
rect 29344 25060 29392 25116
rect 29448 25060 29476 25116
rect 29156 23548 29476 25060
rect 31724 24388 31780 32844
rect 31724 24322 31780 24332
rect 33818 32172 34138 33684
rect 33818 32116 33846 32172
rect 33902 32116 33950 32172
rect 34006 32116 34054 32172
rect 34110 32116 34138 32172
rect 33818 30604 34138 32116
rect 33818 30548 33846 30604
rect 33902 30548 33950 30604
rect 34006 30548 34054 30604
rect 34110 30548 34138 30604
rect 33818 29036 34138 30548
rect 33818 28980 33846 29036
rect 33902 28980 33950 29036
rect 34006 28980 34054 29036
rect 34110 28980 34138 29036
rect 33818 27468 34138 28980
rect 33818 27412 33846 27468
rect 33902 27412 33950 27468
rect 34006 27412 34054 27468
rect 34110 27412 34138 27468
rect 33818 25900 34138 27412
rect 33818 25844 33846 25900
rect 33902 25844 33950 25900
rect 34006 25844 34054 25900
rect 34110 25844 34138 25900
rect 33818 24332 34138 25844
rect 29156 23492 29184 23548
rect 29240 23492 29288 23548
rect 29344 23492 29392 23548
rect 29448 23492 29476 23548
rect 29156 21980 29476 23492
rect 29156 21924 29184 21980
rect 29240 21924 29288 21980
rect 29344 21924 29392 21980
rect 29448 21924 29476 21980
rect 29156 20412 29476 21924
rect 29156 20356 29184 20412
rect 29240 20356 29288 20412
rect 29344 20356 29392 20412
rect 29448 20356 29476 20412
rect 29156 18844 29476 20356
rect 29156 18788 29184 18844
rect 29240 18788 29288 18844
rect 29344 18788 29392 18844
rect 29448 18788 29476 18844
rect 29156 17276 29476 18788
rect 24494 16436 24522 16492
rect 24578 16436 24626 16492
rect 24682 16436 24730 16492
rect 24786 16436 24814 16492
rect 24494 14924 24814 16436
rect 25452 17220 25508 17230
rect 25452 16100 25508 17164
rect 25452 16034 25508 16044
rect 29156 17220 29184 17276
rect 29240 17220 29288 17276
rect 29344 17220 29392 17276
rect 29448 17220 29476 17276
rect 24494 14868 24522 14924
rect 24578 14868 24626 14924
rect 24682 14868 24730 14924
rect 24786 14868 24814 14924
rect 24494 13356 24814 14868
rect 24494 13300 24522 13356
rect 24578 13300 24626 13356
rect 24682 13300 24730 13356
rect 24786 13300 24814 13356
rect 24494 11788 24814 13300
rect 24494 11732 24522 11788
rect 24578 11732 24626 11788
rect 24682 11732 24730 11788
rect 24786 11732 24814 11788
rect 24494 10220 24814 11732
rect 24494 10164 24522 10220
rect 24578 10164 24626 10220
rect 24682 10164 24730 10220
rect 24786 10164 24814 10220
rect 24494 8652 24814 10164
rect 24494 8596 24522 8652
rect 24578 8596 24626 8652
rect 24682 8596 24730 8652
rect 24786 8596 24814 8652
rect 24494 7084 24814 8596
rect 24494 7028 24522 7084
rect 24578 7028 24626 7084
rect 24682 7028 24730 7084
rect 24786 7028 24814 7084
rect 24494 5516 24814 7028
rect 24494 5460 24522 5516
rect 24578 5460 24626 5516
rect 24682 5460 24730 5516
rect 24786 5460 24814 5516
rect 24494 3948 24814 5460
rect 24494 3892 24522 3948
rect 24578 3892 24626 3948
rect 24682 3892 24730 3948
rect 24786 3892 24814 3948
rect 24494 3076 24814 3892
rect 29156 15708 29476 17220
rect 29156 15652 29184 15708
rect 29240 15652 29288 15708
rect 29344 15652 29392 15708
rect 29448 15652 29476 15708
rect 29156 14140 29476 15652
rect 29156 14084 29184 14140
rect 29240 14084 29288 14140
rect 29344 14084 29392 14140
rect 29448 14084 29476 14140
rect 29156 12572 29476 14084
rect 33818 24276 33846 24332
rect 33902 24276 33950 24332
rect 34006 24276 34054 24332
rect 34110 24276 34138 24332
rect 33818 22764 34138 24276
rect 33818 22708 33846 22764
rect 33902 22708 33950 22764
rect 34006 22708 34054 22764
rect 34110 22708 34138 22764
rect 33818 21196 34138 22708
rect 33818 21140 33846 21196
rect 33902 21140 33950 21196
rect 34006 21140 34054 21196
rect 34110 21140 34138 21196
rect 33818 19628 34138 21140
rect 35308 34804 35364 34814
rect 35308 20244 35364 34748
rect 35420 34468 35476 34478
rect 35420 31780 35476 34412
rect 35644 33908 35700 34972
rect 35644 33012 35700 33852
rect 35644 32946 35700 32956
rect 38480 34524 38800 36036
rect 38480 34468 38508 34524
rect 38564 34468 38612 34524
rect 38668 34468 38716 34524
rect 38772 34468 38800 34524
rect 38480 32956 38800 34468
rect 35420 31714 35476 31724
rect 38480 32900 38508 32956
rect 38564 32900 38612 32956
rect 38668 32900 38716 32956
rect 38772 32900 38800 32956
rect 37100 31444 37156 31454
rect 37100 29652 37156 31388
rect 38480 31388 38800 32900
rect 38480 31332 38508 31388
rect 38564 31332 38612 31388
rect 38668 31332 38716 31388
rect 38772 31332 38800 31388
rect 37100 29586 37156 29596
rect 37660 31108 37716 31118
rect 37660 28420 37716 31052
rect 37660 28354 37716 28364
rect 38480 29820 38800 31332
rect 38480 29764 38508 29820
rect 38564 29764 38612 29820
rect 38668 29764 38716 29820
rect 38772 29764 38800 29820
rect 38480 28252 38800 29764
rect 38480 28196 38508 28252
rect 38564 28196 38612 28252
rect 38668 28196 38716 28252
rect 38772 28196 38800 28252
rect 38480 26684 38800 28196
rect 38480 26628 38508 26684
rect 38564 26628 38612 26684
rect 38668 26628 38716 26684
rect 38772 26628 38800 26684
rect 35420 25508 35476 25518
rect 35420 24052 35476 25452
rect 35420 23986 35476 23996
rect 35644 25396 35700 25406
rect 35644 24052 35700 25340
rect 35644 23986 35700 23996
rect 38480 25116 38800 26628
rect 38480 25060 38508 25116
rect 38564 25060 38612 25116
rect 38668 25060 38716 25116
rect 38772 25060 38800 25116
rect 35308 20178 35364 20188
rect 38480 23548 38800 25060
rect 38480 23492 38508 23548
rect 38564 23492 38612 23548
rect 38668 23492 38716 23548
rect 38772 23492 38800 23548
rect 38480 21980 38800 23492
rect 38480 21924 38508 21980
rect 38564 21924 38612 21980
rect 38668 21924 38716 21980
rect 38772 21924 38800 21980
rect 38480 20412 38800 21924
rect 38480 20356 38508 20412
rect 38564 20356 38612 20412
rect 38668 20356 38716 20412
rect 38772 20356 38800 20412
rect 33818 19572 33846 19628
rect 33902 19572 33950 19628
rect 34006 19572 34054 19628
rect 34110 19572 34138 19628
rect 33818 18060 34138 19572
rect 33818 18004 33846 18060
rect 33902 18004 33950 18060
rect 34006 18004 34054 18060
rect 34110 18004 34138 18060
rect 33818 16492 34138 18004
rect 33818 16436 33846 16492
rect 33902 16436 33950 16492
rect 34006 16436 34054 16492
rect 34110 16436 34138 16492
rect 33818 14924 34138 16436
rect 38480 18844 38800 20356
rect 38480 18788 38508 18844
rect 38564 18788 38612 18844
rect 38668 18788 38716 18844
rect 38772 18788 38800 18844
rect 38480 17276 38800 18788
rect 38480 17220 38508 17276
rect 38564 17220 38612 17276
rect 38668 17220 38716 17276
rect 38772 17220 38800 17276
rect 38480 15708 38800 17220
rect 38480 15652 38508 15708
rect 38564 15652 38612 15708
rect 38668 15652 38716 15708
rect 38772 15652 38800 15708
rect 33818 14868 33846 14924
rect 33902 14868 33950 14924
rect 34006 14868 34054 14924
rect 34110 14868 34138 14924
rect 31612 13748 31668 13758
rect 31612 12740 31668 13692
rect 31612 12674 31668 12684
rect 33628 13636 33684 13646
rect 33628 12740 33684 13580
rect 33628 12674 33684 12684
rect 33818 13356 34138 14868
rect 33818 13300 33846 13356
rect 33902 13300 33950 13356
rect 34006 13300 34054 13356
rect 34110 13300 34138 13356
rect 29156 12516 29184 12572
rect 29240 12516 29288 12572
rect 29344 12516 29392 12572
rect 29448 12516 29476 12572
rect 29156 11004 29476 12516
rect 29156 10948 29184 11004
rect 29240 10948 29288 11004
rect 29344 10948 29392 11004
rect 29448 10948 29476 11004
rect 29156 9436 29476 10948
rect 29156 9380 29184 9436
rect 29240 9380 29288 9436
rect 29344 9380 29392 9436
rect 29448 9380 29476 9436
rect 29156 7868 29476 9380
rect 29156 7812 29184 7868
rect 29240 7812 29288 7868
rect 29344 7812 29392 7868
rect 29448 7812 29476 7868
rect 29156 6300 29476 7812
rect 29156 6244 29184 6300
rect 29240 6244 29288 6300
rect 29344 6244 29392 6300
rect 29448 6244 29476 6300
rect 29156 4732 29476 6244
rect 29156 4676 29184 4732
rect 29240 4676 29288 4732
rect 29344 4676 29392 4732
rect 29448 4676 29476 4732
rect 29156 3164 29476 4676
rect 29156 3108 29184 3164
rect 29240 3108 29288 3164
rect 29344 3108 29392 3164
rect 29448 3108 29476 3164
rect 29156 3076 29476 3108
rect 33818 11788 34138 13300
rect 34300 15092 34356 15102
rect 34300 12852 34356 15036
rect 34300 12786 34356 12796
rect 38480 14140 38800 15652
rect 38480 14084 38508 14140
rect 38564 14084 38612 14140
rect 38668 14084 38716 14140
rect 38772 14084 38800 14140
rect 33818 11732 33846 11788
rect 33902 11732 33950 11788
rect 34006 11732 34054 11788
rect 34110 11732 34138 11788
rect 33818 10220 34138 11732
rect 33818 10164 33846 10220
rect 33902 10164 33950 10220
rect 34006 10164 34054 10220
rect 34110 10164 34138 10220
rect 33818 8652 34138 10164
rect 33818 8596 33846 8652
rect 33902 8596 33950 8652
rect 34006 8596 34054 8652
rect 34110 8596 34138 8652
rect 33818 7084 34138 8596
rect 33818 7028 33846 7084
rect 33902 7028 33950 7084
rect 34006 7028 34054 7084
rect 34110 7028 34138 7084
rect 33818 5516 34138 7028
rect 33818 5460 33846 5516
rect 33902 5460 33950 5516
rect 34006 5460 34054 5516
rect 34110 5460 34138 5516
rect 33818 3948 34138 5460
rect 33818 3892 33846 3948
rect 33902 3892 33950 3948
rect 34006 3892 34054 3948
rect 34110 3892 34138 3948
rect 33818 3076 34138 3892
rect 38480 12572 38800 14084
rect 38480 12516 38508 12572
rect 38564 12516 38612 12572
rect 38668 12516 38716 12572
rect 38772 12516 38800 12572
rect 38480 11004 38800 12516
rect 38480 10948 38508 11004
rect 38564 10948 38612 11004
rect 38668 10948 38716 11004
rect 38772 10948 38800 11004
rect 38480 9436 38800 10948
rect 38480 9380 38508 9436
rect 38564 9380 38612 9436
rect 38668 9380 38716 9436
rect 38772 9380 38800 9436
rect 38480 7868 38800 9380
rect 38480 7812 38508 7868
rect 38564 7812 38612 7868
rect 38668 7812 38716 7868
rect 38772 7812 38800 7868
rect 38480 6300 38800 7812
rect 38480 6244 38508 6300
rect 38564 6244 38612 6300
rect 38668 6244 38716 6300
rect 38772 6244 38800 6300
rect 38480 4732 38800 6244
rect 38480 4676 38508 4732
rect 38564 4676 38612 4732
rect 38668 4676 38716 4732
rect 38772 4676 38800 4732
rect 38480 3164 38800 4676
rect 38480 3108 38508 3164
rect 38564 3108 38612 3164
rect 38668 3108 38716 3164
rect 38772 3108 38800 3164
rect 38480 3076 38800 3108
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0562_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751534193
transform 1 0 22960 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _0563_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752061876
transform 1 0 19152 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_8  _0564_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752063767
transform 1 0 18144 0 -1 14112
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0565_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751889408
transform 1 0 20048 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0566_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753182340
transform 1 0 19712 0 1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0567_
timestamp 1751534193
transform 1 0 29120 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0568_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751740063
transform -1 0 23520 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0569_
timestamp 1753182340
transform 1 0 22512 0 1 14112
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0570_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753441877
transform -1 0 21616 0 -1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0571_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752063729
transform 1 0 21392 0 -1 20384
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0572_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751914308
transform 1 0 21168 0 1 15680
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0573_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532043
transform 1 0 31136 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0574_
timestamp 1751889408
transform 1 0 29008 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0575_
timestamp 1751889408
transform 1 0 31360 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0576_
timestamp 1751534193
transform -1 0 31360 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0577_
timestamp 1751534193
transform -1 0 23184 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0578_
timestamp 1751534193
transform 1 0 21616 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0579_
timestamp 1751532043
transform -1 0 20160 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0580_
timestamp 1751534193
transform 1 0 23408 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0581_
timestamp 1751534193
transform 1 0 24080 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0582_
timestamp 1751534193
transform 1 0 18032 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0583_
timestamp 1751534193
transform -1 0 20832 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0584_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753868718
transform 1 0 21840 0 -1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0585_
timestamp 1751889408
transform 1 0 23744 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0586_
timestamp 1751914308
transform 1 0 21616 0 -1 15680
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0587_
timestamp 1751889408
transform -1 0 23968 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0588_
timestamp 1751914308
transform 1 0 21168 0 1 14112
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0589_
timestamp 1751889408
transform 1 0 24080 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0590_
timestamp 1751534193
transform -1 0 28112 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0591_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752345181
transform 1 0 24528 0 1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0592_
timestamp 1751740063
transform 1 0 25088 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0593_
timestamp 1751534193
transform -1 0 19488 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0594_
timestamp 1751534193
transform -1 0 17024 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0595_
timestamp 1751534193
transform 1 0 14336 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0596_
timestamp 1751534193
transform 1 0 28112 0 1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0597_
timestamp 1751534193
transform -1 0 37968 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0598_
timestamp 1751532043
transform -1 0 29680 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0599_
timestamp 1752063729
transform -1 0 38304 0 -1 29792
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0600_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751889808
transform -1 0 35280 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0601_
timestamp 1751740063
transform -1 0 29792 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0602_
timestamp 1751889408
transform 1 0 23184 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0603_
timestamp 1751532043
transform -1 0 22064 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0604_
timestamp 1751532043
transform -1 0 21616 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0605_
timestamp 1753868718
transform 1 0 20160 0 -1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0606_
timestamp 1751534193
transform 1 0 26096 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0607_
timestamp 1751532043
transform 1 0 25312 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0608_
timestamp 1753182340
transform 1 0 25760 0 1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0609_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753172561
transform -1 0 28336 0 -1 23520
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0610_
timestamp 1751534193
transform 1 0 30464 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0611_
timestamp 1753182340
transform 1 0 33376 0 1 25088
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0612_
timestamp 1751914308
transform 1 0 31360 0 -1 28224
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0613_
timestamp 1751889408
transform -1 0 36512 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0614_
timestamp 1752063729
transform -1 0 35280 0 -1 32928
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0615_
timestamp 1751534193
transform 1 0 29232 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0616_
timestamp 1751534193
transform 1 0 29792 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0617_
timestamp 1751534193
transform 1 0 33376 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0618_
timestamp 1751889408
transform -1 0 33936 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0619_
timestamp 1751534193
transform -1 0 35840 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0620_
timestamp 1751534193
transform 1 0 34496 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0621_
timestamp 1752063729
transform -1 0 37296 0 -1 25088
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0622_
timestamp 1751534193
transform -1 0 31920 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0623_
timestamp 1751534193
transform -1 0 32592 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0624_
timestamp 1751740063
transform 1 0 31136 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0625_
timestamp 1753172561
transform 1 0 31696 0 1 21952
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0626_
timestamp 1751914308
transform 1 0 33264 0 1 21952
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0627_
timestamp 1752063729
transform 1 0 33936 0 -1 21952
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0628_
timestamp 1751889408
transform 1 0 34608 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0629_
timestamp 1751534193
transform -1 0 19712 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0630_
timestamp 1751534193
transform 1 0 19040 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _0631_
timestamp 1752061876
transform 1 0 30352 0 -1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0632_
timestamp 1751534193
transform 1 0 31920 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0633_
timestamp 1752345181
transform 1 0 31472 0 -1 21952
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0634_
timestamp 1751914308
transform 1 0 33152 0 -1 20384
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0635_
timestamp 1752063729
transform 1 0 35952 0 -1 21952
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0636_
timestamp 1751534193
transform -1 0 30912 0 1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0637_
timestamp 1751889408
transform 1 0 30464 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _0638_
timestamp 1752061876
transform 1 0 31472 0 -1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0639_
timestamp 1752345181
transform -1 0 32144 0 1 26656
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0640_
timestamp 1751889808
transform -1 0 30912 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0641_
timestamp 1751914308
transform 1 0 31248 0 1 28224
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0642_
timestamp 1751534193
transform -1 0 30464 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0643_
timestamp 1751889408
transform 1 0 32816 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0644_
timestamp 1752345181
transform -1 0 33376 0 1 25088
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0645_
timestamp 1751914308
transform 1 0 32928 0 -1 28224
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0646_
timestamp 1752063729
transform 1 0 33600 0 -1 26656
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0647_
timestamp 1753182340
transform -1 0 32144 0 1 25088
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0648_
timestamp 1751914308
transform -1 0 34272 0 -1 31360
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0649_
timestamp 1751889408
transform 1 0 31920 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0650_
timestamp 1751534193
transform 1 0 37296 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0651_
timestamp 1751534193
transform -1 0 14000 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0652_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751531619
transform -1 0 31248 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0653_
timestamp 1753182340
transform 1 0 29680 0 1 25088
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0654_
timestamp 1751914308
transform 1 0 29904 0 1 28224
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0655_
timestamp 1751889408
transform 1 0 30912 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0656_
timestamp 1751534193
transform 1 0 31696 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0657_
timestamp 1751889408
transform 1 0 29344 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0658_
timestamp 1752345181
transform 1 0 30912 0 -1 26656
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0659_
timestamp 1751889808
transform 1 0 32144 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0660_
timestamp 1751914308
transform 1 0 36848 0 1 29792
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0661_
timestamp 1751534193
transform -1 0 34720 0 1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0662_
timestamp 1751532043
transform -1 0 29456 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0663_
timestamp 1751534193
transform 1 0 27776 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0664_
timestamp 1751531619
transform 1 0 23744 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0665_
timestamp 1751889408
transform 1 0 26656 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0666_
timestamp 1751531619
transform -1 0 26096 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0667_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753960525
transform -1 0 26096 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0668_
timestamp 1751534193
transform -1 0 18256 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0669_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753371985
transform 1 0 19824 0 1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0670_
timestamp 1751889408
transform 1 0 23408 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0671_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753277515
transform -1 0 25648 0 1 15680
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0672_
timestamp 1751889408
transform -1 0 25424 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0673_
timestamp 1751534193
transform 1 0 25760 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0674_
timestamp 1751914308
transform -1 0 37520 0 -1 23520
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0675_
timestamp 1751532043
transform 1 0 35728 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0676_
timestamp 1753371985
transform -1 0 36400 0 1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0677_
timestamp 1753960525
transform 1 0 35504 0 1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0678_
timestamp 1751914308
transform 1 0 36848 0 1 32928
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0679_
timestamp 1751914308
transform 1 0 36848 0 1 20384
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0680_
timestamp 1751914308
transform -1 0 38192 0 1 26656
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0681_
timestamp 1751914308
transform 1 0 36848 0 1 31360
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0682_
timestamp 1751914308
transform 1 0 34720 0 1 32928
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0683_
timestamp 1751914308
transform 1 0 36848 0 1 28224
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0684_
timestamp 1751914308
transform -1 0 38192 0 1 25088
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0685_
timestamp 1751914308
transform -1 0 38192 0 1 23520
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _0686_
timestamp 1752061876
transform 1 0 18704 0 1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0687_
timestamp 1751740063
transform -1 0 22288 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0688_
timestamp 1753868718
transform 1 0 20272 0 -1 17248
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0689_
timestamp 1753960525
transform 1 0 25424 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0690_
timestamp 1753960525
transform -1 0 30016 0 -1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0691_
timestamp 1751531619
transform 1 0 28448 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0692_
timestamp 1753441877
transform 1 0 30576 0 1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0693_
timestamp 1753371985
transform 1 0 26096 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0694_
timestamp 1752345181
transform -1 0 28784 0 1 15680
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0695_
timestamp 1753277515
transform 1 0 21168 0 1 10976
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0696_
timestamp 1753277515
transform 1 0 21168 0 1 12544
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0697_
timestamp 1751532043
transform 1 0 22288 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0698_
timestamp 1751914308
transform 1 0 22176 0 -1 14112
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0699_
timestamp 1751532043
transform 1 0 23744 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _0700_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751905124
transform -1 0 31136 0 -1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _0701_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753891287
transform -1 0 30800 0 -1 17248
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0702_
timestamp 1753441877
transform 1 0 29680 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _0703_
timestamp 1753891287
transform -1 0 30576 0 1 15680
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0704_
timestamp 1751532043
transform -1 0 25536 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0705_
timestamp 1753172561
transform -1 0 23632 0 1 18816
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0706_
timestamp 1751534193
transform -1 0 11088 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0707_
timestamp 1751889408
transform 1 0 9856 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0708_
timestamp 1751740063
transform -1 0 35504 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0709_
timestamp 1751534193
transform -1 0 30576 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0710_
timestamp 1753172561
transform 1 0 25984 0 -1 21952
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0711_
timestamp 1751531619
transform -1 0 22960 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0712_
timestamp 1751534193
transform 1 0 14672 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0713_
timestamp 1753371985
transform -1 0 14448 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_4  _0714_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751546029
transform -1 0 10304 0 1 12544
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0715_
timestamp 1751914308
transform 1 0 11760 0 1 10976
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0716_
timestamp 1751889408
transform -1 0 14336 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0717_
timestamp 1752063729
transform 1 0 14336 0 -1 10976
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0718_
timestamp 1751534193
transform -1 0 14336 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0719_
timestamp 1751889408
transform 1 0 8400 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0720_
timestamp 1751914308
transform 1 0 9408 0 -1 10976
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0721_
timestamp 1751889408
transform -1 0 12096 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0722_
timestamp 1752063729
transform 1 0 10416 0 1 9408
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0723_
timestamp 1752345181
transform 1 0 25536 0 1 21952
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0724_
timestamp 1751531619
transform -1 0 29120 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_4  _0725_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751882821
transform 1 0 27104 0 1 21952
box -86 -86 1542 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0726_
timestamp 1752063729
transform -1 0 17024 0 -1 9408
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0727_
timestamp 1751914308
transform -1 0 14672 0 1 7840
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0728_
timestamp 1751889408
transform -1 0 14112 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0729_
timestamp 1752063729
transform 1 0 12768 0 -1 9408
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0730_
timestamp 1751914308
transform 1 0 9632 0 -1 6272
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0731_
timestamp 1751889408
transform -1 0 12208 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0732_
timestamp 1752063729
transform 1 0 11088 0 1 6272
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0733_
timestamp 1751914308
transform -1 0 14672 0 1 6272
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0734_
timestamp 1751889408
transform -1 0 13776 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0735_
timestamp 1752063729
transform -1 0 13104 0 1 4704
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0736_
timestamp 1751534193
transform 1 0 19712 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0737_
timestamp 1751534193
transform -1 0 21840 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0738_
timestamp 1751914308
transform 1 0 15680 0 -1 4704
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0739_
timestamp 1751889408
transform -1 0 18032 0 -1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0740_
timestamp 1752063729
transform -1 0 15456 0 1 4704
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0741_
timestamp 1752063729
transform -1 0 20160 0 1 9408
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0742_
timestamp 1751914308
transform -1 0 16464 0 1 6272
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0743_
timestamp 1751889408
transform -1 0 17024 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0744_
timestamp 1752063729
transform 1 0 16464 0 1 6272
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0745_
timestamp 1751914308
transform 1 0 18704 0 1 6272
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0746_
timestamp 1751889408
transform 1 0 20048 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0747_
timestamp 1752063729
transform -1 0 20720 0 -1 9408
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0748_
timestamp 1751914308
transform -1 0 21616 0 -1 7840
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0749_
timestamp 1751889408
transform 1 0 20160 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0750_
timestamp 1752063729
transform -1 0 20944 0 1 4704
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0751_
timestamp 1751534193
transform 1 0 22176 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0752_
timestamp 1751914308
transform 1 0 21280 0 -1 6272
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0753_
timestamp 1751889408
transform 1 0 22624 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0754_
timestamp 1752063729
transform -1 0 23744 0 1 4704
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _0755_
timestamp 1751905124
transform 1 0 30576 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0756_
timestamp 1751534193
transform -1 0 31024 0 -1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0757_
timestamp 1751889408
transform -1 0 27440 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0758_
timestamp 1753960525
transform -1 0 30912 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0759_
timestamp 1752345181
transform -1 0 31024 0 -1 21952
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_4  _0760_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752061857
transform 1 0 30240 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0761_
timestamp 1752063729
transform -1 0 32144 0 1 7840
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0762_
timestamp 1751914308
transform -1 0 26544 0 -1 7840
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0763_
timestamp 1751889408
transform -1 0 23632 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0764_
timestamp 1752063729
transform -1 0 24080 0 1 6272
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0765_
timestamp 1751914308
transform 1 0 26544 0 -1 7840
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0766_
timestamp 1751914308
transform -1 0 29232 0 -1 6272
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0767_
timestamp 1751889408
transform 1 0 24080 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0768_
timestamp 1752063729
transform 1 0 24640 0 1 6272
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0769_
timestamp 1751914308
transform -1 0 30576 0 -1 6272
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0770_
timestamp 1751914308
transform -1 0 29232 0 -1 7840
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0771_
timestamp 1751889408
transform 1 0 25984 0 -1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0772_
timestamp 1752063729
transform 1 0 26656 0 1 6272
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0773_
timestamp 1751534193
transform 1 0 29008 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0774_
timestamp 1751914308
transform 1 0 29344 0 1 6272
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0775_
timestamp 1751914308
transform 1 0 30576 0 -1 6272
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0776_
timestamp 1751889408
transform 1 0 30688 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0777_
timestamp 1752063729
transform -1 0 31920 0 -1 4704
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0778_
timestamp 1751534193
transform 1 0 32144 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0779_
timestamp 1751914308
transform -1 0 34272 0 -1 6272
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0780_
timestamp 1752063729
transform 1 0 30688 0 -1 9408
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0781_
timestamp 1751914308
transform 1 0 33152 0 1 6272
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0782_
timestamp 1751889408
transform 1 0 31920 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0783_
timestamp 1752063729
transform 1 0 32928 0 -1 4704
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0784_
timestamp 1751914308
transform 1 0 34944 0 -1 4704
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0785_
timestamp 1751914308
transform 1 0 36848 0 1 6272
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0786_
timestamp 1751889408
transform 1 0 34608 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0787_
timestamp 1752063729
transform 1 0 34608 0 1 6272
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0788_
timestamp 1751914308
transform 1 0 34160 0 -1 7840
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0789_
timestamp 1751914308
transform 1 0 36848 0 1 7840
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0790_
timestamp 1751889408
transform 1 0 34160 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0791_
timestamp 1752063729
transform 1 0 35504 0 -1 7840
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0792_
timestamp 1751534193
transform -1 0 28784 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0793_
timestamp 1751914308
transform 1 0 34944 0 1 7840
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0794_
timestamp 1751914308
transform 1 0 36848 0 1 9408
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0795_
timestamp 1751889408
transform 1 0 32592 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0796_
timestamp 1752063729
transform 1 0 33376 0 1 9408
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0797_
timestamp 1751740063
transform -1 0 30352 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0798_
timestamp 1751740063
transform 1 0 28784 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0799_
timestamp 1751531619
transform 1 0 28784 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0800_
timestamp 1751534193
transform -1 0 30128 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0801_
timestamp 1751889408
transform -1 0 26656 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0802_
timestamp 1751889408
transform 1 0 32032 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0803_
timestamp 1753172561
transform 1 0 29792 0 -1 20384
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0804_
timestamp 1753371985
transform 1 0 30912 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0805_
timestamp 1751534193
transform -1 0 32256 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0806_
timestamp 1751914308
transform -1 0 26992 0 1 9408
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0807_
timestamp 1751889408
transform -1 0 26656 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0808_
timestamp 1751534193
transform -1 0 23968 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0809_
timestamp 1751914308
transform -1 0 27104 0 -1 9408
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0810_
timestamp 1751914308
transform 1 0 26992 0 1 9408
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0811_
timestamp 1751889408
transform -1 0 27888 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0812_
timestamp 1751534193
transform -1 0 27328 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0813_
timestamp 1751914308
transform -1 0 29232 0 -1 9408
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0814_
timestamp 1751914308
transform -1 0 30576 0 -1 9408
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0815_
timestamp 1751889408
transform 1 0 29008 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0816_
timestamp 1751534193
transform 1 0 30128 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0817_
timestamp 1751534193
transform 1 0 14112 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0818_
timestamp 1751534193
transform 1 0 15344 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0819_
timestamp 1751914308
transform 1 0 29792 0 -1 10976
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0820_
timestamp 1751914308
transform 1 0 31024 0 -1 12544
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0821_
timestamp 1751889408
transform -1 0 31584 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0822_
timestamp 1751534193
transform -1 0 30016 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0823_
timestamp 1751534193
transform 1 0 31472 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0824_
timestamp 1751914308
transform 1 0 33040 0 1 12544
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0825_
timestamp 1751534193
transform 1 0 32816 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0826_
timestamp 1751914308
transform 1 0 33712 0 -1 15680
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0827_
timestamp 1751889408
transform -1 0 34832 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0828_
timestamp 1751534193
transform -1 0 34608 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0829_
timestamp 1751914308
transform 1 0 34496 0 1 12544
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0830_
timestamp 1751914308
transform 1 0 36848 0 1 12544
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0831_
timestamp 1751889408
transform 1 0 35840 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0832_
timestamp 1751534193
transform 1 0 37408 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0833_
timestamp 1751914308
transform -1 0 37408 0 -1 14112
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0834_
timestamp 1751914308
transform 1 0 35280 0 1 14112
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0835_
timestamp 1751889408
transform 1 0 36848 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0836_
timestamp 1751534193
transform -1 0 34496 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0837_
timestamp 1751534193
transform -1 0 9072 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0838_
timestamp 1751914308
transform -1 0 36400 0 -1 15680
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0839_
timestamp 1751914308
transform -1 0 36176 0 1 15680
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0840_
timestamp 1751889408
transform 1 0 33936 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0841_
timestamp 1751534193
transform 1 0 34720 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0842_
timestamp 1751532043
transform -1 0 24864 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0843_
timestamp 1751532043
transform -1 0 29344 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0844_
timestamp 1751534193
transform -1 0 25648 0 1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0845_
timestamp 1753441877
transform 1 0 26432 0 -1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0846_
timestamp 1751534193
transform -1 0 24864 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0847_
timestamp 1751534193
transform -1 0 28112 0 1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0848_
timestamp 1753441877
transform 1 0 24864 0 1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0849_
timestamp 1751534193
transform 1 0 27216 0 1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0850_
timestamp 1752345181
transform 1 0 19712 0 1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0851_
timestamp 1752063729
transform 1 0 10976 0 1 25088
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0852_
timestamp 1752063729
transform -1 0 15344 0 1 25088
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0853_
timestamp 1751534193
transform -1 0 15232 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0854_
timestamp 1751532043
transform -1 0 28896 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0855_
timestamp 1751889408
transform 1 0 19936 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0856_
timestamp 1751889408
transform 1 0 21168 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0857_
timestamp 1752345181
transform -1 0 12768 0 1 32928
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0858_
timestamp 1753172561
transform -1 0 16912 0 -1 36064
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0859_
timestamp 1752345181
transform -1 0 20496 0 1 34496
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0860_
timestamp 1753182340
transform 1 0 17920 0 -1 32928
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0861_
timestamp 1751534193
transform 1 0 20272 0 1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0862_
timestamp 1753172561
transform -1 0 24640 0 1 31360
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _0863_
timestamp 1752061876
transform 1 0 23744 0 -1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0864_
timestamp 1753277515
transform -1 0 26656 0 -1 28224
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0865_
timestamp 1751534193
transform -1 0 25760 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0866_
timestamp 1751889408
transform -1 0 25760 0 1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0867_
timestamp 1751534193
transform 1 0 24192 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _0868_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753579406
transform 1 0 20272 0 -1 18816
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0869_
timestamp 1753182340
transform -1 0 19712 0 1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0870_
timestamp 1751534193
transform 1 0 19712 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0871_
timestamp 1751534193
transform 1 0 26208 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0872_
timestamp 1753182340
transform -1 0 25984 0 1 26656
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0873_
timestamp 1753960525
transform 1 0 25088 0 -1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0874_
timestamp 1751889408
transform -1 0 27552 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0875_
timestamp 1753960525
transform 1 0 26656 0 -1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0876_
timestamp 1751534193
transform 1 0 27776 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0877_
timestamp 1751889408
transform 1 0 26992 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0878_
timestamp 1751914308
transform 1 0 27328 0 -1 15680
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0879_
timestamp 1751534193
transform -1 0 28672 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0880_
timestamp 1751534193
transform 1 0 16688 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0881_
timestamp 1751889408
transform -1 0 16800 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0882_
timestamp 1751534193
transform -1 0 16576 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _0883_
timestamp 1752061876
transform -1 0 24976 0 1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0884_
timestamp 1751531619
transform -1 0 29792 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_4  _0885_
timestamp 1751882821
transform -1 0 26544 0 -1 23520
box -86 -86 1542 870
use gf180mcu_as_sc_mcu7t3v3__buff_8  _0886_
timestamp 1752063767
transform -1 0 13888 0 -1 21952
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_8  _0887_
timestamp 1752063767
transform -1 0 7840 0 -1 25088
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0888_
timestamp 1751914308
transform 1 0 13328 0 1 23520
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0889_
timestamp 1751889408
transform 1 0 14560 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0890_
timestamp 1752063729
transform 1 0 14000 0 1 21952
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0891_
timestamp 1751531619
transform -1 0 28784 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0892_
timestamp 1751889808
transform 1 0 27552 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0893_
timestamp 1751914308
transform -1 0 31696 0 1 32928
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0894_
timestamp 1751889808
transform 1 0 28000 0 1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0895_
timestamp 1752063729
transform 1 0 29008 0 1 34496
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0896_
timestamp 1753172561
transform 1 0 26432 0 1 23520
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _0897_
timestamp 1752061876
transform -1 0 28560 0 1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0898_
timestamp 1751914308
transform 1 0 29008 0 1 32928
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0899_
timestamp 1751889808
transform 1 0 29008 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0900_
timestamp 1751534193
transform 1 0 31696 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0901_
timestamp 1752345181
transform 1 0 25424 0 -1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0902_
timestamp 1751914308
transform -1 0 26768 0 1 14112
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0903_
timestamp 1751534193
transform -1 0 25760 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0904_
timestamp 1751914308
transform -1 0 10752 0 -1 23520
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0905_
timestamp 1751889408
transform -1 0 8288 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0906_
timestamp 1752063729
transform 1 0 8176 0 1 20384
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0907_
timestamp 1751914308
transform -1 0 9184 0 -1 25088
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0908_
timestamp 1751889408
transform -1 0 7168 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0909_
timestamp 1752063729
transform 1 0 7168 0 -1 23520
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0910_
timestamp 1751534193
transform -1 0 6160 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0911_
timestamp 1751914308
transform -1 0 7056 0 1 25088
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0912_
timestamp 1751889408
transform -1 0 5264 0 1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0913_
timestamp 1752063729
transform 1 0 4368 0 -1 28224
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_8  _0914_
timestamp 1752063767
transform -1 0 5040 0 1 23520
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0915_
timestamp 1751914308
transform 1 0 1568 0 1 29792
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0916_
timestamp 1751889408
transform 1 0 4368 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0917_
timestamp 1752063729
transform -1 0 4928 0 1 29792
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0918_
timestamp 1751914308
transform 1 0 1680 0 -1 31360
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0919_
timestamp 1751889408
transform 1 0 6048 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0920_
timestamp 1752063729
transform -1 0 4368 0 1 31360
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0921_
timestamp 1751914308
transform -1 0 5824 0 -1 29792
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0922_
timestamp 1751889408
transform -1 0 3584 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0923_
timestamp 1752063729
transform 1 0 2464 0 -1 29792
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0924_
timestamp 1751534193
transform -1 0 4704 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0925_
timestamp 1751914308
transform 1 0 2800 0 -1 26656
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0926_
timestamp 1751889408
transform 1 0 5040 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0927_
timestamp 1752063729
transform -1 0 4032 0 1 25088
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_8  _0928_
timestamp 1752063767
transform -1 0 5264 0 1 21952
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0929_
timestamp 1751914308
transform -1 0 6384 0 -1 21952
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0930_
timestamp 1751889408
transform -1 0 3248 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0931_
timestamp 1752063729
transform 1 0 2016 0 1 20384
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0932_
timestamp 1751914308
transform -1 0 8176 0 1 20384
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0933_
timestamp 1751889408
transform -1 0 4144 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0934_
timestamp 1752063729
transform 1 0 3248 0 1 18816
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0935_
timestamp 1751914308
transform -1 0 6832 0 1 20384
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0936_
timestamp 1751889408
transform -1 0 5264 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0937_
timestamp 1752063729
transform 1 0 5488 0 1 18816
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0938_
timestamp 1751534193
transform -1 0 12544 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0939_
timestamp 1751534193
transform -1 0 11424 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0940_
timestamp 1751914308
transform 1 0 7168 0 -1 20384
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0941_
timestamp 1751889408
transform 1 0 9408 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0942_
timestamp 1752063729
transform -1 0 9744 0 1 17248
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0943_
timestamp 1751534193
transform -1 0 14560 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0944_
timestamp 1751914308
transform -1 0 12656 0 -1 18816
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0945_
timestamp 1751889408
transform -1 0 11312 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0946_
timestamp 1752063729
transform 1 0 9856 0 -1 17248
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0947_
timestamp 1751914308
transform 1 0 12208 0 -1 17248
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0948_
timestamp 1751889408
transform 1 0 13328 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0949_
timestamp 1752063729
transform 1 0 13328 0 1 15680
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0950_
timestamp 1751914308
transform 1 0 11760 0 1 18816
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0951_
timestamp 1751889408
transform 1 0 12880 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0952_
timestamp 1752063729
transform 1 0 13776 0 -1 18816
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0953_
timestamp 1751534193
transform 1 0 10752 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0954_
timestamp 1751914308
transform -1 0 14672 0 1 20384
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0955_
timestamp 1751889408
transform -1 0 11872 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0956_
timestamp 1752063729
transform 1 0 11088 0 1 20384
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0957_
timestamp 1751914308
transform -1 0 13104 0 1 23520
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0958_
timestamp 1751889408
transform 1 0 11872 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0959_
timestamp 1751534193
transform -1 0 12768 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0960_
timestamp 1751532043
transform -1 0 9968 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0961_
timestamp 1751532043
transform 1 0 10528 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0962_
timestamp 1751534193
transform 1 0 19600 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0963_
timestamp 1751534193
transform 1 0 17360 0 1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0964_
timestamp 1751534193
transform -1 0 17920 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0965_
timestamp 1753441877
transform 1 0 11088 0 -1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0966_
timestamp 1751534193
transform -1 0 11760 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0967_
timestamp 1751531619
transform -1 0 10976 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0968_
timestamp 1753960525
transform -1 0 11088 0 -1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0969_
timestamp 1753371985
transform -1 0 11088 0 1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0970_
timestamp 1751740063
transform -1 0 8176 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0971_
timestamp 1751534193
transform 1 0 6720 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0972_
timestamp 1751914308
transform 1 0 7504 0 -1 28224
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0973_
timestamp 1751534193
transform -1 0 10864 0 -1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0974_
timestamp 1753441877
transform -1 0 9072 0 1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0975_
timestamp 1753868718
transform -1 0 9408 0 1 28224
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0976_
timestamp 1751889408
transform -1 0 8736 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0977_
timestamp 1752063729
transform -1 0 7168 0 -1 34496
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0978_
timestamp 1751531619
transform 1 0 9408 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0979_
timestamp 1751740063
transform -1 0 7840 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0980_
timestamp 1751914308
transform 1 0 6720 0 1 29792
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0981_
timestamp 1752063729
transform -1 0 14224 0 -1 28224
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0982_
timestamp 1753441877
transform -1 0 10416 0 1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0983_
timestamp 1753868718
transform -1 0 9296 0 1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0984_
timestamp 1751889408
transform -1 0 8624 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0985_
timestamp 1752063729
transform -1 0 4144 0 1 34496
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0986_
timestamp 1751534193
transform -1 0 10864 0 1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0987_
timestamp 1751534193
transform -1 0 12320 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0988_
timestamp 1751534193
transform -1 0 11536 0 1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0989_
timestamp 1751740063
transform -1 0 7840 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0990_
timestamp 1751914308
transform 1 0 6944 0 1 31360
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0991_
timestamp 1753441877
transform -1 0 10528 0 -1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0992_
timestamp 1753868718
transform -1 0 10864 0 1 31360
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0993_
timestamp 1751889408
transform -1 0 9184 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _0994_
timestamp 1752063729
transform 1 0 9408 0 -1 34496
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0995_
timestamp 1751534193
transform -1 0 12544 0 -1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0996_
timestamp 1751532043
transform 1 0 7168 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0997_
timestamp 1751889808
transform 1 0 8400 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0998_
timestamp 1751740063
transform 1 0 7616 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0999_
timestamp 1751914308
transform 1 0 8288 0 1 31360
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1000_
timestamp 1751534193
transform 1 0 10864 0 -1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1001_
timestamp 1753441877
transform -1 0 11984 0 1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1002_
timestamp 1753868718
transform -1 0 10640 0 -1 32928
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1003_
timestamp 1751889408
transform -1 0 9632 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1004_
timestamp 1751534193
transform -1 0 9184 0 1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1005_
timestamp 1751531619
transform 1 0 10640 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1006_
timestamp 1751740063
transform 1 0 11424 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1007_
timestamp 1752061876
transform 1 0 11984 0 1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1008_
timestamp 1751914308
transform -1 0 12768 0 -1 31360
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1009_
timestamp 1751532043
transform -1 0 13776 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1010_
timestamp 1753441877
transform 1 0 11984 0 1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1011_
timestamp 1753868718
transform 1 0 13328 0 1 31360
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1012_
timestamp 1751889408
transform -1 0 14112 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _1013_
timestamp 1752063729
transform -1 0 14224 0 -1 32928
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1014_
timestamp 1751889808
transform 1 0 14560 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1015_
timestamp 1751914308
transform 1 0 13888 0 1 29792
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1016_
timestamp 1751740063
transform 1 0 16128 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1017_
timestamp 1751531619
transform 1 0 14224 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1018_
timestamp 1753371985
transform 1 0 15456 0 -1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1019_
timestamp 1751740063
transform 1 0 15456 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1020_
timestamp 1753182340
transform -1 0 18480 0 -1 34496
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1021_
timestamp 1751534193
transform -1 0 17472 0 1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1022_
timestamp 1751534193
transform 1 0 22960 0 1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1023_
timestamp 1751532043
transform -1 0 17024 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1024_
timestamp 1751740063
transform -1 0 17024 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1025_
timestamp 1751889408
transform -1 0 16128 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1026_
timestamp 1751914308
transform 1 0 12880 0 -1 29792
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1027_
timestamp 1753441877
transform 1 0 13104 0 -1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1028_
timestamp 1753868718
transform 1 0 14224 0 -1 31360
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1029_
timestamp 1751889408
transform 1 0 14224 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _1030_
timestamp 1752063729
transform 1 0 13888 0 1 34496
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1031_
timestamp 1751534193
transform 1 0 16352 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1032_
timestamp 1751531619
transform -1 0 18032 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1033_
timestamp 1753441877
transform -1 0 18256 0 1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1034_
timestamp 1753182340
transform -1 0 15904 0 -1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1035_
timestamp 1751914308
transform -1 0 15120 0 1 26656
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1036_
timestamp 1751889408
transform -1 0 17024 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1037_
timestamp 1753960525
transform 1 0 16016 0 1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1038_
timestamp 1751534193
transform 1 0 17584 0 1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1039_
timestamp 1751534193
transform -1 0 23184 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1040_
timestamp 1753960525
transform 1 0 19152 0 -1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1041_
timestamp 1753441877
transform 1 0 20272 0 -1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1042_
timestamp 1751532043
transform 1 0 9408 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1043_
timestamp 1751534193
transform -1 0 19712 0 1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1044_
timestamp 1751914308
transform 1 0 18816 0 1 28224
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1045_
timestamp 1753371985
transform 1 0 21168 0 1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1046_
timestamp 1751889408
transform 1 0 21392 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1047_
timestamp 1751534193
transform 1 0 22288 0 1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1048_
timestamp 1751532043
transform -1 0 18816 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1049_
timestamp 1753441877
transform 1 0 18592 0 -1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1050_
timestamp 1752061876
transform -1 0 22512 0 -1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1051_
timestamp 1751914308
transform 1 0 15120 0 1 26656
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1052_
timestamp 1751889408
transform -1 0 19152 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1053_
timestamp 1753960525
transform 1 0 19040 0 -1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1054_
timestamp 1751534193
transform 1 0 23968 0 1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1055_
timestamp 1751531619
transform -1 0 20944 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1056_
timestamp 1751740063
transform -1 0 18144 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1057_
timestamp 1751534193
transform 1 0 17248 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1058_
timestamp 1751914308
transform 1 0 17360 0 1 23520
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1059_
timestamp 1751889408
transform -1 0 19376 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1060_
timestamp 1751534193
transform 1 0 17920 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1061_
timestamp 1753441877
transform -1 0 19824 0 1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1062_
timestamp 1753868718
transform 1 0 18144 0 -1 25088
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1063_
timestamp 1751534193
transform 1 0 20384 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1064_
timestamp 1751532043
transform -1 0 18704 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1065_
timestamp 1751889408
transform -1 0 20496 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1066_
timestamp 1751889408
transform 1 0 17808 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1067_
timestamp 1753960525
transform 1 0 18704 0 1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1068_
timestamp 1751889408
transform -1 0 20608 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1069_
timestamp 1751532043
transform 1 0 20496 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1070_
timestamp 1753441877
transform 1 0 19152 0 1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1071_
timestamp 1753868718
transform 1 0 19376 0 -1 25088
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1072_
timestamp 1751534193
transform 1 0 20608 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1073_
timestamp 1751534193
transform -1 0 24192 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1074_
timestamp 1753441877
transform 1 0 19936 0 -1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1075_
timestamp 1751531619
transform 1 0 21056 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1076_
timestamp 1751531619
transform -1 0 21952 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1077_
timestamp 1751532043
transform 1 0 18144 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1078_
timestamp 1751532043
transform -1 0 22960 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _1079_
timestamp 1752345181
transform -1 0 21392 0 -1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1080_
timestamp 1751914308
transform 1 0 19264 0 -1 26656
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1081_
timestamp 1751740063
transform -1 0 21616 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1082_
timestamp 1753960525
transform 1 0 21392 0 1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1083_
timestamp 1751534193
transform 1 0 23408 0 -1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1084_
timestamp 1751532043
transform 1 0 15008 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1085_
timestamp 1751532043
transform -1 0 23744 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _1086_
timestamp 1753172561
transform -1 0 23520 0 -1 31360
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1087_
timestamp 1751914308
transform 1 0 15232 0 1 29792
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1088_
timestamp 1751889808
transform 1 0 21168 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1089_
timestamp 1753960525
transform -1 0 23072 0 1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1090_
timestamp 1753441877
transform 1 0 21952 0 1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1091_
timestamp 1753371985
transform 1 0 22176 0 -1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1092_
timestamp 1751531619
transform 1 0 15344 0 1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1093_
timestamp 1753960525
transform 1 0 23968 0 1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1094_
timestamp 1751889808
transform 1 0 25984 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1095_
timestamp 1753441877
transform 1 0 23632 0 1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1096_
timestamp 1753441877
transform 1 0 24640 0 1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1097_
timestamp 1751531619
transform 1 0 25200 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1098_
timestamp 1753371985
transform 1 0 25312 0 -1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1099_
timestamp 1751534193
transform -1 0 10976 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1100_
timestamp 1751889408
transform -1 0 14672 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1101_
timestamp 1751914308
transform -1 0 12432 0 -1 12544
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1102_
timestamp 1751889408
transform 1 0 10976 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _1103_
timestamp 1752063729
transform 1 0 11088 0 1 12544
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1104_
timestamp 1751889408
transform -1 0 11088 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1105_
timestamp 1751914308
transform -1 0 10864 0 -1 14112
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1106_
timestamp 1751889408
transform -1 0 9184 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _1107_
timestamp 1752063729
transform -1 0 9184 0 -1 14112
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1108_
timestamp 1751534193
transform -1 0 7728 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1109_
timestamp 1751889408
transform -1 0 10192 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_4  _1110_
timestamp 1751546029
transform -1 0 13888 0 -1 12544
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1111_
timestamp 1751914308
transform 1 0 7728 0 -1 12544
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1112_
timestamp 1751889408
transform -1 0 9632 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _1113_
timestamp 1752063729
transform -1 0 8064 0 -1 10976
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1114_
timestamp 1751889408
transform 1 0 8400 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1115_
timestamp 1751914308
transform -1 0 9856 0 1 9408
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1116_
timestamp 1751889408
transform -1 0 8400 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _1117_
timestamp 1752063729
transform -1 0 7168 0 -1 9408
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1118_
timestamp 1751889408
transform 1 0 7056 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1119_
timestamp 1751914308
transform 1 0 7504 0 1 7840
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1120_
timestamp 1751889408
transform -1 0 9632 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _1121_
timestamp 1752063729
transform -1 0 8176 0 1 6272
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1122_
timestamp 1751889408
transform 1 0 9408 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1123_
timestamp 1751914308
transform 1 0 7840 0 -1 7840
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1124_
timestamp 1751889408
transform -1 0 10976 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  _1125_
timestamp 1752063729
transform -1 0 10192 0 1 6272
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751632746
transform -1 0 17360 0 1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1127_
timestamp 1751632746
transform -1 0 12544 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1128_
timestamp 1751632746
transform -1 0 15232 0 -1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1129_
timestamp 1751632746
transform 1 0 10976 0 -1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1130_
timestamp 1751632746
transform 1 0 12544 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1131_
timestamp 1751632746
transform 1 0 15456 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1132_
timestamp 1751632746
transform 1 0 17248 0 -1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1133_
timestamp 1751632746
transform 1 0 17920 0 1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1134_
timestamp 1751632746
transform 1 0 18480 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1135_
timestamp 1751632746
transform -1 0 24528 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1136_
timestamp 1751632746
transform 1 0 21840 0 -1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1137_
timestamp 1751632746
transform 1 0 24752 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1138_
timestamp 1751632746
transform 1 0 26880 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1139_
timestamp 1751632746
transform 1 0 29904 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1140_
timestamp 1751632746
transform 1 0 32928 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1141_
timestamp 1751632746
transform 1 0 35392 0 -1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1142_
timestamp 1751632746
transform -1 0 38416 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1143_
timestamp 1751632746
transform 1 0 33936 0 -1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1144_
timestamp 1751632746
transform 1 0 22400 0 1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1145_
timestamp 1751632746
transform 1 0 25088 0 -1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1146_
timestamp 1751632746
transform -1 0 32032 0 1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1147_
timestamp 1751632746
transform 1 0 30016 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1148_
timestamp 1751632746
transform 1 0 33040 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1149_
timestamp 1751632746
transform -1 0 38416 0 -1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1150_
timestamp 1751632746
transform 1 0 34496 0 -1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1151_
timestamp 1751632746
transform 1 0 33600 0 1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1152_
timestamp 1751632746
transform 1 0 24976 0 1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1153_
timestamp 1751632746
transform -1 0 28336 0 -1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1154_
timestamp 1751632746
transform 1 0 25760 0 1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1155_
timestamp 1751632746
transform 1 0 17248 0 -1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1156_
timestamp 1751632746
transform 1 0 28784 0 -1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1157_
timestamp 1751632746
transform 1 0 27216 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1158_
timestamp 1751632746
transform 1 0 19600 0 -1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1159_
timestamp 1751632746
transform 1 0 17920 0 1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1160_
timestamp 1751632746
transform 1 0 16912 0 1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1161_
timestamp 1751632746
transform 1 0 17248 0 -1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1162_
timestamp 1751632746
transform 1 0 25088 0 -1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1163_
timestamp 1751632746
transform 1 0 15008 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1164_
timestamp 1751632746
transform 1 0 34272 0 -1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1165_
timestamp 1751632746
transform 1 0 34720 0 -1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1166_
timestamp 1751632746
transform -1 0 38416 0 -1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1167_
timestamp 1751632746
transform 1 0 16016 0 1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1168_
timestamp 1751632746
transform 1 0 31696 0 1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1169_
timestamp 1751632746
transform 1 0 32928 0 -1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1170_
timestamp 1751632746
transform 1 0 35280 0 -1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1171_
timestamp 1751632746
transform -1 0 36624 0 1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1172_
timestamp 1751632746
transform 1 0 29344 0 -1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1173_
timestamp 1751632746
transform 1 0 31024 0 1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1174_
timestamp 1751632746
transform -1 0 31696 0 -1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1175_
timestamp 1751632746
transform 1 0 23520 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1176_
timestamp 1751632746
transform 1 0 8288 0 1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1177_
timestamp 1751632746
transform -1 0 9968 0 1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1178_
timestamp 1751632746
transform 1 0 4480 0 -1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1179_
timestamp 1751632746
transform 1 0 3024 0 -1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1180_
timestamp 1751632746
transform 1 0 2352 0 -1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1181_
timestamp 1751632746
transform 1 0 2240 0 1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1182_
timestamp 1751632746
transform 1 0 2016 0 -1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1183_
timestamp 1751632746
transform 1 0 2016 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1184_
timestamp 1751632746
transform 1 0 4144 0 -1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1185_
timestamp 1751632746
transform 1 0 5712 0 -1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1186_
timestamp 1751632746
transform 1 0 7952 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1187_
timestamp 1751632746
transform 1 0 9968 0 1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1188_
timestamp 1751632746
transform 1 0 13664 0 -1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1189_
timestamp 1751632746
transform 1 0 14448 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1190_
timestamp 1751632746
transform 1 0 11984 0 -1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1191_
timestamp 1751632746
transform 1 0 11536 0 -1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1192_
timestamp 1751632746
transform 1 0 9072 0 1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1193_
timestamp 1751632746
transform 1 0 5488 0 1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1194_
timestamp 1751632746
transform 1 0 2464 0 -1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1195_
timestamp 1751632746
transform 1 0 10080 0 1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1196_
timestamp 1751632746
transform 1 0 6160 0 -1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1197_
timestamp 1751632746
transform 1 0 12320 0 -1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1198_
timestamp 1751632746
transform 1 0 15904 0 1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1199_
timestamp 1751632746
transform 1 0 17248 0 -1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1200_
timestamp 1751632746
transform 1 0 17248 0 1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1201_
timestamp 1751632746
transform -1 0 23744 0 -1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1202_
timestamp 1751632746
transform -1 0 23632 0 1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1203_
timestamp 1751632746
transform 1 0 21168 0 1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1204_
timestamp 1751632746
transform 1 0 21280 0 -1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1205_
timestamp 1751632746
transform 1 0 23744 0 1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1206_
timestamp 1751632746
transform 1 0 21840 0 -1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1207_
timestamp 1751632746
transform 1 0 25984 0 -1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1208_
timestamp 1751632746
transform -1 0 14224 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1209_
timestamp 1751632746
transform 1 0 7056 0 1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1210_
timestamp 1751632746
transform 1 0 5824 0 1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1211_
timestamp 1751632746
transform 1 0 5488 0 1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1212_
timestamp 1751632746
transform 1 0 5824 0 -1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1213_
timestamp 1751632746
transform -1 0 11088 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1222_
timestamp 1751534193
transform 1 0 31024 0 1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1223_
timestamp 1751534193
transform -1 0 35392 0 1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1224_
timestamp 1751534193
transform -1 0 35504 0 1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1225_
timestamp 1751534193
transform 1 0 35728 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1226_
timestamp 1751534193
transform 1 0 35392 0 1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1227_
timestamp 1751534193
transform 1 0 36400 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1228_
timestamp 1751534193
transform -1 0 9968 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1229_
timestamp 1751534193
transform -1 0 3584 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1230_
timestamp 1751534193
transform -1 0 6160 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1231_
timestamp 1751534193
transform -1 0 6720 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1232_
timestamp 1751534193
transform -1 0 7392 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1233_
timestamp 1751534193
transform -1 0 8064 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0563__A dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532392
transform 1 0 19936 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0569__B
timestamp 1751532392
transform 1 0 24416 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0569__C
timestamp 1751532392
transform 1 0 24416 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0572__A
timestamp 1751532392
transform 1 0 23408 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0582__A
timestamp 1751532392
transform -1 0 18928 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0586__A
timestamp 1751532392
transform -1 0 24528 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0588__A
timestamp 1751532392
transform 1 0 23968 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0593__A
timestamp 1751532392
transform 1 0 19712 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0595__A
timestamp 1751532392
transform 1 0 15008 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0596__A
timestamp 1751532392
transform 1 0 24640 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0609__A
timestamp 1751532392
transform -1 0 28784 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0613__A
timestamp 1751532392
transform 1 0 35952 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0616__A
timestamp 1751532392
transform 1 0 30240 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0629__A
timestamp 1751532392
transform 1 0 18816 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0633__A
timestamp 1751532392
transform 1 0 31248 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0649__A
timestamp 1751532392
transform 1 0 36624 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0651__A
timestamp 1751532392
transform 1 0 14224 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0654__B
timestamp 1751532392
transform 1 0 29568 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0655__A
timestamp 1751532392
transform 1 0 36288 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0662__A
timestamp 1751532392
transform -1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0666__A
timestamp 1751532392
transform -1 0 25984 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0685__S
timestamp 1751532392
transform 1 0 38192 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0687__B
timestamp 1751532392
transform 1 0 22960 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0690__A
timestamp 1751532392
transform 1 0 31024 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0692__B
timestamp 1751532392
transform 1 0 31920 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0694__B
timestamp 1751532392
transform 1 0 27328 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0696__A
timestamp 1751532392
transform 1 0 23296 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0696__B
timestamp 1751532392
transform 1 0 22848 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0701__A
timestamp 1751532392
transform 1 0 31024 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0706__A
timestamp 1751532392
transform 1 0 13552 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0708__A
timestamp 1751532392
transform 1 0 34496 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0713__A
timestamp 1751532392
transform -1 0 15120 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0713__C
timestamp 1751532392
transform 1 0 15680 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0715__A
timestamp 1751532392
transform -1 0 12880 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0716__A
timestamp 1751532392
transform -1 0 14560 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0718__A
timestamp 1751532392
transform -1 0 15008 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0719__A
timestamp 1751532392
transform 1 0 10080 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0726__A
timestamp 1751532392
transform 1 0 17472 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0727__B
timestamp 1751532392
transform -1 0 15120 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0741__A
timestamp 1751532392
transform 1 0 20384 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0798__A
timestamp 1751532392
transform 1 0 29568 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0804__C
timestamp 1751532392
transform 1 0 32256 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0818__A
timestamp 1751532392
transform -1 0 15344 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0821__A
timestamp 1751532392
transform 1 0 30576 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0827__A
timestamp 1751532392
transform -1 0 34048 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0831__A
timestamp 1751532392
transform -1 0 35392 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0835__A
timestamp 1751532392
transform 1 0 36400 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0837__A
timestamp 1751532392
transform 1 0 9632 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0840__A
timestamp 1751532392
transform 1 0 33712 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0844__A
timestamp 1751532392
transform 1 0 24640 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0847__A
timestamp 1751532392
transform -1 0 28336 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0851__A
timestamp 1751532392
transform 1 0 12992 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0855__A
timestamp 1751532392
transform 1 0 20944 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0863__A
timestamp 1751532392
transform 1 0 24416 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0866__A
timestamp 1751532392
transform -1 0 26656 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0872__B
timestamp 1751532392
transform 1 0 27104 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0872__C
timestamp 1751532392
transform 1 0 27776 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0874__A
timestamp 1751532392
transform 1 0 28224 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0878__B
timestamp 1751532392
transform -1 0 29456 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0881__B
timestamp 1751532392
transform 1 0 17584 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0883__B
timestamp 1751532392
transform -1 0 26208 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0889__B
timestamp 1751532392
transform -1 0 16240 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0893__A
timestamp 1751532392
transform 1 0 36176 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0898__B
timestamp 1751532392
transform 1 0 24192 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0902__A
timestamp 1751532392
transform -1 0 27216 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0904__B
timestamp 1751532392
transform 1 0 10752 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0905__B
timestamp 1751532392
transform 1 0 8288 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0908__B
timestamp 1751532392
transform -1 0 6384 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0910__A
timestamp 1751532392
transform 1 0 6384 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0924__A
timestamp 1751532392
transform 1 0 4928 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0925__A
timestamp 1751532392
transform 1 0 4144 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0929__B
timestamp 1751532392
transform 1 0 6608 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0939__A
timestamp 1751532392
transform 1 0 11648 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0953__A
timestamp 1751532392
transform 1 0 11424 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0966__A
timestamp 1751532392
transform 1 0 12656 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0968__D
timestamp 1751532392
transform -1 0 11424 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0971__A
timestamp 1751532392
transform -1 0 6720 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0986__A
timestamp 1751532392
transform -1 0 10192 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0995__A
timestamp 1751532392
transform 1 0 13552 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1000__A
timestamp 1751532392
transform -1 0 11536 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1010__C
timestamp 1751532392
transform -1 0 11984 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1015__A
timestamp 1751532392
transform 1 0 14448 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1027__C
timestamp 1751532392
transform -1 0 15456 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1037__B
timestamp 1751532392
transform -1 0 17696 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1039__A
timestamp 1751532392
transform 1 0 23408 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1044__A
timestamp 1751532392
transform -1 0 18816 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1053__B
timestamp 1751532392
transform 1 0 18144 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1056__A
timestamp 1751532392
transform 1 0 18032 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1059__A
timestamp 1751532392
transform -1 0 19600 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1076__A
timestamp 1751532392
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1082__B
timestamp 1751532392
transform 1 0 22064 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1093__D
timestamp 1751532392
transform -1 0 27216 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1097__A
timestamp 1751532392
transform 1 0 26992 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1099__A
timestamp 1751532392
transform -1 0 12208 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1100__A
timestamp 1751532392
transform 1 0 14112 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1108__A
timestamp 1751532392
transform 1 0 7728 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1120__A
timestamp 1751532392
transform 1 0 9856 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1124__A
timestamp 1751532392
transform 1 0 10976 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1126__CLK
timestamp 1751532392
transform 1 0 17472 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1128__CLK
timestamp 1751532392
transform 1 0 15456 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1131__CLK
timestamp 1751532392
transform 1 0 18704 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1132__CLK
timestamp 1751532392
transform 1 0 17024 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1133__CLK
timestamp 1751532392
transform 1 0 17696 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1134__CLK
timestamp 1751532392
transform 1 0 18256 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1140__CLK
timestamp 1751532392
transform -1 0 37296 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1141__CLK
timestamp 1751532392
transform -1 0 36400 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1142__CLK
timestamp 1751532392
transform 1 0 35168 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1143__CLK
timestamp 1751532392
transform 1 0 37184 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1146__CLK
timestamp 1751532392
transform 1 0 32256 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1148__CLK
timestamp 1751532392
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1149__CLK
timestamp 1751532392
transform 1 0 35168 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1150__CLK
timestamp 1751532392
transform 1 0 33600 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1151__CLK
timestamp 1751532392
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1152__CLK
timestamp 1751532392
transform 1 0 20720 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1154__CLK
timestamp 1751532392
transform 1 0 29120 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1158__D
timestamp 1751532392
transform 1 0 22960 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1159__D
timestamp 1751532392
transform -1 0 21168 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1160__D
timestamp 1751532392
transform -1 0 18144 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1161__D
timestamp 1751532392
transform 1 0 23856 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1163__CLK
timestamp 1751532392
transform 1 0 18256 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1166__CLK
timestamp 1751532392
transform 1 0 35168 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1167__CLK
timestamp 1751532392
transform 1 0 15792 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1171__CLK
timestamp 1751532392
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1176__CLK
timestamp 1751532392
transform 1 0 7280 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1177__CLK
timestamp 1751532392
transform 1 0 10192 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1178__CLK
timestamp 1751532392
transform 1 0 7728 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1179__CLK
timestamp 1751532392
transform 1 0 6048 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1180__CLK
timestamp 1751532392
transform 1 0 5600 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1181__CLK
timestamp 1751532392
transform 1 0 5712 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1182__CLK
timestamp 1751532392
transform 1 0 4256 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1183__CLK
timestamp 1751532392
transform 1 0 5712 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1184__CLK
timestamp 1751532392
transform 1 0 7728 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1185__CLK
timestamp 1751532392
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1186__CLK
timestamp 1751532392
transform 1 0 11200 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1187__CLK
timestamp 1751532392
transform -1 0 15232 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1188__CLK
timestamp 1751532392
transform 1 0 17472 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1189__CLK
timestamp 1751532392
transform 1 0 17696 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1190__CLK
timestamp 1751532392
transform 1 0 15232 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1191__CLK
timestamp 1751532392
transform 1 0 15568 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1192__CLK
timestamp 1751532392
transform 1 0 13552 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1193__CLK
timestamp 1751532392
transform 1 0 9408 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1194__CLK
timestamp 1751532392
transform -1 0 5936 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1195__CLK
timestamp 1751532392
transform 1 0 9856 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1196__CLK
timestamp 1751532392
transform -1 0 9856 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1197__CLK
timestamp 1751532392
transform -1 0 11088 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1198__CLK
timestamp 1751532392
transform 1 0 13664 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1199__CLK
timestamp 1751532392
transform 1 0 18704 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1200__CLK
timestamp 1751532392
transform 1 0 17024 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1201__CLK
timestamp 1751532392
transform 1 0 23968 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1202__CLK
timestamp 1751532392
transform 1 0 23856 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1203__CLK
timestamp 1751532392
transform -1 0 24640 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1204__CLK
timestamp 1751532392
transform 1 0 24528 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1205__CLK
timestamp 1751532392
transform 1 0 28672 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1206__CLK
timestamp 1751532392
transform 1 0 24640 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1207__CLK
timestamp 1751532392
transform 1 0 29232 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1208__CLK
timestamp 1751532392
transform 1 0 14448 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1223__A
timestamp 1751532392
transform 1 0 36288 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1229__A
timestamp 1751532392
transform -1 0 2912 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_0_clk_i_A
timestamp 1751532392
transform -1 0 24192 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_0__f_clk_i_A
timestamp 1751532392
transform 1 0 12880 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_1__f_clk_i_A
timestamp 1751532392
transform -1 0 18368 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_2__f_clk_i_A
timestamp 1751532392
transform 1 0 10080 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_3__f_clk_i_A
timestamp 1751532392
transform 1 0 14896 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_4__f_clk_i_A
timestamp 1751532392
transform 1 0 28000 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_5__f_clk_i_A
timestamp 1751532392
transform 1 0 32256 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_6__f_clk_i_A
timestamp 1751532392
transform 1 0 25424 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_7__f_clk_i_A
timestamp 1751532392
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload1_A
timestamp 1751532392
transform 1 0 15008 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload2_A
timestamp 1751532392
transform 1 0 12768 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload4_A
timestamp 1751532392
transform 1 0 33712 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload5_A
timestamp 1751532392
transform 1 0 24192 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_fanout58_A
timestamp 1751532392
transform 1 0 21392 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input1_A
timestamp 1751532392
transform -1 0 37968 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input2_A
timestamp 1751532392
transform -1 0 37744 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input3_A
timestamp 1751532392
transform -1 0 37744 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input4_A
timestamp 1751532392
transform -1 0 37744 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input5_A
timestamp 1751532392
transform -1 0 37744 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input6_A
timestamp 1751532392
transform -1 0 37744 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input7_A
timestamp 1751532392
transform -1 0 37744 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input8_A
timestamp 1751532392
transform -1 0 38416 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input9_A
timestamp 1751532392
transform -1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input10_A
timestamp 1751532392
transform -1 0 38416 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input11_A
timestamp 1751532392
transform -1 0 38416 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input12_A
timestamp 1751532392
transform 1 0 29120 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input13_A
timestamp 1751532392
transform 1 0 29568 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input14_A
timestamp 1751532392
transform 1 0 30800 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input15_A
timestamp 1751532392
transform 1 0 31584 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input16_A
timestamp 1751532392
transform -1 0 33488 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input17_A
timestamp 1751532392
transform 1 0 35392 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input18_A
timestamp 1751532392
transform -1 0 37072 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input19_A
timestamp 1751532392
transform -1 0 37968 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_output29_A
timestamp 1751532392
transform 1 0 36064 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_output30_A
timestamp 1751532392
transform -1 0 20720 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_output33_A
timestamp 1751532392
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0_clk_i dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751661108
transform -1 0 23968 0 1 20384
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_0__f_clk_i
timestamp 1751661108
transform 1 0 10752 0 -1 10976
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_1__f_clk_i
timestamp 1751661108
transform 1 0 15344 0 1 9408
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_2__f_clk_i
timestamp 1751661108
transform -1 0 9856 0 1 25088
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_3__f_clk_i
timestamp 1751661108
transform 1 0 11872 0 -1 26656
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_4__f_clk_i
timestamp 1751661108
transform 1 0 28224 0 -1 12544
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_5__f_clk_i
timestamp 1751661108
transform 1 0 32480 0 1 14112
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_6__f_clk_i
timestamp 1751661108
transform 1 0 25648 0 -1 29792
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_7__f_clk_i
timestamp 1751661108
transform -1 0 32928 0 1 29792
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload0 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751896485
transform 1 0 10640 0 1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_4  clkload1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751633659
transform 1 0 15232 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  clkload2
timestamp 1751532043
transform 1 0 12096 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload3
timestamp 1751896485
transform -1 0 28784 0 1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  clkload4
timestamp 1751532043
transform 1 0 32928 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkload5
timestamp 1751661108
transform 1 0 25648 0 1 31360
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkload6
timestamp 1751661108
transform 1 0 29904 0 -1 31360
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout58
timestamp 1751534193
transform -1 0 20496 0 1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout59
timestamp 1751534193
transform -1 0 19936 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout60
timestamp 1751534193
transform -1 0 17920 0 -1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout61
timestamp 1751534193
transform -1 0 13776 0 1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout62
timestamp 1751534193
transform -1 0 8848 0 1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout63
timestamp 1751534193
transform 1 0 10416 0 1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout64
timestamp 1751534193
transform 1 0 11760 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_8  fanout65
timestamp 1752063767
transform -1 0 19264 0 -1 12544
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_8  fanout66
timestamp 1752063767
transform -1 0 20944 0 1 12544
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__buff_8  fanout67
timestamp 1752063767
transform 1 0 20160 0 -1 14112
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532246
transform 1 0 1568 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_6 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532440
transform 1 0 2016 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_8 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532423
transform 1 0 2240 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_36
timestamp 1751532423
transform 1 0 5376 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_70
timestamp 1751532423
transform 1 0 9184 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_138
timestamp 1751532246
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_142
timestamp 1751532440
transform 1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_144
timestamp 1751532423
transform 1 0 17472 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_172
timestamp 1751532440
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_174
timestamp 1751532423
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_200
timestamp 1751532246
transform 1 0 23744 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_237
timestamp 1751532423
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_246
timestamp 1751532440
transform 1 0 28896 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_250
timestamp 1751532440
transform 1 0 29344 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_254
timestamp 1751532423
transform 1 0 29792 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_261
timestamp 1751532440
transform 1 0 30576 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_265
timestamp 1751532246
transform 1 0 31024 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_269
timestamp 1751532423
transform 1 0 31472 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_280
timestamp 1751532246
transform 1 0 32704 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_284
timestamp 1751532423
transform 1 0 33152 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_0_293 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532312
transform 1 0 34160 0 1 3136
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_301
timestamp 1751532440
transform 1 0 35056 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_303
timestamp 1751532423
transform 1 0 35280 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_314
timestamp 1751532440
transform 1 0 36512 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_316
timestamp 1751532423
transform 1 0 36736 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_1_2
timestamp 1751532312
transform 1 0 1568 0 -1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_10
timestamp 1751532440
transform 1 0 2464 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_72
timestamp 1751532440
transform 1 0 9408 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_74
timestamp 1751532423
transform 1 0 9632 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_127
timestamp 1751532423
transform 1 0 15568 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_149
timestamp 1751532440
transform 1 0 18032 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_207
timestamp 1751532440
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_209
timestamp 1751532423
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_1_212
timestamp 1751532312
transform 1 0 25088 0 -1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_227
timestamp 1751532423
transform 1 0 26768 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_273
timestamp 1751532246
transform 1 0 31920 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_277
timestamp 1751532440
transform 1 0 32368 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_279
timestamp 1751532423
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_1_312
timestamp 1751532312
transform 1 0 36288 0 -1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_320
timestamp 1751532246
transform 1 0 37184 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_324
timestamp 1751532423
transform 1 0 37632 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_327
timestamp 1751532440
transform 1 0 37968 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_2_27
timestamp 1751532312
transform 1 0 4368 0 1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_2_37
timestamp 1751532246
transform 1 0 5488 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_41
timestamp 1751532423
transform 1 0 5936 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_107
timestamp 1751532423
transform 1 0 13328 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_153
timestamp 1751532440
transform 1 0 18480 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_2_177
timestamp 1751532246
transform 1 0 21168 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_181
timestamp 1751532423
transform 1 0 21616 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_2_200
timestamp 1751532312
transform 1 0 23744 0 1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_208
timestamp 1751532423
transform 1 0 24640 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_2_236
timestamp 1751532312
transform 1 0 27776 0 1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_244
timestamp 1751532423
transform 1 0 28672 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_2_247
timestamp 1751532312
transform 1 0 29008 0 1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_309
timestamp 1751532440
transform 1 0 35952 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_313
timestamp 1751532440
transform 1 0 36400 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_317
timestamp 1751532440
transform 1 0 36848 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_321
timestamp 1751532440
transform 1 0 37296 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532351
transform 1 0 1568 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_18
timestamp 1751532351
transform 1 0 3360 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_34
timestamp 1751532246
transform 1 0 5152 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_38
timestamp 1751532440
transform 1 0 5600 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_67
timestamp 1751532440
transform 1 0 8848 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_69
timestamp 1751532423
transform 1 0 9072 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_72
timestamp 1751532440
transform 1 0 9408 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_138
timestamp 1751532440
transform 1 0 16800 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_142
timestamp 1751532423
transform 1 0 17248 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_175
timestamp 1751532440
transform 1 0 20944 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_177
timestamp 1751532423
transform 1 0 21168 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_197
timestamp 1751532246
transform 1 0 23408 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_201
timestamp 1751532440
transform 1 0 23856 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_294
timestamp 1751532440
transform 1 0 34272 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_296
timestamp 1751532423
transform 1 0 34496 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_2
timestamp 1751532351
transform 1 0 1568 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_18
timestamp 1751532351
transform 1 0 3360 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_34
timestamp 1751532423
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_4_37
timestamp 1751532246
transform 1 0 5488 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_41
timestamp 1751532440
transform 1 0 5936 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_86
timestamp 1751532423
transform 1 0 10976 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_4_119
timestamp 1751532246
transform 1 0 14672 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_153
timestamp 1751532440
transform 1 0 18480 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_174
timestamp 1751532423
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_183
timestamp 1751532440
transform 1 0 21840 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_4_203
timestamp 1751532246
transform 1 0 24080 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_207
timestamp 1751532423
transform 1 0 24528 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_244
timestamp 1751532423
transform 1 0 28672 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_247
timestamp 1751532440
transform 1 0 29008 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_249
timestamp 1751532423
transform 1 0 29232 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_4_269
timestamp 1751532312
transform 1 0 31472 0 1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_4_277
timestamp 1751532246
transform 1 0 32368 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_281
timestamp 1751532440
transform 1 0 32816 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_283
timestamp 1751532423
transform 1 0 33040 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_296
timestamp 1751532423
transform 1 0 34496 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_329
timestamp 1751532440
transform 1 0 38192 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_2
timestamp 1751532351
transform 1 0 1568 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_18
timestamp 1751532351
transform 1 0 3360 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_34
timestamp 1751532351
transform 1 0 5152 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_50
timestamp 1751532423
transform 1 0 6944 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_79
timestamp 1751532246
transform 1 0 10192 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_83
timestamp 1751532440
transform 1 0 10640 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_85
timestamp 1751532423
transform 1 0 10864 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_88
timestamp 1751532440
transform 1 0 11200 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_124
timestamp 1751532440
transform 1 0 15232 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_128
timestamp 1751532246
transform 1 0 15680 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_132
timestamp 1751532423
transform 1 0 16128 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_181
timestamp 1751532440
transform 1 0 21616 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_212
timestamp 1751532423
transform 1 0 25088 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_5_249
timestamp 1751532312
transform 1 0 29232 0 -1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_257
timestamp 1751532440
transform 1 0 30128 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_5_265
timestamp 1751532312
transform 1 0 31024 0 -1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_273
timestamp 1751532246
transform 1 0 31920 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_277
timestamp 1751532440
transform 1 0 32368 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_279
timestamp 1751532423
transform 1 0 32592 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_5_282
timestamp 1751532312
transform 1 0 32928 0 -1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_290
timestamp 1751532440
transform 1 0 33824 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_292
timestamp 1751532423
transform 1 0 34048 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_323
timestamp 1751532440
transform 1 0 37520 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_2
timestamp 1751532351
transform 1 0 1568 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_18
timestamp 1751532351
transform 1 0 3360 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_34
timestamp 1751532423
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_37
timestamp 1751532351
transform 1 0 5488 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_53
timestamp 1751532440
transform 1 0 7280 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_74
timestamp 1751532440
transform 1 0 9632 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_78
timestamp 1751532312
transform 1 0 10080 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_86
timestamp 1751532440
transform 1 0 10976 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_88
timestamp 1751532423
transform 1 0 11200 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_96
timestamp 1751532312
transform 1 0 12096 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_104
timestamp 1751532423
transform 1 0 12992 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_119
timestamp 1751532440
transform 1 0 14672 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_123
timestamp 1751532351
transform 1 0 15120 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_139
timestamp 1751532423
transform 1 0 16912 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_142
timestamp 1751532246
transform 1 0 17248 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_177
timestamp 1751532312
transform 1 0 21168 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_185
timestamp 1751532423
transform 1 0 22064 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_199
timestamp 1751532351
transform 1 0 23632 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_215
timestamp 1751532246
transform 1 0 25424 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_233
timestamp 1751532312
transform 1 0 27440 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_241
timestamp 1751532246
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_253
timestamp 1751532246
transform 1 0 29680 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_281
timestamp 1751532312
transform 1 0 32816 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_289
timestamp 1751532246
transform 1 0 33712 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_312
timestamp 1751532440
transform 1 0 36288 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_314
timestamp 1751532423
transform 1 0 36512 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_329
timestamp 1751532440
transform 1 0 38192 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_2
timestamp 1751532351
transform 1 0 1568 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_18
timestamp 1751532351
transform 1 0 3360 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_52
timestamp 1751532246
transform 1 0 7168 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_72
timestamp 1751532423
transform 1 0 9408 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_100
timestamp 1751532440
transform 1 0 12544 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_120
timestamp 1751532440
transform 1 0 14784 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_142
timestamp 1751532440
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_146
timestamp 1751532246
transform 1 0 17696 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_152
timestamp 1751532440
transform 1 0 18368 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_154
timestamp 1751532423
transform 1 0 18592 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_173
timestamp 1751532351
transform 1 0 20720 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_189
timestamp 1751532351
transform 1 0 22512 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_205
timestamp 1751532246
transform 1 0 24304 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_209
timestamp 1751532423
transform 1 0 24752 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_212
timestamp 1751532246
transform 1 0 25088 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_216
timestamp 1751532440
transform 1 0 25536 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_261
timestamp 1751532423
transform 1 0 30576 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_282
timestamp 1751532351
transform 1 0 32928 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_298
timestamp 1751532246
transform 1 0 34720 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_2
timestamp 1751532351
transform 1 0 1568 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_18
timestamp 1751532351
transform 1 0 3360 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_34
timestamp 1751532423
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_76
timestamp 1751532440
transform 1 0 9856 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_80
timestamp 1751532423
transform 1 0 10304 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_99
timestamp 1751532246
transform 1 0 12432 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_114
timestamp 1751532440
transform 1 0 14112 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_118
timestamp 1751532440
transform 1 0 14560 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_122
timestamp 1751532440
transform 1 0 15008 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_124
timestamp 1751532423
transform 1 0 15232 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_168
timestamp 1751532440
transform 1 0 20160 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_172
timestamp 1751532440
transform 1 0 20608 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_174
timestamp 1751532423
transform 1 0 20832 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_8_177
timestamp 1751532312
transform 1 0 21168 0 1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_185
timestamp 1751532440
transform 1 0 22064 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_187
timestamp 1751532423
transform 1 0 22288 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_215
timestamp 1751532440
transform 1 0 25424 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_241
timestamp 1751532246
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_274
timestamp 1751532440
transform 1 0 32032 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_278
timestamp 1751532423
transform 1 0 32480 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_8_304
timestamp 1751532312
transform 1 0 35392 0 1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_312
timestamp 1751532440
transform 1 0 36288 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_314
timestamp 1751532423
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_329
timestamp 1751532440
transform 1 0 38192 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_2
timestamp 1751532351
transform 1 0 1568 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_18
timestamp 1751532351
transform 1 0 3360 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_9_34
timestamp 1751532312
transform 1 0 5152 0 -1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_60
timestamp 1751532440
transform 1 0 8064 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_62
timestamp 1751532423
transform 1 0 8288 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_109
timestamp 1751532423
transform 1 0 13552 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_134
timestamp 1751532246
transform 1 0 16352 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_138
timestamp 1751532440
transform 1 0 16800 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_142
timestamp 1751532440
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_9_146
timestamp 1751532312
transform 1 0 17696 0 -1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_154
timestamp 1751532440
transform 1 0 18592 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_170
timestamp 1751532246
transform 1 0 20384 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_174
timestamp 1751532423
transform 1 0 20832 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_177
timestamp 1751532351
transform 1 0 21168 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_193
timestamp 1751532440
transform 1 0 22960 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_195
timestamp 1751532423
transform 1 0 23184 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_9_202
timestamp 1751532312
transform 1 0 23968 0 -1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_245
timestamp 1751532440
transform 1 0 28784 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_9_266
timestamp 1751532312
transform 1 0 31136 0 -1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_274
timestamp 1751532246
transform 1 0 32032 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_278
timestamp 1751532440
transform 1 0 32480 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_9_282
timestamp 1751532312
transform 1 0 32928 0 -1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_290
timestamp 1751532423
transform 1 0 33824 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_318
timestamp 1751532440
transform 1 0 36960 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_9_322
timestamp 1751532312
transform 1 0 37408 0 -1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_330
timestamp 1751532423
transform 1 0 38304 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_2
timestamp 1751532351
transform 1 0 1568 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_18
timestamp 1751532351
transform 1 0 3360 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_34
timestamp 1751532423
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_37
timestamp 1751532440
transform 1 0 5488 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_39
timestamp 1751532423
transform 1 0 5712 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_74
timestamp 1751532440
transform 1 0 9632 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_107
timestamp 1751532440
transform 1 0 13328 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_143
timestamp 1751532440
transform 1 0 17360 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_147
timestamp 1751532423
transform 1 0 17808 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_191
timestamp 1751532440
transform 1 0 22736 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_195
timestamp 1751532351
transform 1 0 23184 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_10_211
timestamp 1751532312
transform 1 0 24976 0 1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_232
timestamp 1751532246
transform 1 0 27328 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_236
timestamp 1751532440
transform 1 0 27776 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_240
timestamp 1751532246
transform 1 0 28224 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_244
timestamp 1751532423
transform 1 0 28672 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_247
timestamp 1751532246
transform 1 0 29008 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_263
timestamp 1751532351
transform 1 0 30800 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_279
timestamp 1751532351
transform 1 0 32592 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_295
timestamp 1751532246
transform 1 0 34384 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_299
timestamp 1751532440
transform 1 0 34832 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_301
timestamp 1751532423
transform 1 0 35056 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_10_304
timestamp 1751532312
transform 1 0 35392 0 1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_312
timestamp 1751532440
transform 1 0 36288 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_314
timestamp 1751532423
transform 1 0 36512 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_317
timestamp 1751532246
transform 1 0 36848 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_321
timestamp 1751532440
transform 1 0 37296 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_2
timestamp 1751532351
transform 1 0 1568 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_18
timestamp 1751532351
transform 1 0 3360 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_34
timestamp 1751532351
transform 1 0 5152 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_50
timestamp 1751532423
transform 1 0 6944 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_69
timestamp 1751532423
transform 1 0 9072 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_79
timestamp 1751532440
transform 1 0 10192 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_99
timestamp 1751532440
transform 1 0 12432 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_119
timestamp 1751532440
transform 1 0 14672 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_121
timestamp 1751532423
transform 1 0 14896 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_138
timestamp 1751532440
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_160
timestamp 1751532440
transform 1 0 19264 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_162
timestamp 1751532423
transform 1 0 19488 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_190
timestamp 1751532440
transform 1 0 22624 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_194
timestamp 1751532440
transform 1 0 23072 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_11_198
timestamp 1751532312
transform 1 0 23520 0 -1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_206
timestamp 1751532246
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_239
timestamp 1751532423
transform 1 0 28112 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_277
timestamp 1751532440
transform 1 0 32368 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_279
timestamp 1751532423
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_11_282
timestamp 1751532312
transform 1 0 32928 0 -1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_299
timestamp 1751532440
transform 1 0 34832 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_301
timestamp 1751532423
transform 1 0 35056 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_12_2
timestamp 1751532351
transform 1 0 1568 0 1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_12_18
timestamp 1751532351
transform 1 0 3360 0 1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_34
timestamp 1751532423
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_12_37
timestamp 1751532351
transform 1 0 5488 0 1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_53
timestamp 1751532246
transform 1 0 7280 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_59
timestamp 1751532246
transform 1 0 7952 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_70
timestamp 1751532423
transform 1 0 9184 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_107
timestamp 1751532440
transform 1 0 13328 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_111
timestamp 1751532440
transform 1 0 13776 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_113
timestamp 1751532423
transform 1 0 14000 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_149
timestamp 1751532440
transform 1 0 18032 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_153
timestamp 1751532246
transform 1 0 18480 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_225
timestamp 1751532312
transform 1 0 26544 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_233
timestamp 1751532440
transform 1 0 27440 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_247
timestamp 1751532440
transform 1 0 29008 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_249
timestamp 1751532423
transform 1 0 29232 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_295
timestamp 1751532423
transform 1 0 34384 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_329
timestamp 1751532440
transform 1 0 38192 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_2
timestamp 1751532351
transform 1 0 1568 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_18
timestamp 1751532351
transform 1 0 3360 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_34
timestamp 1751532351
transform 1 0 5152 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_50
timestamp 1751532440
transform 1 0 6944 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_72
timestamp 1751532423
transform 1 0 9408 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_85
timestamp 1751532440
transform 1 0 10864 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_87
timestamp 1751532423
transform 1 0 11088 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_115
timestamp 1751532440
transform 1 0 14224 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_119
timestamp 1751532440
transform 1 0 14672 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_121
timestamp 1751532423
transform 1 0 14896 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_124
timestamp 1751532246
transform 1 0 15232 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_128
timestamp 1751532440
transform 1 0 15680 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_136
timestamp 1751532246
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_142
timestamp 1751532246
transform 1 0 17248 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_146
timestamp 1751532440
transform 1 0 17696 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_198
timestamp 1751532440
transform 1 0 23520 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_204
timestamp 1751532440
transform 1 0 24192 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_208
timestamp 1751532440
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_224
timestamp 1751532246
transform 1 0 26432 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_228
timestamp 1751532440
transform 1 0 26880 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_230
timestamp 1751532423
transform 1 0 27104 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_258
timestamp 1751532440
transform 1 0 30240 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_260
timestamp 1751532423
transform 1 0 30464 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_276
timestamp 1751532246
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_282
timestamp 1751532423
transform 1 0 32928 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_328
timestamp 1751532440
transform 1 0 38080 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_330
timestamp 1751532423
transform 1 0 38304 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_2
timestamp 1751532351
transform 1 0 1568 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_18
timestamp 1751532351
transform 1 0 3360 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_34
timestamp 1751532423
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_14_37
timestamp 1751532312
transform 1 0 5488 0 1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_45
timestamp 1751532246
transform 1 0 6384 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_49
timestamp 1751532440
transform 1 0 6832 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_78
timestamp 1751532440
transform 1 0 10080 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_93
timestamp 1751532440
transform 1 0 11760 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_14_97
timestamp 1751532312
transform 1 0 12208 0 1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_113
timestamp 1751532440
transform 1 0 14000 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_117
timestamp 1751532351
transform 1 0 14448 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_133
timestamp 1751532246
transform 1 0 16240 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_137
timestamp 1751532440
transform 1 0 16688 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_166
timestamp 1751532423
transform 1 0 19936 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_174
timestamp 1751532423
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_200
timestamp 1751532440
transform 1 0 23744 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_204
timestamp 1751532440
transform 1 0 24192 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_227
timestamp 1751532440
transform 1 0 26768 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_231
timestamp 1751532246
transform 1 0 27216 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_235
timestamp 1751532440
transform 1 0 27664 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_237
timestamp 1751532423
transform 1 0 27888 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_244
timestamp 1751532423
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_247
timestamp 1751532440
transform 1 0 29008 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_251
timestamp 1751532351
transform 1 0 29456 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_267
timestamp 1751532440
transform 1 0 31248 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_275
timestamp 1751532440
transform 1 0 32144 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_277
timestamp 1751532423
transform 1 0 32368 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_317
timestamp 1751532440
transform 1 0 36848 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_321
timestamp 1751532440
transform 1 0 37296 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_2
timestamp 1751532351
transform 1 0 1568 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_18
timestamp 1751532351
transform 1 0 3360 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_34
timestamp 1751532351
transform 1 0 5152 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_50
timestamp 1751532351
transform 1 0 6944 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_66
timestamp 1751532246
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_72
timestamp 1751532351
transform 1 0 9408 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_88
timestamp 1751532246
transform 1 0 11200 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_92
timestamp 1751532440
transform 1 0 11648 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_100
timestamp 1751532351
transform 1 0 12544 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_116
timestamp 1751532246
transform 1 0 14336 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_120
timestamp 1751532440
transform 1 0 14784 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_122
timestamp 1751532423
transform 1 0 15008 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_125
timestamp 1751532312
transform 1 0 15344 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_133
timestamp 1751532246
transform 1 0 16240 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_137
timestamp 1751532440
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_139
timestamp 1751532423
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_169
timestamp 1751532440
transform 1 0 20272 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_199
timestamp 1751532440
transform 1 0 23632 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_203
timestamp 1751532440
transform 1 0 24080 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_207
timestamp 1751532440
transform 1 0 24528 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_209
timestamp 1751532423
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_212
timestamp 1751532440
transform 1 0 25088 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_218
timestamp 1751532312
transform 1 0 25760 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_226
timestamp 1751532246
transform 1 0 26656 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_230
timestamp 1751532440
transform 1 0 27104 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_244
timestamp 1751532423
transform 1 0 28672 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_272
timestamp 1751532246
transform 1 0 31808 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_278
timestamp 1751532440
transform 1 0 32480 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_286
timestamp 1751532440
transform 1 0 33376 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_288
timestamp 1751532423
transform 1 0 33600 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_313
timestamp 1751532351
transform 1 0 36400 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_329
timestamp 1751532440
transform 1 0 38192 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_2
timestamp 1751532351
transform 1 0 1568 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_18
timestamp 1751532351
transform 1 0 3360 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_34
timestamp 1751532423
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_37
timestamp 1751532351
transform 1 0 5488 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_53
timestamp 1751532351
transform 1 0 7280 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_69
timestamp 1751532312
transform 1 0 9072 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_77
timestamp 1751532246
transform 1 0 9968 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_81
timestamp 1751532440
transform 1 0 10416 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_83
timestamp 1751532423
transform 1 0 10640 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_90
timestamp 1751532440
transform 1 0 11424 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_94
timestamp 1751532312
transform 1 0 11872 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_102
timestamp 1751532440
transform 1 0 12768 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_104
timestamp 1751532423
transform 1 0 12992 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_131
timestamp 1751532351
transform 1 0 16016 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_147
timestamp 1751532440
transform 1 0 17808 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_195
timestamp 1751532440
transform 1 0 23184 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_199
timestamp 1751532246
transform 1 0 23632 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_217
timestamp 1751532312
transform 1 0 25648 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_225
timestamp 1751532246
transform 1 0 26544 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_229
timestamp 1751532440
transform 1 0 26992 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_231
timestamp 1751532423
transform 1 0 27216 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_271
timestamp 1751532440
transform 1 0 31696 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_275
timestamp 1751532246
transform 1 0 32144 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_279
timestamp 1751532440
transform 1 0 32592 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_287
timestamp 1751532440
transform 1 0 33488 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_297
timestamp 1751532440
transform 1 0 34608 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_311
timestamp 1751532440
transform 1 0 36176 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_324
timestamp 1751532246
transform 1 0 37632 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_328
timestamp 1751532440
transform 1 0 38080 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_330
timestamp 1751532423
transform 1 0 38304 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_2
timestamp 1751532351
transform 1 0 1568 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_18
timestamp 1751532351
transform 1 0 3360 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_34
timestamp 1751532351
transform 1 0 5152 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_50
timestamp 1751532312
transform 1 0 6944 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_58
timestamp 1751532246
transform 1 0 7840 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_62
timestamp 1751532423
transform 1 0 8288 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_69
timestamp 1751532423
transform 1 0 9072 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_72
timestamp 1751532440
transform 1 0 9408 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_94
timestamp 1751532440
transform 1 0 11872 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_96
timestamp 1751532423
transform 1 0 12096 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_109
timestamp 1751532423
transform 1 0 13552 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_137
timestamp 1751532440
transform 1 0 16688 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_139
timestamp 1751532423
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_142
timestamp 1751532440
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_146
timestamp 1751532312
transform 1 0 17696 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_154
timestamp 1751532423
transform 1 0 18592 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_157
timestamp 1751532440
transform 1 0 18928 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_191
timestamp 1751532440
transform 1 0 22736 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_195
timestamp 1751532440
transform 1 0 23184 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_204
timestamp 1751532246
transform 1 0 24192 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_208
timestamp 1751532440
transform 1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_212
timestamp 1751532440
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_214
timestamp 1751532423
transform 1 0 25312 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_225
timestamp 1751532312
transform 1 0 26544 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_233
timestamp 1751532440
transform 1 0 27440 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_235
timestamp 1751532423
transform 1 0 27664 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_263
timestamp 1751532440
transform 1 0 30800 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_267
timestamp 1751532312
transform 1 0 31248 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_275
timestamp 1751532246
transform 1 0 32144 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_279
timestamp 1751532423
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_282
timestamp 1751532246
transform 1 0 32928 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_286
timestamp 1751532440
transform 1 0 33376 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_323
timestamp 1751532312
transform 1 0 37520 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_2
timestamp 1751532351
transform 1 0 1568 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_18
timestamp 1751532351
transform 1 0 3360 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_34
timestamp 1751532423
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_37
timestamp 1751532351
transform 1 0 5488 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_53
timestamp 1751532246
transform 1 0 7280 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_75
timestamp 1751532440
transform 1 0 9744 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_104
timestamp 1751532423
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_120
timestamp 1751532440
transform 1 0 14784 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_124
timestamp 1751532351
transform 1 0 15232 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_140
timestamp 1751532246
transform 1 0 17024 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_144
timestamp 1751532423
transform 1 0 17472 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_18_151
timestamp 1751532312
transform 1 0 18256 0 1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_159
timestamp 1751532246
transform 1 0 19152 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_163
timestamp 1751532440
transform 1 0 19600 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_165
timestamp 1751532423
transform 1 0 19824 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_174
timestamp 1751532423
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_177
timestamp 1751532351
transform 1 0 21168 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_193
timestamp 1751532246
transform 1 0 22960 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_197
timestamp 1751532440
transform 1 0 23408 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_199
timestamp 1751532423
transform 1 0 23632 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_207
timestamp 1751532246
transform 1 0 24528 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_18_231
timestamp 1751532312
transform 1 0 27216 0 1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_239
timestamp 1751532246
transform 1 0 28112 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_251
timestamp 1751532440
transform 1 0 29456 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_263
timestamp 1751532440
transform 1 0 30800 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_267
timestamp 1751532351
transform 1 0 31248 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_283
timestamp 1751532246
transform 1 0 33040 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_287
timestamp 1751532423
transform 1 0 33488 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_317
timestamp 1751532440
transform 1 0 36848 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_321
timestamp 1751532440
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_19_2
timestamp 1751532351
transform 1 0 1568 0 -1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_19_18
timestamp 1751532351
transform 1 0 3360 0 -1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_34
timestamp 1751532246
transform 1 0 5152 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_38
timestamp 1751532423
transform 1 0 5600 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_66
timestamp 1751532440
transform 1 0 8736 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_79
timestamp 1751532440
transform 1 0 10192 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_81
timestamp 1751532423
transform 1 0 10416 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_101
timestamp 1751532440
transform 1 0 12656 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_110
timestamp 1751532423
transform 1 0 13664 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_19_129
timestamp 1751532312
transform 1 0 15792 0 -1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_137
timestamp 1751532440
transform 1 0 16688 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_139
timestamp 1751532423
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_194
timestamp 1751532423
transform 1 0 23072 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_202
timestamp 1751532423
transform 1 0 23968 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_212
timestamp 1751532440
transform 1 0 25088 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_214
timestamp 1751532423
transform 1 0 25312 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_239
timestamp 1751532246
transform 1 0 28112 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_243
timestamp 1751532440
transform 1 0 28560 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_245
timestamp 1751532423
transform 1 0 28784 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_19_270
timestamp 1751532312
transform 1 0 31584 0 -1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_278
timestamp 1751532440
transform 1 0 32480 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_282
timestamp 1751532246
transform 1 0 32928 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_286
timestamp 1751532440
transform 1 0 33376 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_288
timestamp 1751532423
transform 1 0 33600 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_304
timestamp 1751532440
transform 1 0 35392 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_306
timestamp 1751532423
transform 1 0 35616 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_19_311
timestamp 1751532351
transform 1 0 36176 0 -1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_327
timestamp 1751532246
transform 1 0 37968 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_20_2
timestamp 1751532312
transform 1 0 1568 0 1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_10
timestamp 1751532246
transform 1 0 2464 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_14
timestamp 1751532440
transform 1 0 2912 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_16
timestamp 1751532423
transform 1 0 3136 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_55
timestamp 1751532440
transform 1 0 7504 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_86
timestamp 1751532440
transform 1 0 10976 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_90
timestamp 1751532440
transform 1 0 11424 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_92
timestamp 1751532423
transform 1 0 11648 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_144
timestamp 1751532440
transform 1 0 17472 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_148
timestamp 1751532246
transform 1 0 17920 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_152
timestamp 1751532423
transform 1 0 18368 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_199
timestamp 1751532423
transform 1 0 23632 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_20_236
timestamp 1751532312
transform 1 0 27776 0 1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_244
timestamp 1751532423
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_247
timestamp 1751532423
transform 1 0 29008 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_274
timestamp 1751532440
transform 1 0 32032 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_278
timestamp 1751532351
transform 1 0 32480 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_294
timestamp 1751532351
transform 1 0 34272 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_310
timestamp 1751532246
transform 1 0 36064 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_314
timestamp 1751532423
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_317
timestamp 1751532440
transform 1 0 36848 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_321
timestamp 1751532440
transform 1 0 37296 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_2
timestamp 1751532351
transform 1 0 1568 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_64
timestamp 1751532246
transform 1 0 8512 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_68
timestamp 1751532440
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_76
timestamp 1751532351
transform 1 0 9856 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_92
timestamp 1751532440
transform 1 0 11648 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_94
timestamp 1751532423
transform 1 0 11872 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_122
timestamp 1751532440
transform 1 0 15008 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_126
timestamp 1751532440
transform 1 0 15456 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_130
timestamp 1751532312
transform 1 0 15904 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_138
timestamp 1751532440
transform 1 0 16800 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_142
timestamp 1751532351
transform 1 0 17248 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_158
timestamp 1751532246
transform 1 0 19040 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_162
timestamp 1751532440
transform 1 0 19488 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_209
timestamp 1751532423
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_216
timestamp 1751532440
transform 1 0 25536 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_220
timestamp 1751532351
transform 1 0 25984 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_236
timestamp 1751532312
transform 1 0 27776 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_244
timestamp 1751532440
transform 1 0 28672 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_246
timestamp 1751532423
transform 1 0 28896 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_275
timestamp 1751532246
transform 1 0 32144 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_279
timestamp 1751532423
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_282
timestamp 1751532440
transform 1 0 32928 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_296
timestamp 1751532246
transform 1 0 34496 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_300
timestamp 1751532440
transform 1 0 34944 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_2
timestamp 1751532246
transform 1 0 1568 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_24
timestamp 1751532246
transform 1 0 4032 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_22_79
timestamp 1751532312
transform 1 0 10192 0 1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_119
timestamp 1751532440
transform 1 0 14672 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_123
timestamp 1751532351
transform 1 0 15120 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_139
timestamp 1751532351
transform 1 0 16912 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_155
timestamp 1751532440
transform 1 0 18704 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_157
timestamp 1751532423
transform 1 0 18928 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_212
timestamp 1751532440
transform 1 0 25088 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_227
timestamp 1751532440
transform 1 0 26768 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_22_231
timestamp 1751532312
transform 1 0 27216 0 1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_239
timestamp 1751532246
transform 1 0 28112 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_243
timestamp 1751532440
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_22_247
timestamp 1751532312
transform 1 0 29008 0 1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_255
timestamp 1751532440
transform 1 0 29904 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_257
timestamp 1751532423
transform 1 0 30128 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_281
timestamp 1751532246
transform 1 0 32816 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_285
timestamp 1751532440
transform 1 0 33264 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_287
timestamp 1751532423
transform 1 0 33488 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_329
timestamp 1751532440
transform 1 0 38192 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_2
timestamp 1751532246
transform 1 0 1568 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_45
timestamp 1751532440
transform 1 0 6384 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_49
timestamp 1751532312
transform 1 0 6832 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_57
timestamp 1751532246
transform 1 0 7728 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_61
timestamp 1751532423
transform 1 0 8176 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_64
timestamp 1751532246
transform 1 0 8512 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_68
timestamp 1751532440
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_72
timestamp 1751532312
transform 1 0 9408 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_80
timestamp 1751532246
transform 1 0 10304 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_84
timestamp 1751532440
transform 1 0 10752 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_86
timestamp 1751532423
transform 1 0 10976 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_118
timestamp 1751532312
transform 1 0 14560 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_126
timestamp 1751532440
transform 1 0 15456 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_128
timestamp 1751532423
transform 1 0 15680 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_131
timestamp 1751532312
transform 1 0 16016 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_139
timestamp 1751532423
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_142
timestamp 1751532312
transform 1 0 17248 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_154
timestamp 1751532440
transform 1 0 18592 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_162
timestamp 1751532440
transform 1 0 19488 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_166
timestamp 1751532312
transform 1 0 19936 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_174
timestamp 1751532246
transform 1 0 20832 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_178
timestamp 1751532440
transform 1 0 21280 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_180
timestamp 1751532423
transform 1 0 21504 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_187
timestamp 1751532312
transform 1 0 22288 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_195
timestamp 1751532246
transform 1 0 23184 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_199
timestamp 1751532440
transform 1 0 23632 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_201
timestamp 1751532423
transform 1 0 23856 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_204
timestamp 1751532246
transform 1 0 24192 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_208
timestamp 1751532440
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_219
timestamp 1751532423
transform 1 0 25872 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_248
timestamp 1751532246
transform 1 0 29120 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_252
timestamp 1751532440
transform 1 0 29568 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_265
timestamp 1751532440
transform 1 0 31024 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_282
timestamp 1751532440
transform 1 0 32928 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_327
timestamp 1751532246
transform 1 0 37968 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_2
timestamp 1751532312
transform 1 0 1568 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_37
timestamp 1751532440
transform 1 0 5488 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_41
timestamp 1751532312
transform 1 0 5936 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_49
timestamp 1751532246
transform 1 0 6832 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_89
timestamp 1751532246
transform 1 0 11312 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_93
timestamp 1751532423
transform 1 0 11760 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_101
timestamp 1751532246
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_107
timestamp 1751532246
transform 1 0 13328 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_111
timestamp 1751532440
transform 1 0 13776 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_158
timestamp 1751532440
transform 1 0 19040 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_160
timestamp 1751532423
transform 1 0 19264 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_169
timestamp 1751532246
transform 1 0 20272 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_173
timestamp 1751532440
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_24_177
timestamp 1751532351
transform 1 0 21168 0 1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_193
timestamp 1751532440
transform 1 0 22960 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_202
timestamp 1751532312
transform 1 0 23968 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_210
timestamp 1751532246
transform 1 0 24864 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_214
timestamp 1751532440
transform 1 0 25312 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_227
timestamp 1751532440
transform 1 0 26768 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_229
timestamp 1751532423
transform 1 0 26992 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_243
timestamp 1751532440
transform 1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_254
timestamp 1751532423
transform 1 0 29792 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_304
timestamp 1751532312
transform 1 0 35392 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_312
timestamp 1751532440
transform 1 0 36288 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_314
timestamp 1751532423
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_317
timestamp 1751532312
transform 1 0 36848 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_325
timestamp 1751532246
transform 1 0 37744 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_2
timestamp 1751532351
transform 1 0 1568 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_18
timestamp 1751532246
transform 1 0 3360 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_22
timestamp 1751532440
transform 1 0 3808 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_30
timestamp 1751532440
transform 1 0 4704 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_25_34
timestamp 1751532312
transform 1 0 5152 0 -1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_42
timestamp 1751532423
transform 1 0 6048 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_90
timestamp 1751532423
transform 1 0 11424 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_125
timestamp 1751532440
transform 1 0 15344 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_129
timestamp 1751532440
transform 1 0 15792 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_133
timestamp 1751532423
transform 1 0 16240 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_142
timestamp 1751532246
transform 1 0 17248 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_146
timestamp 1751532423
transform 1 0 17696 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_161
timestamp 1751532440
transform 1 0 19376 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_163
timestamp 1751532423
transform 1 0 19600 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_25_176
timestamp 1751532312
transform 1 0 21056 0 -1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_184
timestamp 1751532440
transform 1 0 21952 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_193
timestamp 1751532351
transform 1 0 22960 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_209
timestamp 1751532423
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_225
timestamp 1751532440
transform 1 0 26544 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_241
timestamp 1751532440
transform 1 0 28336 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_279
timestamp 1751532423
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_25_282
timestamp 1751532312
transform 1 0 32928 0 -1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_290
timestamp 1751532246
transform 1 0 33824 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_294
timestamp 1751532440
transform 1 0 34272 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_308
timestamp 1751532440
transform 1 0 35840 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_310
timestamp 1751532423
transform 1 0 36064 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_323
timestamp 1751532440
transform 1 0 37520 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_26_2
timestamp 1751532312
transform 1 0 1568 0 1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_10
timestamp 1751532246
transform 1 0 2464 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_14
timestamp 1751532423
transform 1 0 2912 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_33
timestamp 1751532440
transform 1 0 5040 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_43
timestamp 1751532440
transform 1 0 6160 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_47
timestamp 1751532440
transform 1 0 6608 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_49
timestamp 1751532423
transform 1 0 6832 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_77
timestamp 1751532440
transform 1 0 9968 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_81
timestamp 1751532440
transform 1 0 10416 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_83
timestamp 1751532423
transform 1 0 10640 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_86
timestamp 1751532246
transform 1 0 10976 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_92
timestamp 1751532423
transform 1 0 11648 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_26_125
timestamp 1751532312
transform 1 0 15344 0 1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_133
timestamp 1751532246
transform 1 0 16240 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_172
timestamp 1751532440
transform 1 0 20608 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_174
timestamp 1751532423
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_204
timestamp 1751532440
transform 1 0 24192 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_208
timestamp 1751532246
transform 1 0 24640 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_218
timestamp 1751532246
transform 1 0 25760 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_222
timestamp 1751532440
transform 1 0 26208 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_247
timestamp 1751532246
transform 1 0 29008 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_251
timestamp 1751532423
transform 1 0 29456 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_254
timestamp 1751532246
transform 1 0 29792 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_26_279
timestamp 1751532351
transform 1 0 32592 0 1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_295
timestamp 1751532423
transform 1 0 34384 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_329
timestamp 1751532440
transform 1 0 38192 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_27_2
timestamp 1751532246
transform 1 0 1568 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_72
timestamp 1751532351
transform 1 0 9408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_27_88
timestamp 1751532312
transform 1 0 11200 0 -1 25088
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_102
timestamp 1751532440
transform 1 0 12768 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_106
timestamp 1751532351
transform 1 0 13216 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_27_126
timestamp 1751532312
transform 1 0 15456 0 -1 25088
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_27_134
timestamp 1751532246
transform 1 0 16352 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_138
timestamp 1751532440
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_142
timestamp 1751532423
transform 1 0 17248 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_205
timestamp 1751532440
transform 1 0 24304 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_209
timestamp 1751532423
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_212
timestamp 1751532351
transform 1 0 25088 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_228
timestamp 1751532351
transform 1 0 26880 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_244
timestamp 1751532423
transform 1 0 28672 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_252
timestamp 1751532440
transform 1 0 29568 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_279
timestamp 1751532423
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_27_282
timestamp 1751532246
transform 1 0 32928 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_27_292
timestamp 1751532246
transform 1 0 34048 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_327
timestamp 1751532440
transform 1 0 37968 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_28_2
timestamp 1751532246
transform 1 0 1568 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_24
timestamp 1751532440
transform 1 0 4032 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_37
timestamp 1751532440
transform 1 0 5488 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_76
timestamp 1751532440
transform 1 0 9856 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_80
timestamp 1751532440
transform 1 0 10304 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_104
timestamp 1751532423
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_132
timestamp 1751532351
transform 1 0 16128 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_148
timestamp 1751532423
transform 1 0 17920 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_177
timestamp 1751532440
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_181
timestamp 1751532351
transform 1 0 21616 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_28_197
timestamp 1751532246
transform 1 0 23408 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_218
timestamp 1751532440
transform 1 0 25760 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_222
timestamp 1751532440
transform 1 0 26208 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_28_226
timestamp 1751532246
transform 1 0 26656 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_230
timestamp 1751532440
transform 1 0 27104 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_232
timestamp 1751532423
transform 1 0 27328 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_243
timestamp 1751532440
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_247
timestamp 1751532440
transform 1 0 29008 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_28_297
timestamp 1751532246
transform 1 0 34608 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_301
timestamp 1751532440
transform 1 0 35056 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_313
timestamp 1751532440
transform 1 0 36400 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_329
timestamp 1751532440
transform 1 0 38192 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_29_2
timestamp 1751532312
transform 1 0 1568 0 -1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_10
timestamp 1751532440
transform 1 0 2464 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_12
timestamp 1751532423
transform 1 0 2688 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_25
timestamp 1751532440
transform 1 0 4144 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_27
timestamp 1751532423
transform 1 0 4368 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_55
timestamp 1751532440
transform 1 0 7504 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_29_59
timestamp 1751532312
transform 1 0 7952 0 -1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_67
timestamp 1751532440
transform 1 0 8848 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_69
timestamp 1751532423
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_72
timestamp 1751532246
transform 1 0 9408 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_76
timestamp 1751532440
transform 1 0 9856 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_78
timestamp 1751532423
transform 1 0 10080 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_86
timestamp 1751532440
transform 1 0 10976 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_90
timestamp 1751532246
transform 1 0 11424 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_119
timestamp 1751532440
transform 1 0 14672 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_29_123
timestamp 1751532312
transform 1 0 15120 0 -1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_131
timestamp 1751532440
transform 1 0 16016 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_133
timestamp 1751532423
transform 1 0 16240 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_29_148
timestamp 1751532312
transform 1 0 17920 0 -1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_156
timestamp 1751532246
transform 1 0 18816 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_172
timestamp 1751532440
transform 1 0 20608 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_29_181
timestamp 1751532351
transform 1 0 21616 0 -1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_197
timestamp 1751532246
transform 1 0 23408 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_201
timestamp 1751532440
transform 1 0 23856 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_203
timestamp 1751532423
transform 1 0 24080 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_228
timestamp 1751532440
transform 1 0 26880 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_232
timestamp 1751532246
transform 1 0 27328 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_236
timestamp 1751532440
transform 1 0 27776 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_238
timestamp 1751532423
transform 1 0 28000 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_29_241
timestamp 1751532351
transform 1 0 28336 0 -1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_275
timestamp 1751532246
transform 1 0 32144 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_279
timestamp 1751532423
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_282
timestamp 1751532440
transform 1 0 32928 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_286
timestamp 1751532440
transform 1 0 33376 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_2
timestamp 1751532351
transform 1 0 1568 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_18
timestamp 1751532246
transform 1 0 3360 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_22
timestamp 1751532440
transform 1 0 3808 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_24
timestamp 1751532423
transform 1 0 4032 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_30_27
timestamp 1751532312
transform 1 0 4368 0 1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_37
timestamp 1751532351
transform 1 0 5488 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_53
timestamp 1751532246
transform 1 0 7280 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_57
timestamp 1751532440
transform 1 0 7728 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_100
timestamp 1751532440
transform 1 0 12544 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_104
timestamp 1751532423
transform 1 0 12992 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_107
timestamp 1751532440
transform 1 0 13328 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_30_135
timestamp 1751532312
transform 1 0 16464 0 1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_149
timestamp 1751532440
transform 1 0 18032 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_151
timestamp 1751532423
transform 1 0 18256 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_169
timestamp 1751532246
transform 1 0 20272 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_30_184
timestamp 1751532312
transform 1 0 21952 0 1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_192
timestamp 1751532246
transform 1 0 22848 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_196
timestamp 1751532440
transform 1 0 23296 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_198
timestamp 1751532423
transform 1 0 23520 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_234
timestamp 1751532440
transform 1 0 27552 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_238
timestamp 1751532440
transform 1 0 28000 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_242
timestamp 1751532440
transform 1 0 28448 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_244
timestamp 1751532423
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_247
timestamp 1751532440
transform 1 0 29008 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_251
timestamp 1751532246
transform 1 0 29456 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_255
timestamp 1751532440
transform 1 0 29904 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_257
timestamp 1751532423
transform 1 0 30128 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_307
timestamp 1751532246
transform 1 0 35728 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_311
timestamp 1751532440
transform 1 0 36176 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_329
timestamp 1751532440
transform 1 0 38192 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_31_2
timestamp 1751532312
transform 1 0 1568 0 -1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_10
timestamp 1751532440
transform 1 0 2464 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_12
timestamp 1751532423
transform 1 0 2688 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_20
timestamp 1751532246
transform 1 0 3584 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_24
timestamp 1751532440
transform 1 0 4032 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_26
timestamp 1751532423
transform 1 0 4256 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_31_45
timestamp 1751532312
transform 1 0 6384 0 -1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_53
timestamp 1751532440
transform 1 0 7280 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_67
timestamp 1751532440
transform 1 0 8848 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_69
timestamp 1751532423
transform 1 0 9072 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_72
timestamp 1751532423
transform 1 0 9408 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_115
timestamp 1751532440
transform 1 0 14224 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_117
timestamp 1751532423
transform 1 0 14448 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_31_124
timestamp 1751532312
transform 1 0 15232 0 -1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_132
timestamp 1751532423
transform 1 0 16128 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_164
timestamp 1751532440
transform 1 0 19712 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_183
timestamp 1751532440
transform 1 0 21840 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_31_187
timestamp 1751532312
transform 1 0 22288 0 -1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_195
timestamp 1751532246
transform 1 0 23184 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_199
timestamp 1751532423
transform 1 0 23632 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_246
timestamp 1751532440
transform 1 0 28896 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_250
timestamp 1751532440
transform 1 0 29344 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_267
timestamp 1751532423
transform 1 0 31248 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_294
timestamp 1751532246
transform 1 0 34272 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_32_2
timestamp 1751532246
transform 1 0 1568 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_6
timestamp 1751532440
transform 1 0 2016 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_37
timestamp 1751532440
transform 1 0 5488 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_32_41
timestamp 1751532246
transform 1 0 5936 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_45
timestamp 1751532423
transform 1 0 6384 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_32_72
timestamp 1751532246
transform 1 0 9408 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_76
timestamp 1751532423
transform 1 0 9856 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_99
timestamp 1751532440
transform 1 0 12432 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_103
timestamp 1751532440
transform 1 0 12880 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_107
timestamp 1751532440
transform 1 0 13328 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_111
timestamp 1751532351
transform 1 0 13776 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_32_127
timestamp 1751532246
transform 1 0 15568 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_151
timestamp 1751532423
transform 1 0 18256 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_177
timestamp 1751532440
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_195
timestamp 1751532440
transform 1 0 23184 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_32_199
timestamp 1751532246
transform 1 0 23632 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_203
timestamp 1751532440
transform 1 0 24080 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_205
timestamp 1751532423
transform 1 0 24304 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_247
timestamp 1751532440
transform 1 0 29008 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_279
timestamp 1751532440
transform 1 0 32592 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_288
timestamp 1751532440
transform 1 0 33600 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_329
timestamp 1751532440
transform 1 0 38192 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_33_2
timestamp 1751532312
transform 1 0 1568 0 -1 29792
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_33_40
timestamp 1751532312
transform 1 0 5824 0 -1 29792
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_48
timestamp 1751532440
transform 1 0 6720 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_50
timestamp 1751532423
transform 1 0 6944 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_58
timestamp 1751532423
transform 1 0 7840 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_66
timestamp 1751532246
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_91
timestamp 1751532440
transform 1 0 11536 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_93
timestamp 1751532423
transform 1 0 11760 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_100
timestamp 1751532440
transform 1 0 12544 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_102
timestamp 1751532423
transform 1 0 12768 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_115
timestamp 1751532440
transform 1 0 14224 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_33_130
timestamp 1751532312
transform 1 0 15904 0 -1 29792
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_138
timestamp 1751532440
transform 1 0 16800 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_142
timestamp 1751532440
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_146
timestamp 1751532246
transform 1 0 17696 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_152
timestamp 1751532440
transform 1 0 18368 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_156
timestamp 1751532440
transform 1 0 18816 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_193
timestamp 1751532246
transform 1 0 22960 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_203
timestamp 1751532246
transform 1 0 24080 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_207
timestamp 1751532423
transform 1 0 24528 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_212
timestamp 1751532440
transform 1 0 25088 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_214
timestamp 1751532423
transform 1 0 25312 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_242
timestamp 1751532440
transform 1 0 28448 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_277
timestamp 1751532440
transform 1 0 32368 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_279
timestamp 1751532423
transform 1 0 32592 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_282
timestamp 1751532440
transform 1 0 32928 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_286
timestamp 1751532423
transform 1 0 33376 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_330
timestamp 1751532423
transform 1 0 38304 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_32
timestamp 1751532440
transform 1 0 4928 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_34
timestamp 1751532423
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_37
timestamp 1751532246
transform 1 0 5488 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_41
timestamp 1751532423
transform 1 0 5936 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_44
timestamp 1751532246
transform 1 0 6272 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_87
timestamp 1751532440
transform 1 0 11088 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_91
timestamp 1751532440
transform 1 0 11536 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_111
timestamp 1751532423
transform 1 0 13776 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_136
timestamp 1751532246
transform 1 0 16576 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_142
timestamp 1751532440
transform 1 0 17248 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_144
timestamp 1751532423
transform 1 0 17472 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_151
timestamp 1751532246
transform 1 0 18256 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_155
timestamp 1751532440
transform 1 0 18704 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_157
timestamp 1751532423
transform 1 0 18928 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_171
timestamp 1751532246
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_194
timestamp 1751532246
transform 1 0 23072 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_198
timestamp 1751532440
transform 1 0 23520 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_227
timestamp 1751532440
transform 1 0 26768 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_231
timestamp 1751532440
transform 1 0 27216 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_247
timestamp 1751532440
transform 1 0 29008 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_249
timestamp 1751532423
transform 1 0 29232 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_307
timestamp 1751532440
transform 1 0 35728 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_311
timestamp 1751532246
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_329
timestamp 1751532440
transform 1 0 38192 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_2
timestamp 1751532423
transform 1 0 1568 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_49
timestamp 1751532440
transform 1 0 6832 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_65
timestamp 1751532246
transform 1 0 8624 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_69
timestamp 1751532423
transform 1 0 9072 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_35_82
timestamp 1751532312
transform 1 0 10528 0 -1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_102
timestamp 1751532440
transform 1 0 12768 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_104
timestamp 1751532423
transform 1 0 12992 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_35_149
timestamp 1751532312
transform 1 0 18032 0 -1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_157
timestamp 1751532440
transform 1 0 18928 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_159
timestamp 1751532423
transform 1 0 19152 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_173
timestamp 1751532440
transform 1 0 20720 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_204
timestamp 1751532246
transform 1 0 24192 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_212
timestamp 1751532423
transform 1 0 25088 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_254
timestamp 1751532423
transform 1 0 29792 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_327
timestamp 1751532246
transform 1 0 37968 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_36_2
timestamp 1751532246
transform 1 0 1568 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_6
timestamp 1751532440
transform 1 0 2016 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_8
timestamp 1751532423
transform 1 0 2240 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_34
timestamp 1751532423
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_36_37
timestamp 1751532312
transform 1 0 5488 0 1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_36_45
timestamp 1751532246
transform 1 0 6384 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_49
timestamp 1751532423
transform 1 0 6832 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_139
timestamp 1751532440
transform 1 0 16912 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_141
timestamp 1751532423
transform 1 0 17136 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_36_177
timestamp 1751532246
transform 1 0 21168 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_181
timestamp 1751532440
transform 1 0 21616 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_183
timestamp 1751532423
transform 1 0 21840 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_208
timestamp 1751532440
transform 1 0 24640 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_210
timestamp 1751532423
transform 1 0 24864 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_242
timestamp 1751532440
transform 1 0 28448 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_244
timestamp 1751532423
transform 1 0 28672 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_254
timestamp 1751532423
transform 1 0 29792 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_305
timestamp 1751532440
transform 1 0 35504 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_314
timestamp 1751532423
transform 1 0 36512 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_329
timestamp 1751532440
transform 1 0 38192 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_37_2
timestamp 1751532246
transform 1 0 1568 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_6
timestamp 1751532440
transform 1 0 2016 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_8
timestamp 1751532423
transform 1 0 2240 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_36
timestamp 1751532440
transform 1 0 5376 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_37_40
timestamp 1751532312
transform 1 0 5824 0 -1 32928
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_37_48
timestamp 1751532246
transform 1 0 6720 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_122
timestamp 1751532440
transform 1 0 15008 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_37_200
timestamp 1751532246
transform 1 0 23744 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_212
timestamp 1751532440
transform 1 0 25088 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_234
timestamp 1751532440
transform 1 0 27552 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_236
timestamp 1751532423
transform 1 0 27776 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_262
timestamp 1751532440
transform 1 0 30688 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_271
timestamp 1751532440
transform 1 0 31696 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_282
timestamp 1751532440
transform 1 0 32928 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_284
timestamp 1751532423
transform 1 0 33152 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_330
timestamp 1751532423
transform 1 0 38304 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_2
timestamp 1751532351
transform 1 0 1568 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_18
timestamp 1751532351
transform 1 0 3360 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_34
timestamp 1751532423
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_37
timestamp 1751532351
transform 1 0 5488 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_38_53
timestamp 1751532312
transform 1 0 7280 0 1 32928
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_74
timestamp 1751532440
transform 1 0 9632 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_76
timestamp 1751532423
transform 1 0 9856 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_102
timestamp 1751532440
transform 1 0 12768 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_104
timestamp 1751532423
transform 1 0 12992 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_114
timestamp 1751532423
transform 1 0 14112 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_172
timestamp 1751532440
transform 1 0 20608 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_174
timestamp 1751532423
transform 1 0 20832 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_38_199
timestamp 1751532246
transform 1 0 23632 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_203
timestamp 1751532423
transform 1 0 24080 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_206
timestamp 1751532440
transform 1 0 24416 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_310
timestamp 1751532440
transform 1 0 36064 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_314
timestamp 1751532423
transform 1 0 36512 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_329
timestamp 1751532440
transform 1 0 38192 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_39_2
timestamp 1751532351
transform 1 0 1568 0 -1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_39_18
timestamp 1751532351
transform 1 0 3360 0 -1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_39_52
timestamp 1751532312
transform 1 0 7168 0 -1 34496
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_60
timestamp 1751532440
transform 1 0 8064 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_62
timestamp 1751532423
transform 1 0 8288 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_153
timestamp 1751532440
transform 1 0 18480 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_182
timestamp 1751532423
transform 1 0 21728 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_212
timestamp 1751532440
transform 1 0 25088 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_241
timestamp 1751532440
transform 1 0 28336 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_243
timestamp 1751532423
transform 1 0 28560 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_277
timestamp 1751532440
transform 1 0 32368 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_279
timestamp 1751532423
transform 1 0 32592 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_309
timestamp 1751532440
transform 1 0 35952 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_313
timestamp 1751532440
transform 1 0 36400 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_317
timestamp 1751532440
transform 1 0 36848 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_40_2
timestamp 1751532246
transform 1 0 1568 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_6
timestamp 1751532423
transform 1 0 2016 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_40_25
timestamp 1751532312
transform 1 0 4144 0 1 34496
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_33
timestamp 1751532440
transform 1 0 5040 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_70
timestamp 1751532440
transform 1 0 9184 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_74
timestamp 1751532440
transform 1 0 9632 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_107
timestamp 1751532440
transform 1 0 13328 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_109
timestamp 1751532423
transform 1 0 13552 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_157
timestamp 1751532440
transform 1 0 18928 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_159
timestamp 1751532423
transform 1 0 19152 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_171
timestamp 1751532440
transform 1 0 20496 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_208
timestamp 1751532440
transform 1 0 24640 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_210
timestamp 1751532423
transform 1 0 24864 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_310
timestamp 1751532440
transform 1 0 36064 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_314
timestamp 1751532423
transform 1 0 36512 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_40_317
timestamp 1751532312
transform 1 0 36848 0 1 34496
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_327
timestamp 1751532440
transform 1 0 37968 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_41_2
timestamp 1751532312
transform 1 0 1568 0 -1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_37
timestamp 1751532440
transform 1 0 5488 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_41
timestamp 1751532440
transform 1 0 5936 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_72
timestamp 1751532440
transform 1 0 9408 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_41_76
timestamp 1751532312
transform 1 0 9856 0 -1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_84
timestamp 1751532423
transform 1 0 10752 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_91
timestamp 1751532423
transform 1 0 11536 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_139
timestamp 1751532423
transform 1 0 16912 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_169
timestamp 1751532440
transform 1 0 20272 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_200
timestamp 1751532440
transform 1 0 23744 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_268
timestamp 1751532440
transform 1 0 31360 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_270
timestamp 1751532423
transform 1 0 31584 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_277
timestamp 1751532440
transform 1 0 32368 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_279
timestamp 1751532423
transform 1 0 32592 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_41_319
timestamp 1751532312
transform 1 0 37072 0 -1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_41_327
timestamp 1751532246
transform 1 0 37968 0 -1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_42_2
timestamp 1751532312
transform 1 0 1568 0 1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_10
timestamp 1751532246
transform 1 0 2464 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_14
timestamp 1751532440
transform 1 0 2912 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_16
timestamp 1751532423
transform 1 0 3136 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_21
timestamp 1751532246
transform 1 0 3696 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_25
timestamp 1751532440
transform 1 0 4144 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_31
timestamp 1751532440
transform 1 0 4816 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_33
timestamp 1751532423
transform 1 0 5040 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_36
timestamp 1751532423
transform 1 0 5376 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_41
timestamp 1751532246
transform 1 0 5936 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_45
timestamp 1751532440
transform 1 0 6384 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_51
timestamp 1751532246
transform 1 0 7056 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_55
timestamp 1751532440
transform 1 0 7504 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_61
timestamp 1751532440
transform 1 0 8176 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_63
timestamp 1751532423
transform 1 0 8400 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_70
timestamp 1751532440
transform 1 0 9184 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_72
timestamp 1751532423
transform 1 0 9408 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_104
timestamp 1751532423
transform 1 0 12992 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_144
timestamp 1751532423
transform 1 0 17472 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_199
timestamp 1751532440
transform 1 0 23632 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_203
timestamp 1751532423
transform 1 0 24080 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_237
timestamp 1751532423
transform 1 0 27888 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_271
timestamp 1751532423
transform 1 0 31696 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_305
timestamp 1751532423
transform 1 0 35504 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_308
timestamp 1751532440
transform 1 0 35840 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_42_312
timestamp 1751532312
transform 1 0 36288 0 1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_320
timestamp 1751532440
transform 1 0 37184 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_322
timestamp 1751532423
transform 1 0 37408 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input1
timestamp 1751534193
transform -1 0 37744 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input2
timestamp 1751534193
transform -1 0 38416 0 1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input3
timestamp 1751534193
transform -1 0 38416 0 -1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input4
timestamp 1751534193
transform -1 0 38416 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input5
timestamp 1751534193
transform -1 0 38416 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input6
timestamp 1751534193
transform -1 0 38416 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input7
timestamp 1751534193
transform -1 0 38416 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input8
timestamp 1751534193
transform -1 0 38416 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input9
timestamp 1751534193
transform -1 0 38416 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input10
timestamp 1751534193
transform -1 0 38416 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input11
timestamp 1751534193
transform -1 0 38416 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input12
timestamp 1751534193
transform -1 0 27888 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input13
timestamp 1751534193
transform -1 0 28896 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input14
timestamp 1751534193
transform -1 0 30576 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input15
timestamp 1751534193
transform 1 0 32032 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input16
timestamp 1751534193
transform 1 0 33488 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input17
timestamp 1751534193
transform 1 0 35840 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input18
timestamp 1751534193
transform 1 0 37072 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input19
timestamp 1751534193
transform -1 0 38416 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output20
timestamp 1751661108
transform 1 0 14224 0 -1 34496
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output21
timestamp 1751661108
transform 1 0 15008 0 1 32928
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output22
timestamp 1751661108
transform 1 0 13776 0 1 36064
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output23
timestamp 1751661108
transform 1 0 17808 0 1 32928
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output24
timestamp 1751661108
transform 1 0 18928 0 -1 34496
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output25
timestamp 1751661108
transform -1 0 20384 0 1 36064
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output26
timestamp 1751661108
transform 1 0 21168 0 1 34496
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output27
timestamp 1751661108
transform 1 0 24416 0 1 36064
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output28
timestamp 1751661108
transform 1 0 25088 0 -1 36064
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output29
timestamp 1751661108
transform -1 0 31024 0 1 36064
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output30
timestamp 1751661108
transform 1 0 27888 0 -1 36064
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output31
timestamp 1751661108
transform 1 0 32032 0 1 36064
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output32
timestamp 1751661108
transform 1 0 27888 0 -1 32928
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output33
timestamp 1751661108
transform 1 0 32928 0 1 26656
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output34
timestamp 1751661108
transform 1 0 32704 0 1 31360
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output35
timestamp 1751661108
transform 1 0 32928 0 -1 36064
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output36
timestamp 1751661108
transform -1 0 35728 0 1 29792
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output37
timestamp 1751661108
transform -1 0 36288 0 -1 29792
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output38
timestamp 1751661108
transform -1 0 36624 0 1 28224
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output39
timestamp 1751661108
transform -1 0 32704 0 1 31360
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output40
timestamp 1751661108
transform 1 0 35616 0 -1 26656
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output41
timestamp 1751661108
transform 1 0 11424 0 -1 34496
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output42
timestamp 1751661108
transform 1 0 9968 0 1 36064
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output43
timestamp 1751661108
transform -1 0 4368 0 1 4704
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output44
timestamp 1751661108
transform 1 0 2352 0 1 3136
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output45
timestamp 1751661108
transform -1 0 6384 0 -1 4704
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output46
timestamp 1751661108
transform 1 0 6384 0 -1 4704
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output47
timestamp 1751661108
transform 1 0 6160 0 1 3136
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output48
timestamp 1751661108
transform 1 0 9744 0 -1 4704
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output49
timestamp 1751661108
transform 1 0 25984 0 1 32928
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output50
timestamp 1751661108
transform 1 0 9968 0 1 3136
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output51
timestamp 1751661108
transform 1 0 14000 0 -1 6272
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output52
timestamp 1751661108
transform 1 0 13776 0 1 3136
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output53
timestamp 1751661108
transform 1 0 17360 0 -1 6272
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output54
timestamp 1751661108
transform 1 0 17584 0 1 3136
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output55
timestamp 1751661108
transform 1 0 20944 0 1 3136
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output56
timestamp 1751661108
transform 1 0 24416 0 1 3136
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output57
timestamp 1751661108
transform 1 0 25088 0 -1 6272
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_0_Left_43 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532504
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_0_Right_0
timestamp 1751532504
transform -1 0 38640 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_1_Left_44
timestamp 1751532504
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_1_Right_1
timestamp 1751532504
transform -1 0 38640 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_2_Left_45
timestamp 1751532504
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_2_Right_2
timestamp 1751532504
transform -1 0 38640 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_3_Left_46
timestamp 1751532504
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_3_Right_3
timestamp 1751532504
transform -1 0 38640 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_4_Left_47
timestamp 1751532504
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_4_Right_4
timestamp 1751532504
transform -1 0 38640 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_5_Left_48
timestamp 1751532504
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_5_Right_5
timestamp 1751532504
transform -1 0 38640 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_6_Left_49
timestamp 1751532504
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_6_Right_6
timestamp 1751532504
transform -1 0 38640 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_7_Left_50
timestamp 1751532504
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_7_Right_7
timestamp 1751532504
transform -1 0 38640 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_8_Left_51
timestamp 1751532504
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_8_Right_8
timestamp 1751532504
transform -1 0 38640 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_9_Left_52
timestamp 1751532504
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_9_Right_9
timestamp 1751532504
transform -1 0 38640 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_10_Left_53
timestamp 1751532504
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_10_Right_10
timestamp 1751532504
transform -1 0 38640 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_11_Left_54
timestamp 1751532504
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_11_Right_11
timestamp 1751532504
transform -1 0 38640 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_12_Left_55
timestamp 1751532504
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_12_Right_12
timestamp 1751532504
transform -1 0 38640 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_13_Left_56
timestamp 1751532504
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_13_Right_13
timestamp 1751532504
transform -1 0 38640 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_14_Left_57
timestamp 1751532504
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_14_Right_14
timestamp 1751532504
transform -1 0 38640 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_15_Left_58
timestamp 1751532504
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_15_Right_15
timestamp 1751532504
transform -1 0 38640 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_16_Left_59
timestamp 1751532504
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_16_Right_16
timestamp 1751532504
transform -1 0 38640 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_17_Left_60
timestamp 1751532504
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_17_Right_17
timestamp 1751532504
transform -1 0 38640 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_18_Left_61
timestamp 1751532504
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_18_Right_18
timestamp 1751532504
transform -1 0 38640 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_19_Left_62
timestamp 1751532504
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_19_Right_19
timestamp 1751532504
transform -1 0 38640 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_20_Left_63
timestamp 1751532504
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_20_Right_20
timestamp 1751532504
transform -1 0 38640 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_21_Left_64
timestamp 1751532504
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_21_Right_21
timestamp 1751532504
transform -1 0 38640 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_22_Left_65
timestamp 1751532504
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_22_Right_22
timestamp 1751532504
transform -1 0 38640 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_23_Left_66
timestamp 1751532504
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_23_Right_23
timestamp 1751532504
transform -1 0 38640 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_24_Left_67
timestamp 1751532504
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_24_Right_24
timestamp 1751532504
transform -1 0 38640 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_25_Left_68
timestamp 1751532504
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_25_Right_25
timestamp 1751532504
transform -1 0 38640 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_26_Left_69
timestamp 1751532504
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_26_Right_26
timestamp 1751532504
transform -1 0 38640 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_27_Left_70
timestamp 1751532504
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_27_Right_27
timestamp 1751532504
transform -1 0 38640 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_28_Left_71
timestamp 1751532504
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_28_Right_28
timestamp 1751532504
transform -1 0 38640 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_29_Left_72
timestamp 1751532504
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_29_Right_29
timestamp 1751532504
transform -1 0 38640 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_30_Left_73
timestamp 1751532504
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_30_Right_30
timestamp 1751532504
transform -1 0 38640 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_31_Left_74
timestamp 1751532504
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_31_Right_31
timestamp 1751532504
transform -1 0 38640 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_32_Left_75
timestamp 1751532504
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_32_Right_32
timestamp 1751532504
transform -1 0 38640 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_33_Left_76
timestamp 1751532504
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_33_Right_33
timestamp 1751532504
transform -1 0 38640 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_34_Left_77
timestamp 1751532504
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_34_Right_34
timestamp 1751532504
transform -1 0 38640 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_35_Left_78
timestamp 1751532504
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_35_Right_35
timestamp 1751532504
transform -1 0 38640 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_36_Left_79
timestamp 1751532504
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_36_Right_36
timestamp 1751532504
transform -1 0 38640 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_37_Left_80
timestamp 1751532504
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_37_Right_37
timestamp 1751532504
transform -1 0 38640 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_38_Left_81
timestamp 1751532504
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_38_Right_38
timestamp 1751532504
transform -1 0 38640 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_39_Left_82
timestamp 1751532504
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_39_Right_39
timestamp 1751532504
transform -1 0 38640 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_40_Left_83
timestamp 1751532504
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_40_Right_40
timestamp 1751532504
transform -1 0 38640 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_41_Left_84
timestamp 1751532504
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_41_Right_41
timestamp 1751532504
transform -1 0 38640 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_42_Left_85
timestamp 1751532504
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_42_Right_42
timestamp 1751532504
transform -1 0 38640 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_86
timestamp 1751532504
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_87
timestamp 1751532504
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_88
timestamp 1751532504
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_89
timestamp 1751532504
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_90
timestamp 1751532504
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_91
timestamp 1751532504
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_92
timestamp 1751532504
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_93
timestamp 1751532504
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_94
timestamp 1751532504
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_95
timestamp 1751532504
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_96
timestamp 1751532504
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_97
timestamp 1751532504
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_98
timestamp 1751532504
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_99
timestamp 1751532504
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_100
timestamp 1751532504
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_101
timestamp 1751532504
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_102
timestamp 1751532504
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_103
timestamp 1751532504
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_104
timestamp 1751532504
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_105
timestamp 1751532504
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_106
timestamp 1751532504
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_107
timestamp 1751532504
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_108
timestamp 1751532504
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_109
timestamp 1751532504
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_110
timestamp 1751532504
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_111
timestamp 1751532504
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_112
timestamp 1751532504
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_113
timestamp 1751532504
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_114
timestamp 1751532504
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_115
timestamp 1751532504
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_116
timestamp 1751532504
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_117
timestamp 1751532504
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_118
timestamp 1751532504
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_119
timestamp 1751532504
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_120
timestamp 1751532504
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_121
timestamp 1751532504
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_122
timestamp 1751532504
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_123
timestamp 1751532504
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_124
timestamp 1751532504
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_125
timestamp 1751532504
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_126
timestamp 1751532504
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_127
timestamp 1751532504
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_128
timestamp 1751532504
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_129
timestamp 1751532504
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_130
timestamp 1751532504
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_131
timestamp 1751532504
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_132
timestamp 1751532504
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_133
timestamp 1751532504
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_134
timestamp 1751532504
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_135
timestamp 1751532504
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_136
timestamp 1751532504
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_137
timestamp 1751532504
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_138
timestamp 1751532504
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_139
timestamp 1751532504
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_140
timestamp 1751532504
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_141
timestamp 1751532504
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_142
timestamp 1751532504
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_143
timestamp 1751532504
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_144
timestamp 1751532504
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_145
timestamp 1751532504
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_146
timestamp 1751532504
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_147
timestamp 1751532504
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_148
timestamp 1751532504
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_149
timestamp 1751532504
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_150
timestamp 1751532504
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_151
timestamp 1751532504
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_152
timestamp 1751532504
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_153
timestamp 1751532504
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_154
timestamp 1751532504
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_155
timestamp 1751532504
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_156
timestamp 1751532504
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_157
timestamp 1751532504
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_158
timestamp 1751532504
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_159
timestamp 1751532504
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_160
timestamp 1751532504
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_161
timestamp 1751532504
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_162
timestamp 1751532504
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_163
timestamp 1751532504
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_164
timestamp 1751532504
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_165
timestamp 1751532504
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_166
timestamp 1751532504
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_167
timestamp 1751532504
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_168
timestamp 1751532504
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_169
timestamp 1751532504
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_170
timestamp 1751532504
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_171
timestamp 1751532504
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_172
timestamp 1751532504
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_173
timestamp 1751532504
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_174
timestamp 1751532504
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_175
timestamp 1751532504
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_176
timestamp 1751532504
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_177
timestamp 1751532504
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_178
timestamp 1751532504
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_179
timestamp 1751532504
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_180
timestamp 1751532504
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_181
timestamp 1751532504
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_182
timestamp 1751532504
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_183
timestamp 1751532504
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_184
timestamp 1751532504
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_185
timestamp 1751532504
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_186
timestamp 1751532504
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_187
timestamp 1751532504
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_188
timestamp 1751532504
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_189
timestamp 1751532504
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_190
timestamp 1751532504
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_191
timestamp 1751532504
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_192
timestamp 1751532504
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_193
timestamp 1751532504
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_194
timestamp 1751532504
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_195
timestamp 1751532504
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_196
timestamp 1751532504
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_197
timestamp 1751532504
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_198
timestamp 1751532504
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_199
timestamp 1751532504
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_200
timestamp 1751532504
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_201
timestamp 1751532504
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_202
timestamp 1751532504
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_203
timestamp 1751532504
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_204
timestamp 1751532504
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_205
timestamp 1751532504
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_206
timestamp 1751532504
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_207
timestamp 1751532504
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_208
timestamp 1751532504
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_209
timestamp 1751532504
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_210
timestamp 1751532504
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_211
timestamp 1751532504
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_212
timestamp 1751532504
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_213
timestamp 1751532504
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_214
timestamp 1751532504
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_215
timestamp 1751532504
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_216
timestamp 1751532504
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_217
timestamp 1751532504
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_218
timestamp 1751532504
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_219
timestamp 1751532504
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_220
timestamp 1751532504
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_221
timestamp 1751532504
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_222
timestamp 1751532504
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_223
timestamp 1751532504
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_224
timestamp 1751532504
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_225
timestamp 1751532504
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_226
timestamp 1751532504
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_227
timestamp 1751532504
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_228
timestamp 1751532504
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_229
timestamp 1751532504
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_230
timestamp 1751532504
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_231
timestamp 1751532504
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_232
timestamp 1751532504
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_233
timestamp 1751532504
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_234
timestamp 1751532504
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_235
timestamp 1751532504
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_236
timestamp 1751532504
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_237
timestamp 1751532504
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_238
timestamp 1751532504
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_239
timestamp 1751532504
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_240
timestamp 1751532504
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_241
timestamp 1751532504
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_242
timestamp 1751532504
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_243
timestamp 1751532504
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_244
timestamp 1751532504
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_245
timestamp 1751532504
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_246
timestamp 1751532504
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_247
timestamp 1751532504
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_248
timestamp 1751532504
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_249
timestamp 1751532504
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_250
timestamp 1751532504
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_251
timestamp 1751532504
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_252
timestamp 1751532504
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_253
timestamp 1751532504
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_254
timestamp 1751532504
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_255
timestamp 1751532504
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_256
timestamp 1751532504
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_257
timestamp 1751532504
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_258
timestamp 1751532504
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_259
timestamp 1751532504
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_260
timestamp 1751532504
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_261
timestamp 1751532504
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_262
timestamp 1751532504
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_263
timestamp 1751532504
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_264
timestamp 1751532504
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_265
timestamp 1751532504
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_266
timestamp 1751532504
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_267
timestamp 1751532504
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_268
timestamp 1751532504
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_269
timestamp 1751532504
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_270
timestamp 1751532504
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_271
timestamp 1751532504
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_272
timestamp 1751532504
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_273
timestamp 1751532504
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_274
timestamp 1751532504
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_275
timestamp 1751532504
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_276
timestamp 1751532504
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_277
timestamp 1751532504
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_278
timestamp 1751532504
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_279
timestamp 1751532504
transform 1 0 5152 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_280
timestamp 1751532504
transform 1 0 8960 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_281
timestamp 1751532504
transform 1 0 12768 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_282
timestamp 1751532504
transform 1 0 16576 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_283
timestamp 1751532504
transform 1 0 20384 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_284
timestamp 1751532504
transform 1 0 24192 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_285
timestamp 1751532504
transform 1 0 28000 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_286
timestamp 1751532504
transform 1 0 31808 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_287
timestamp 1751532504
transform 1 0 35616 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_mc14500_68 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532612
transform 1 0 3248 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_mc14500_69
timestamp 1751532612
transform 1 0 4368 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_mc14500_70
timestamp 1751532612
transform 1 0 5488 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_mc14500_71
timestamp 1751532612
transform 1 0 6608 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_mc14500_72
timestamp 1751532612
transform 1 0 7728 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_mc14500_73
timestamp 1751532612
transform -1 0 8960 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_mc14500_74
timestamp 1751532612
transform -1 0 9968 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_mc14500_75
timestamp 1751532612
transform 1 0 11088 0 -1 36064
box -86 -86 534 870
<< labels >>
flabel metal3 s 39200 31584 40000 31696 0 FreeSans 448 0 0 0 SDI
port 0 nsew signal input
flabel metal3 s 39200 2464 40000 2576 0 FreeSans 448 0 0 0 clk_i
port 1 nsew signal input
flabel metal3 s 39200 37408 40000 37520 0 FreeSans 448 0 0 0 custom_setting
port 2 nsew signal input
flabel metal3 s 39200 8288 40000 8400 0 FreeSans 448 0 0 0 io_in[0]
port 3 nsew signal input
flabel metal3 s 39200 11200 40000 11312 0 FreeSans 448 0 0 0 io_in[1]
port 4 nsew signal input
flabel metal3 s 39200 14112 40000 14224 0 FreeSans 448 0 0 0 io_in[2]
port 5 nsew signal input
flabel metal3 s 39200 17024 40000 17136 0 FreeSans 448 0 0 0 io_in[3]
port 6 nsew signal input
flabel metal3 s 39200 19936 40000 20048 0 FreeSans 448 0 0 0 io_in[4]
port 7 nsew signal input
flabel metal3 s 39200 22848 40000 22960 0 FreeSans 448 0 0 0 io_in[5]
port 8 nsew signal input
flabel metal3 s 39200 25760 40000 25872 0 FreeSans 448 0 0 0 io_in[6]
port 9 nsew signal input
flabel metal3 s 39200 28672 40000 28784 0 FreeSans 448 0 0 0 io_in[7]
port 10 nsew signal input
flabel metal2 s 3136 39200 3248 40000 0 FreeSans 448 90 0 0 io_out[0]
port 11 nsew signal output
flabel metal2 s 14336 39200 14448 40000 0 FreeSans 448 90 0 0 io_out[10]
port 12 nsew signal output
flabel metal2 s 15456 39200 15568 40000 0 FreeSans 448 90 0 0 io_out[11]
port 13 nsew signal output
flabel metal2 s 16576 39200 16688 40000 0 FreeSans 448 90 0 0 io_out[12]
port 14 nsew signal output
flabel metal2 s 17696 39200 17808 40000 0 FreeSans 448 90 0 0 io_out[13]
port 15 nsew signal output
flabel metal2 s 18816 39200 18928 40000 0 FreeSans 448 90 0 0 io_out[14]
port 16 nsew signal output
flabel metal2 s 19936 39200 20048 40000 0 FreeSans 448 90 0 0 io_out[15]
port 17 nsew signal output
flabel metal2 s 21056 39200 21168 40000 0 FreeSans 448 90 0 0 io_out[16]
port 18 nsew signal output
flabel metal2 s 22176 39200 22288 40000 0 FreeSans 448 90 0 0 io_out[17]
port 19 nsew signal output
flabel metal2 s 23296 39200 23408 40000 0 FreeSans 448 90 0 0 io_out[18]
port 20 nsew signal output
flabel metal2 s 24416 39200 24528 40000 0 FreeSans 448 90 0 0 io_out[19]
port 21 nsew signal output
flabel metal2 s 4256 39200 4368 40000 0 FreeSans 448 90 0 0 io_out[1]
port 22 nsew signal output
flabel metal2 s 25536 39200 25648 40000 0 FreeSans 448 90 0 0 io_out[20]
port 23 nsew signal output
flabel metal2 s 26656 39200 26768 40000 0 FreeSans 448 90 0 0 io_out[21]
port 24 nsew signal output
flabel metal2 s 27776 39200 27888 40000 0 FreeSans 448 90 0 0 io_out[22]
port 25 nsew signal output
flabel metal2 s 28896 39200 29008 40000 0 FreeSans 448 90 0 0 io_out[23]
port 26 nsew signal output
flabel metal2 s 30016 39200 30128 40000 0 FreeSans 448 90 0 0 io_out[24]
port 27 nsew signal output
flabel metal2 s 31136 39200 31248 40000 0 FreeSans 448 90 0 0 io_out[25]
port 28 nsew signal output
flabel metal2 s 32256 39200 32368 40000 0 FreeSans 448 90 0 0 io_out[26]
port 29 nsew signal output
flabel metal2 s 33376 39200 33488 40000 0 FreeSans 448 90 0 0 io_out[27]
port 30 nsew signal output
flabel metal2 s 34496 39200 34608 40000 0 FreeSans 448 90 0 0 io_out[28]
port 31 nsew signal output
flabel metal2 s 35616 39200 35728 40000 0 FreeSans 448 90 0 0 io_out[29]
port 32 nsew signal output
flabel metal2 s 5376 39200 5488 40000 0 FreeSans 448 90 0 0 io_out[2]
port 33 nsew signal output
flabel metal2 s 36736 39200 36848 40000 0 FreeSans 448 90 0 0 io_out[30]
port 34 nsew signal output
flabel metal2 s 6496 39200 6608 40000 0 FreeSans 448 90 0 0 io_out[3]
port 35 nsew signal output
flabel metal2 s 7616 39200 7728 40000 0 FreeSans 448 90 0 0 io_out[4]
port 36 nsew signal output
flabel metal2 s 8736 39200 8848 40000 0 FreeSans 448 90 0 0 io_out[5]
port 37 nsew signal output
flabel metal2 s 9856 39200 9968 40000 0 FreeSans 448 90 0 0 io_out[6]
port 38 nsew signal output
flabel metal2 s 10976 39200 11088 40000 0 FreeSans 448 90 0 0 io_out[7]
port 39 nsew signal output
flabel metal2 s 12096 39200 12208 40000 0 FreeSans 448 90 0 0 io_out[8]
port 40 nsew signal output
flabel metal2 s 13216 39200 13328 40000 0 FreeSans 448 90 0 0 io_out[9]
port 41 nsew signal output
flabel metal3 s 39200 5376 40000 5488 0 FreeSans 448 0 0 0 rst_n
port 42 nsew signal input
flabel metal2 s 1120 0 1232 800 0 FreeSans 448 90 0 0 sram_addr[0]
port 43 nsew signal output
flabel metal2 s 2912 0 3024 800 0 FreeSans 448 90 0 0 sram_addr[1]
port 44 nsew signal output
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 sram_addr[2]
port 45 nsew signal output
flabel metal2 s 6496 0 6608 800 0 FreeSans 448 90 0 0 sram_addr[3]
port 46 nsew signal output
flabel metal2 s 8288 0 8400 800 0 FreeSans 448 90 0 0 sram_addr[4]
port 47 nsew signal output
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 sram_addr[5]
port 48 nsew signal output
flabel metal3 s 39200 34496 40000 34608 0 FreeSans 448 0 0 0 sram_gwe
port 49 nsew signal output
flabel metal2 s 11872 0 11984 800 0 FreeSans 448 90 0 0 sram_in[0]
port 50 nsew signal output
flabel metal2 s 13664 0 13776 800 0 FreeSans 448 90 0 0 sram_in[1]
port 51 nsew signal output
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 sram_in[2]
port 52 nsew signal output
flabel metal2 s 17248 0 17360 800 0 FreeSans 448 90 0 0 sram_in[3]
port 53 nsew signal output
flabel metal2 s 19040 0 19152 800 0 FreeSans 448 90 0 0 sram_in[4]
port 54 nsew signal output
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 sram_in[5]
port 55 nsew signal output
flabel metal2 s 22624 0 22736 800 0 FreeSans 448 90 0 0 sram_in[6]
port 56 nsew signal output
flabel metal2 s 24416 0 24528 800 0 FreeSans 448 90 0 0 sram_in[7]
port 57 nsew signal output
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 sram_out[0]
port 58 nsew signal input
flabel metal2 s 28000 0 28112 800 0 FreeSans 448 90 0 0 sram_out[1]
port 59 nsew signal input
flabel metal2 s 29792 0 29904 800 0 FreeSans 448 90 0 0 sram_out[2]
port 60 nsew signal input
flabel metal2 s 31584 0 31696 800 0 FreeSans 448 90 0 0 sram_out[3]
port 61 nsew signal input
flabel metal2 s 33376 0 33488 800 0 FreeSans 448 90 0 0 sram_out[4]
port 62 nsew signal input
flabel metal2 s 35168 0 35280 800 0 FreeSans 448 90 0 0 sram_out[5]
port 63 nsew signal input
flabel metal2 s 36960 0 37072 800 0 FreeSans 448 90 0 0 sram_out[6]
port 64 nsew signal input
flabel metal2 s 38752 0 38864 800 0 FreeSans 448 90 0 0 sram_out[7]
port 65 nsew signal input
flabel metal4 s 5846 3076 6166 36908 0 FreeSans 1280 90 0 0 vdd
port 66 nsew power bidirectional
flabel metal4 s 15170 3076 15490 36908 0 FreeSans 1280 90 0 0 vdd
port 66 nsew power bidirectional
flabel metal4 s 24494 3076 24814 36908 0 FreeSans 1280 90 0 0 vdd
port 66 nsew power bidirectional
flabel metal4 s 33818 3076 34138 36908 0 FreeSans 1280 90 0 0 vdd
port 66 nsew power bidirectional
flabel metal4 s 10508 3076 10828 36908 0 FreeSans 1280 90 0 0 vss
port 67 nsew ground bidirectional
flabel metal4 s 19832 3076 20152 36908 0 FreeSans 1280 90 0 0 vss
port 67 nsew ground bidirectional
flabel metal4 s 29156 3076 29476 36908 0 FreeSans 1280 90 0 0 vss
port 67 nsew ground bidirectional
flabel metal4 s 38480 3076 38800 36908 0 FreeSans 1280 90 0 0 vss
port 67 nsew ground bidirectional
rlabel metal1 19992 36848 19992 36848 0 vdd
rlabel via1 20072 36064 20072 36064 0 vss
rlabel metal2 30184 31864 30184 31864 0 SCLK
rlabel metal2 37688 34048 37688 34048 0 SDI
rlabel metal2 34440 32928 34440 32928 0 SDO
rlabel metal2 29624 15568 29624 15568 0 _0000_
rlabel metal2 25928 12824 25928 12824 0 _0001_
rlabel metal2 17864 18088 17864 18088 0 _0002_
rlabel metal3 36400 30856 36400 30856 0 _0003_
rlabel metal2 35112 26684 35112 26684 0 _0004_
rlabel metal2 37520 19992 37520 19992 0 _0005_
rlabel metal2 35784 21112 35784 21112 0 _0006_
rlabel metal3 35112 32424 35112 32424 0 _0007_
rlabel metal2 30016 28056 30016 28056 0 _0008_
rlabel metal2 33824 34104 33824 34104 0 _0009_
rlabel metal2 32536 33880 32536 33880 0 _0010_
rlabel metal2 22456 13832 22456 13832 0 _0011_
rlabel metal2 15848 10864 15848 10864 0 _0012_
rlabel metal2 11704 9296 11704 9296 0 _0013_
rlabel metal2 14280 7448 14280 7448 0 _0014_
rlabel metal2 11816 6160 11816 6160 0 _0015_
rlabel metal3 12656 4312 12656 4312 0 _0016_
rlabel metal3 15288 5208 15288 5208 0 _0017_
rlabel metal2 18032 6888 18032 6888 0 _0018_
rlabel metal3 18984 8792 18984 8792 0 _0019_
rlabel metal2 19376 4312 19376 4312 0 _0020_
rlabel metal3 23128 4312 23128 4312 0 _0021_
rlabel metal2 22680 7112 22680 7112 0 _0022_
rlabel metal2 25592 5824 25592 5824 0 _0023_
rlabel metal2 27776 4312 27776 4312 0 _0024_
rlabel metal2 30744 4816 30744 4816 0 _0025_
rlabel metal2 33768 4816 33768 4816 0 _0026_
rlabel metal2 36176 5880 36176 5880 0 _0027_
rlabel metal2 36680 8064 36680 8064 0 _0028_
rlabel metal2 34832 10024 34832 10024 0 _0029_
rlabel metal2 23240 10136 23240 10136 0 _0030_
rlabel metal2 25928 10864 25928 10864 0 _0031_
rlabel metal2 31192 10528 31192 10528 0 _0032_
rlabel metal3 30240 12936 30240 12936 0 _0033_
rlabel metal2 34272 15848 34272 15848 0 _0034_
rlabel metal2 37576 12824 37576 12824 0 _0035_
rlabel metal3 34720 16744 34720 16744 0 _0036_
rlabel metal2 34440 17976 34440 17976 0 _0037_
rlabel metal2 25816 35224 25816 35224 0 _0038_
rlabel metal2 27552 34104 27552 34104 0 _0039_
rlabel metal2 26600 28336 26600 28336 0 _0040_
rlabel metal2 28168 13720 28168 13720 0 _0041_
rlabel metal2 15848 13272 15848 13272 0 _0042_
rlabel metal3 16184 22344 16184 22344 0 _0043_
rlabel metal3 31192 34888 31192 34888 0 _0044_
rlabel metal3 31472 33992 31472 33992 0 _0045_
rlabel metal2 24360 13272 24360 13272 0 _0046_
rlabel metal2 9128 21672 9128 21672 0 _0047_
rlabel metal2 8792 23352 8792 23352 0 _0048_
rlabel metal2 5432 27608 5432 27608 0 _0049_
rlabel metal2 3808 30408 3808 30408 0 _0050_
rlabel metal2 3192 32200 3192 32200 0 _0051_
rlabel metal2 3080 28952 3080 28952 0 _0052_
rlabel metal2 2856 24976 2856 24976 0 _0053_
rlabel metal2 2856 21224 2856 21224 0 _0054_
rlabel metal2 4760 19656 4760 19656 0 _0055_
rlabel metal2 6608 18424 6608 18424 0 _0056_
rlabel metal3 8680 17864 8680 17864 0 _0057_
rlabel metal2 10864 17640 10864 17640 0 _0058_
rlabel metal2 14504 16520 14504 16520 0 _0059_
rlabel metal2 15288 18928 15288 18928 0 _0060_
rlabel metal2 12600 20356 12600 20356 0 _0061_
rlabel metal2 12376 23800 12376 23800 0 _0062_
rlabel metal2 9912 27384 9912 27384 0 _0063_
rlabel metal2 5992 34608 5992 34608 0 _0064_
rlabel metal2 2968 35336 2968 35336 0 _0065_
rlabel metal2 10920 34608 10920 34608 0 _0066_
rlabel metal2 8792 35336 8792 35336 0 _0067_
rlabel metal2 13104 32760 13104 32760 0 _0068_
rlabel metal2 16744 35616 16744 35616 0 _0069_
rlabel metal2 15512 35112 15512 35112 0 _0070_
rlabel metal2 18032 30408 18032 30408 0 _0071_
rlabel metal2 22736 33544 22736 33544 0 _0072_
rlabel metal2 24360 35448 24360 35448 0 _0073_
rlabel metal2 20776 23632 20776 23632 0 _0074_
rlabel metal3 21560 24584 21560 24584 0 _0075_
rlabel metal3 24192 29624 24192 29624 0 _0076_
rlabel metal2 23016 32872 23016 32872 0 _0077_
rlabel metal2 26824 31080 26824 31080 0 _0078_
rlabel metal2 12600 13216 12600 13216 0 _0079_
rlabel metal2 7952 13944 7952 13944 0 _0080_
rlabel metal2 6608 11368 6608 11368 0 _0081_
rlabel metal2 5992 9520 5992 9520 0 _0082_
rlabel metal2 6664 6160 6664 6160 0 _0083_
rlabel metal3 9632 5208 9632 5208 0 _0084_
rlabel metal3 20664 16072 20664 16072 0 _0085_
rlabel metal2 20776 18368 20776 18368 0 _0086_
rlabel metal2 21392 14728 21392 14728 0 _0087_
rlabel metal2 20804 14728 20804 14728 0 _0088_
rlabel metal2 20664 18956 20664 18956 0 _0089_
rlabel metal2 29960 19936 29960 19936 0 _0090_
rlabel metal3 21504 15064 21504 15064 0 _0091_
rlabel metal3 21981 14952 21981 14952 0 _0092_
rlabel metal2 21560 19992 21560 19992 0 _0093_
rlabel metal2 24472 20328 24472 20328 0 _0094_
rlabel metal2 22250 16464 22250 16464 0 _0095_
rlabel metal2 30296 18984 30296 18984 0 _0096_
rlabel metal3 30604 19992 30604 19992 0 _0097_
rlabel metal2 31892 19880 31892 19880 0 _0098_
rlabel metal3 22456 21560 22456 21560 0 _0099_
rlabel metal2 22344 17080 22344 17080 0 _0100_
rlabel metal2 19936 20132 19936 20132 0 _0101_
rlabel metal3 23968 19768 23968 19768 0 _0102_
rlabel metal2 23912 17472 23912 17472 0 _0103_
rlabel metal2 21000 16996 21000 16996 0 _0104_
rlabel metal2 20440 17164 20440 17164 0 _0105_
rlabel metal2 23016 19356 23016 19356 0 _0106_
rlabel metal2 24808 18704 24808 18704 0 _0107_
rlabel metal2 24248 17584 24248 17584 0 _0108_
rlabel metal3 23100 18536 23100 18536 0 _0109_
rlabel metal2 22357 14616 22357 14616 0 _0110_
rlabel metal3 28952 18424 28952 18424 0 _0111_
rlabel metal2 25928 18508 25928 18508 0 _0112_
rlabel metal2 25032 19656 25032 19656 0 _0113_
rlabel metal3 19712 23128 19712 23128 0 _0114_
rlabel metal2 15120 14000 15120 14000 0 _0115_
rlabel metal2 14728 12544 14728 12544 0 _0116_
rlabel metal2 37688 30072 37688 30072 0 _0117_
rlabel metal2 32536 24864 32536 24864 0 _0118_
rlabel metal3 31752 25480 31752 25480 0 _0119_
rlabel metal3 36120 24696 36120 24696 0 _0120_
rlabel metal2 33880 25396 33880 25396 0 _0121_
rlabel metal2 23464 22736 23464 22736 0 _0122_
rlabel metal3 24724 22344 24724 22344 0 _0123_
rlabel metal3 21084 19432 21084 19432 0 _0124_
rlabel metal2 21364 19432 21364 19432 0 _0125_
rlabel metal3 23968 20776 23968 20776 0 _0126_
rlabel metal2 26488 20272 26488 20272 0 _0127_
rlabel metal2 26376 18228 26376 18228 0 _0128_
rlabel via1 26600 21579 26600 21579 0 _0129_
rlabel metal2 30464 24696 30464 24696 0 _0130_
rlabel metal2 31640 24774 31640 24774 0 _0131_
rlabel metal2 31472 26488 31472 26488 0 _0132_
rlabel metal2 36344 30520 36344 30520 0 _0133_
rlabel metal3 35588 31864 35588 31864 0 _0134_
rlabel metal2 34104 22456 34104 22456 0 _0135_
rlabel metal3 31808 24808 31808 24808 0 _0136_
rlabel metal2 33768 24976 33768 24976 0 _0137_
rlabel metal2 33376 21728 33376 21728 0 _0138_
rlabel metal3 35000 23128 35000 23128 0 _0139_
rlabel metal2 31864 22176 31864 22176 0 _0140_
rlabel metal2 36008 24192 36008 24192 0 _0141_
rlabel metal2 31080 22624 31080 22624 0 _0142_
rlabel metal2 32032 25480 32032 25480 0 _0143_
rlabel metal3 32256 24584 32256 24584 0 _0144_
rlabel metal3 32816 22456 32816 22456 0 _0145_
rlabel metal2 33992 21896 33992 21896 0 _0146_
rlabel metal2 33488 20300 33488 20300 0 _0147_
rlabel metal2 14168 18032 14168 18032 0 _0148_
rlabel metal3 20496 21000 20496 21000 0 _0149_
rlabel metal2 32032 23912 32032 23912 0 _0150_
rlabel metal2 31752 26208 31752 26208 0 _0151_
rlabel metal2 31976 20776 31976 20776 0 _0152_
rlabel metal2 34234 20216 34234 20216 0 _0153_
rlabel metal2 29288 29484 29288 29484 0 _0154_
rlabel metal2 31024 28056 31024 28056 0 _0155_
rlabel metal2 26824 21616 26824 21616 0 _0156_
rlabel metal3 31136 26712 31136 26712 0 _0157_
rlabel metal3 30660 26376 30660 26376 0 _0158_
rlabel metal2 30408 28168 30408 28168 0 _0159_
rlabel metal2 33264 28196 33264 28196 0 _0160_
rlabel metal2 33040 27832 33040 27832 0 _0161_
rlabel metal2 33833 27608 33833 27608 0 _0162_
rlabel metal2 31864 25508 31864 25508 0 _0163_
rlabel metal2 33190 31136 33190 31136 0 _0164_
rlabel metal2 37352 31024 37352 31024 0 _0165_
rlabel metal2 15036 8344 15036 8344 0 _0166_
rlabel metal2 30856 23436 30856 23436 0 _0167_
rlabel metal2 30576 26040 30576 26040 0 _0168_
rlabel metal2 31145 28840 31145 28840 0 _0169_
rlabel metal3 31668 32648 31668 32648 0 _0170_
rlabel metal3 33544 30184 33544 30184 0 _0171_
rlabel metal3 31808 27272 31808 27272 0 _0172_
rlabel metal2 32732 27272 32732 27272 0 _0173_
rlabel metal3 36353 30072 36353 30072 0 _0174_
rlabel metal2 25760 16940 25760 16940 0 _0175_
rlabel metal2 25760 17388 25760 17388 0 _0176_
rlabel metal2 25592 16912 25592 16912 0 _0177_
rlabel metal3 26180 17640 26180 17640 0 _0178_
rlabel metal2 25928 17864 25928 17864 0 _0179_
rlabel metal3 21700 17640 21700 17640 0 _0180_
rlabel metal2 20720 16184 20720 16184 0 _0181_
rlabel metal3 24285 16072 24285 16072 0 _0182_
rlabel metal2 24808 15512 24808 15512 0 _0183_
rlabel metal2 25816 14056 25816 14056 0 _0184_
rlabel metal2 36335 23240 36335 23240 0 _0185_
rlabel metal2 35952 18788 35952 18788 0 _0186_
rlabel metal2 35672 23968 35672 23968 0 _0187_
rlabel metal3 36876 23912 36876 23912 0 _0188_
rlabel metal2 37352 27384 37352 27384 0 _0189_
rlabel metal2 38033 21000 38033 21000 0 _0190_
rlabel metal2 37352 26180 37352 26180 0 _0191_
rlabel metal2 37744 28616 37744 28616 0 _0192_
rlabel metal2 37184 28924 37184 28924 0 _0193_
rlabel metal2 37772 26152 37772 26152 0 _0194_
rlabel metal2 37856 24220 37856 24220 0 _0195_
rlabel metal2 25928 14560 25928 14560 0 _0196_
rlabel metal2 19656 16548 19656 16548 0 _0197_
rlabel metal2 20776 16940 20776 16940 0 _0198_
rlabel metal3 23660 16856 23660 16856 0 _0199_
rlabel metal3 27468 16856 27468 16856 0 _0200_
rlabel metal2 28952 17528 28952 17528 0 _0201_
rlabel metal2 29064 16380 29064 16380 0 _0202_
rlabel metal2 30408 16111 30408 16111 0 _0203_
rlabel metal2 27944 16744 27944 16744 0 _0204_
rlabel metal3 29176 16184 29176 16184 0 _0205_
rlabel metal2 22568 11592 22568 11592 0 _0206_
rlabel metal2 22484 13160 22484 13160 0 _0207_
rlabel metal3 23529 13720 23529 13720 0 _0208_
rlabel metal3 26852 13944 26852 13944 0 _0209_
rlabel metal2 29960 17752 29960 17752 0 _0210_
rlabel metal2 29512 16389 29512 16389 0 _0211_
rlabel metal2 29356 16279 29356 16279 0 _0212_
rlabel metal2 22456 19320 22456 19320 0 _0213_
rlabel metal2 7672 12208 7672 12208 0 _0214_
rlabel metal3 12544 12264 12544 12264 0 _0215_
rlabel metal3 11256 11368 11256 11368 0 _0216_
rlabel metal2 31416 22848 31416 22848 0 _0217_
rlabel metal3 27888 21560 27888 21560 0 _0218_
rlabel metal2 14392 19572 14392 19572 0 _0219_
rlabel metal2 14672 23912 14672 23912 0 _0220_
rlabel metal2 15008 23688 15008 23688 0 _0221_
rlabel metal2 13832 13440 13832 13440 0 _0222_
rlabel metal2 9520 12712 9520 12712 0 _0223_
rlabel metal3 13449 11368 13449 11368 0 _0224_
rlabel metal2 14392 10920 14392 10920 0 _0225_
rlabel metal3 13384 7448 13384 7448 0 _0226_
rlabel metal2 9744 10444 9744 10444 0 _0227_
rlabel metal3 11153 10024 11153 10024 0 _0228_
rlabel metal2 11508 8456 11508 8456 0 _0229_
rlabel metal2 25592 22792 25592 22792 0 _0230_
rlabel metal2 28168 22120 28168 22120 0 _0231_
rlabel metal2 20496 9744 20496 9744 0 _0232_
rlabel metal2 14504 6328 14504 6328 0 _0233_
rlabel metal2 13711 8456 13711 8456 0 _0234_
rlabel metal2 12824 9352 12824 9352 0 _0235_
rlabel metal2 10714 6048 10714 6048 0 _0236_
rlabel metal2 11200 6664 11200 6664 0 _0237_
rlabel metal2 13496 4872 13496 4872 0 _0238_
rlabel metal2 13188 3752 13188 3752 0 _0239_
rlabel metal2 21784 7448 21784 7448 0 _0240_
rlabel metal2 20328 6160 20328 6160 0 _0241_
rlabel metal3 17257 4312 17257 4312 0 _0242_
rlabel metal3 16436 4424 16436 4424 0 _0243_
rlabel metal2 21504 7448 21504 7448 0 _0244_
rlabel metal3 16063 6888 16063 6888 0 _0245_
rlabel metal2 16520 6944 16520 6944 0 _0246_
rlabel metal3 20057 6664 20057 6664 0 _0247_
rlabel metal2 20636 6664 20636 6664 0 _0248_
rlabel metal2 20440 6496 20440 6496 0 _0249_
rlabel metal2 20888 5376 20888 5376 0 _0250_
rlabel metal2 24136 5824 24136 5824 0 _0251_
rlabel metal2 22904 5768 22904 5768 0 _0252_
rlabel metal3 23436 5096 23436 5096 0 _0253_
rlabel metal2 31192 15736 31192 15736 0 _0254_
rlabel metal2 27048 7924 27048 7924 0 _0255_
rlabel metal2 26208 7644 26208 7644 0 _0256_
rlabel metal2 30044 19432 30044 19432 0 _0257_
rlabel metal2 30632 21336 30632 21336 0 _0258_
rlabel metal2 31696 19320 31696 19320 0 _0259_
rlabel metal2 29064 5824 29064 5824 0 _0260_
rlabel metal2 25462 7616 25462 7616 0 _0261_
rlabel metal3 23464 6664 23464 6664 0 _0262_
rlabel metal2 28896 5964 28896 5964 0 _0263_
rlabel metal3 26255 5880 26255 5880 0 _0264_
rlabel metal2 24668 5992 24668 5992 0 _0265_
rlabel metal2 29494 6048 29494 6048 0 _0266_
rlabel metal2 26264 4592 26264 4592 0 _0267_
rlabel metal2 26628 4424 26628 4424 0 _0268_
rlabel metal2 30744 6608 30744 6608 0 _0269_
rlabel metal2 30912 6076 30912 6076 0 _0270_
rlabel metal2 31658 6048 31658 6048 0 _0271_
rlabel metal2 31864 5432 31864 5432 0 _0272_
rlabel metal2 34104 5768 34104 5768 0 _0273_
rlabel metal2 33190 6048 33190 6048 0 _0274_
rlabel metal2 33320 7728 33320 7728 0 _0275_
rlabel metal2 32200 6216 32200 6216 0 _0276_
rlabel metal2 32928 4312 32928 4312 0 _0277_
rlabel via1 36017 4424 36017 4424 0 _0278_
rlabel metal2 34888 5936 34888 5936 0 _0279_
rlabel metal2 35140 5992 35140 5992 0 _0280_
rlabel metal2 35242 7616 35242 7616 0 _0281_
rlabel metal2 34440 8288 34440 8288 0 _0282_
rlabel metal2 35560 7784 35560 7784 0 _0283_
rlabel metal2 26488 8680 26488 8680 0 _0284_
rlabel via1 36017 8344 36017 8344 0 _0285_
rlabel metal3 35401 9800 35401 9800 0 _0286_
rlabel metal2 33292 9800 33292 9800 0 _0287_
rlabel metal2 29120 23128 29120 23128 0 _0288_
rlabel metal3 28840 23912 28840 23912 0 _0289_
rlabel metal2 31080 19740 31080 19740 0 _0290_
rlabel metal2 26600 9436 26600 9436 0 _0291_
rlabel metal2 26656 10052 26656 10052 0 _0292_
rlabel metal2 30968 20160 30968 20160 0 _0293_
rlabel metal2 30296 19712 30296 19712 0 _0294_
rlabel metal2 32872 16464 32872 16464 0 _0295_
rlabel metal3 26852 9688 26852 9688 0 _0296_
rlabel metal2 26264 8792 26264 8792 0 _0297_
rlabel metal2 26096 8372 26096 8372 0 _0298_
rlabel metal2 27048 9324 27048 9324 0 _0299_
rlabel metal2 27608 9184 27608 9184 0 _0300_
rlabel metal2 27328 9352 27328 9352 0 _0301_
rlabel metal3 29195 9016 29195 9016 0 _0302_
rlabel metal2 29559 9128 29559 9128 0 _0303_
rlabel metal2 29596 10696 29596 10696 0 _0304_
rlabel metal2 6104 23464 6104 23464 0 _0305_
rlabel metal2 15736 14840 15736 14840 0 _0306_
rlabel metal2 30874 10976 30874 10976 0 _0307_
rlabel via1 32097 12264 32097 12264 0 _0308_
rlabel metal2 29960 13216 29960 13216 0 _0309_
rlabel metal3 36568 15400 36568 15400 0 _0310_
rlabel metal3 34225 12824 34225 12824 0 _0311_
rlabel metal2 33880 15624 33880 15624 0 _0312_
rlabel metal2 34897 15064 34897 15064 0 _0313_
rlabel metal2 34496 16072 34496 16072 0 _0314_
rlabel metal3 36381 12936 36381 12936 0 _0315_
rlabel metal2 36120 12880 36120 12880 0 _0316_
rlabel metal2 36400 13328 36400 13328 0 _0317_
rlabel metal2 36326 14000 36326 14000 0 _0318_
rlabel metal3 36736 16072 36736 16072 0 _0319_
rlabel metal3 35924 16296 35924 16296 0 _0320_
rlabel metal2 6888 23184 6888 23184 0 _0321_
rlabel metal2 35318 15568 35318 15568 0 _0322_
rlabel via1 35103 16296 35103 16296 0 _0323_
rlabel metal3 34636 18424 34636 18424 0 _0324_
rlabel metal3 25676 32536 25676 32536 0 _0325_
rlabel metal3 21000 26432 21000 26432 0 _0326_
rlabel metal2 23184 32844 23184 32844 0 _0327_
rlabel metal2 25144 34720 25144 34720 0 _0328_
rlabel metal3 23743 33320 23743 33320 0 _0329_
rlabel metal2 25704 34384 25704 34384 0 _0330_
rlabel metal3 11424 25480 11424 25480 0 _0331_
rlabel metal2 16408 25872 16408 25872 0 _0332_
rlabel metal3 15204 27048 15204 27048 0 _0333_
rlabel metal2 24808 28672 24808 28672 0 _0334_
rlabel metal3 26488 27776 26488 27776 0 _0335_
rlabel metal2 20328 30464 20328 30464 0 _0336_
rlabel metal2 22680 31360 22680 31360 0 _0337_
rlabel metal2 16744 32592 16744 32592 0 _0338_
rlabel metal2 16520 32431 16520 32431 0 _0339_
rlabel metal2 18760 33152 18760 33152 0 _0340_
rlabel metal2 20328 31808 20328 31808 0 _0341_
rlabel metal2 22344 31248 22344 31248 0 _0342_
rlabel metal2 24920 29064 24920 29064 0 _0343_
rlabel metal2 25611 27916 25611 27916 0 _0344_
rlabel metal3 25760 27832 25760 27832 0 _0345_
rlabel metal2 25368 24304 25368 24304 0 _0346_
rlabel metal2 25172 25704 25172 25704 0 _0347_
rlabel metal2 19544 24780 19544 24780 0 _0348_
rlabel metal2 18872 18928 18872 18928 0 _0349_
rlabel metal2 19656 20664 19656 20664 0 _0350_
rlabel metal3 24472 26600 24472 26600 0 _0351_
rlabel metal2 26600 26684 26600 26684 0 _0352_
rlabel metal2 25256 26572 25256 26572 0 _0353_
rlabel metal2 25984 26628 25984 26628 0 _0354_
rlabel metal2 26824 27552 26824 27552 0 _0355_
rlabel metal2 27692 27832 27692 27832 0 _0356_
rlabel metal2 27496 15512 27496 15512 0 _0357_
rlabel metal2 28410 14784 28410 14784 0 _0358_
rlabel metal2 11088 7728 11088 7728 0 _0359_
rlabel metal2 16240 12488 16240 12488 0 _0360_
rlabel metal2 14168 23968 14168 23968 0 _0361_
rlabel metal2 26376 22904 26376 22904 0 _0362_
rlabel metal2 14504 21616 14504 21616 0 _0363_
rlabel metal2 4984 24304 4984 24304 0 _0364_
rlabel metal2 6664 24948 6664 24948 0 _0365_
rlabel metal2 14616 23464 14616 23464 0 _0366_
rlabel metal2 14056 22624 14056 22624 0 _0367_
rlabel metal2 27832 22176 27832 22176 0 _0368_
rlabel metal3 29652 21448 29652 21448 0 _0369_
rlabel metal3 29503 33432 29503 33432 0 _0370_
rlabel metal3 28812 34888 28812 34888 0 _0371_
rlabel metal2 27048 24024 27048 24024 0 _0372_
rlabel metal2 27944 25452 27944 25452 0 _0373_
rlabel metal2 29288 31024 29288 31024 0 _0374_
rlabel metal2 29568 30912 29568 30912 0 _0375_
rlabel metal2 26600 14812 26600 14812 0 _0376_
rlabel metal2 25704 14056 25704 14056 0 _0377_
rlabel metal2 8232 22624 8232 22624 0 _0378_
rlabel metal2 8232 21056 8232 21056 0 _0379_
rlabel metal2 7112 23800 7112 23800 0 _0380_
rlabel metal3 6916 23128 6916 23128 0 _0381_
rlabel metal2 4984 25368 4984 25368 0 _0382_
rlabel metal2 5591 25480 5591 25480 0 _0383_
rlabel metal2 4676 25704 4676 25704 0 _0384_
rlabel metal3 3528 26264 3528 26264 0 _0385_
rlabel metal2 2650 30240 2650 30240 0 _0386_
rlabel metal2 4928 30184 4928 30184 0 _0387_
rlabel metal2 6104 30912 6104 30912 0 _0388_
rlabel metal2 6608 31248 6608 31248 0 _0389_
rlabel metal2 3528 28112 3528 28112 0 _0390_
rlabel metal2 2996 27944 2996 27944 0 _0391_
rlabel metal3 4816 23352 4816 23352 0 _0392_
rlabel metal2 5096 24808 5096 24808 0 _0393_
rlabel metal3 4788 24808 4788 24808 0 _0394_
rlabel metal3 5152 21672 5152 21672 0 _0395_
rlabel metal2 5302 21728 5302 21728 0 _0396_
rlabel metal3 2296 20776 2296 20776 0 _0397_
rlabel metal3 5591 20664 5591 20664 0 _0398_
rlabel metal2 3304 19488 3304 19488 0 _0399_
rlabel metal2 5479 20776 5479 20776 0 _0400_
rlabel metal2 4704 20412 4704 20412 0 _0401_
rlabel metal2 11536 24304 11536 24304 0 _0402_
rlabel metal3 10416 18424 10416 18424 0 _0403_
rlabel metal2 8232 19096 8232 19096 0 _0404_
rlabel metal2 9688 17920 9688 17920 0 _0405_
rlabel metal2 14504 21056 14504 21056 0 _0406_
rlabel metal2 11032 18312 11032 18312 0 _0407_
rlabel metal2 9912 17360 9912 17360 0 _0408_
rlabel metal2 13290 17024 13290 17024 0 _0409_
rlabel metal2 13384 16464 13384 16464 0 _0410_
rlabel metal2 13160 18760 13160 18760 0 _0411_
rlabel metal3 13636 18424 13636 18424 0 _0412_
rlabel metal3 10304 23352 10304 23352 0 _0413_
rlabel metal3 12591 21000 12591 21000 0 _0414_
rlabel metal2 11144 21056 11144 21056 0 _0415_
rlabel metal2 12152 23072 12152 23072 0 _0416_
rlabel metal2 12460 22568 12460 22568 0 _0417_
rlabel metal2 9744 28336 9744 28336 0 _0418_
rlabel metal2 10752 25872 10752 25872 0 _0419_
rlabel metal2 10472 26320 10472 26320 0 _0420_
rlabel metal2 17808 27832 17808 27832 0 _0421_
rlabel metal2 17528 27552 17528 27552 0 _0422_
rlabel metal2 11928 28056 11928 28056 0 _0423_
rlabel metal2 11256 28840 11256 28840 0 _0424_
rlabel metal2 10248 26824 10248 26824 0 _0425_
rlabel metal2 10192 28000 10192 28000 0 _0426_
rlabel metal2 7672 28364 7672 28364 0 _0427_
rlabel metal3 7784 31640 7784 31640 0 _0428_
rlabel metal2 8801 27944 8801 27944 0 _0429_
rlabel metal3 9520 29176 9520 29176 0 _0430_
rlabel via2 8904 28602 8904 28602 0 _0431_
rlabel metal2 8428 28840 8428 28840 0 _0432_
rlabel metal2 8148 29512 8148 29512 0 _0433_
rlabel metal2 9688 29260 9688 29260 0 _0434_
rlabel metal2 7224 29512 7224 29512 0 _0435_
rlabel via2 9016 30170 9016 30170 0 _0436_
rlabel metal2 13048 28728 13048 28728 0 _0437_
rlabel metal2 8792 30100 8792 30100 0 _0438_
rlabel metal2 8288 30688 8288 30688 0 _0439_
rlabel metal2 8064 31304 8064 31304 0 _0440_
rlabel metal2 9464 33544 9464 33544 0 _0441_
rlabel metal2 11144 32592 11144 32592 0 _0442_
rlabel metal2 14616 31528 14616 31528 0 _0443_
rlabel metal2 7448 31220 7448 31220 0 _0444_
rlabel via2 10584 31738 10584 31738 0 _0445_
rlabel metal2 9688 31080 9688 31080 0 _0446_
rlabel metal2 9856 32144 9856 32144 0 _0447_
rlabel metal3 9044 34104 9044 34104 0 _0448_
rlabel metal2 22120 31696 22120 31696 0 _0449_
rlabel metal3 7924 32536 7924 32536 0 _0450_
rlabel metal3 10332 32312 10332 32312 0 _0451_
rlabel metal2 8624 31836 8624 31836 0 _0452_
rlabel metal2 9370 32032 9370 32032 0 _0453_
rlabel metal2 11256 29792 11256 29792 0 _0454_
rlabel metal2 10136 32326 10136 32326 0 _0455_
rlabel metal2 9632 32704 9632 32704 0 _0456_
rlabel metal2 9100 33544 9100 33544 0 _0457_
rlabel metal2 11256 32396 11256 32396 0 _0458_
rlabel metal3 13552 31752 13552 31752 0 _0459_
rlabel metal2 12432 31164 12432 31164 0 _0460_
rlabel metal2 11686 31136 11686 31136 0 _0461_
rlabel metal3 12908 30184 12908 30184 0 _0462_
rlabel metal2 13832 31668 13832 31668 0 _0463_
rlabel metal2 14308 31976 14308 31976 0 _0464_
rlabel metal2 13944 32536 13944 32536 0 _0465_
rlabel metal2 15176 30240 15176 30240 0 _0466_
rlabel metal2 16632 31002 16632 31002 0 _0467_
rlabel metal2 17864 33843 17864 33843 0 _0468_
rlabel metal2 15736 31276 15736 31276 0 _0469_
rlabel metal2 16240 31080 16240 31080 0 _0470_
rlabel metal3 16856 32424 16856 32424 0 _0471_
rlabel metal2 17416 35896 17416 35896 0 _0472_
rlabel metal3 21504 32648 21504 32648 0 _0473_
rlabel metal2 16800 30576 16800 30576 0 _0474_
rlabel metal2 16408 32144 16408 32144 0 _0475_
rlabel metal2 15568 31360 15568 31360 0 _0476_
rlabel metal2 13897 29512 13897 29512 0 _0477_
rlabel metal2 14728 30926 14728 30926 0 _0478_
rlabel metal2 15232 31248 15232 31248 0 _0479_
rlabel metal2 14364 33544 14364 33544 0 _0480_
rlabel metal2 16688 26488 16688 26488 0 _0481_
rlabel metal2 17752 30268 17752 30268 0 _0482_
rlabel metal3 17024 28616 17024 28616 0 _0483_
rlabel metal2 14784 27244 14784 27244 0 _0484_
rlabel metal2 16744 27552 16744 27552 0 _0485_
rlabel metal2 16464 28056 16464 28056 0 _0486_
rlabel metal2 16940 28840 16940 28840 0 _0487_
rlabel metal2 21336 33236 21336 33236 0 _0488_
rlabel metal3 20300 32536 20300 32536 0 _0489_
rlabel metal2 21112 32480 21112 32480 0 _0490_
rlabel metal2 9632 20132 9632 20132 0 _0491_
rlabel metal2 19152 28700 19152 28700 0 _0492_
rlabel metal2 20001 28840 20001 28840 0 _0493_
rlabel metal2 21784 32536 21784 32536 0 _0494_
rlabel metal2 21980 32312 21980 32312 0 _0495_
rlabel metal2 18872 28112 18872 28112 0 _0496_
rlabel metal2 19432 28448 19432 28448 0 _0497_
rlabel metal3 15652 27048 15652 27048 0 _0498_
rlabel metal3 17537 27048 17537 27048 0 _0499_
rlabel metal2 18592 27440 18592 27440 0 _0500_
rlabel metal3 19124 29512 19124 29512 0 _0501_
rlabel metal2 19544 25704 19544 25704 0 _0502_
rlabel metal2 17696 24276 17696 24276 0 _0503_
rlabel metal3 18368 23912 18368 23912 0 _0504_
rlabel via1 18433 24136 18433 24136 0 _0505_
rlabel metal2 18788 23240 18788 23240 0 _0506_
rlabel metal2 25032 29232 25032 29232 0 _0507_
rlabel metal2 18872 25172 18872 25172 0 _0508_
rlabel metal2 20496 23128 20496 23128 0 _0509_
rlabel metal2 19040 24276 19040 24276 0 _0510_
rlabel metal2 20552 25424 20552 25424 0 _0511_
rlabel metal2 18368 23408 18368 23408 0 _0512_
rlabel metal2 19628 24136 19628 24136 0 _0513_
rlabel metal2 20020 24136 20020 24136 0 _0514_
rlabel metal3 20020 25704 20020 25704 0 _0515_
rlabel metal2 20104 24836 20104 24836 0 _0516_
rlabel metal2 20524 24696 20524 24696 0 _0517_
rlabel metal2 22904 29232 22904 29232 0 _0518_
rlabel metal2 21560 27776 21560 27776 0 _0519_
rlabel metal2 21672 27972 21672 27972 0 _0520_
rlabel metal2 21336 26740 21336 26740 0 _0521_
rlabel metal2 18368 22064 18368 22064 0 _0522_
rlabel metal3 21980 29400 21980 29400 0 _0523_
rlabel metal2 19600 26460 19600 26460 0 _0524_
rlabel metal2 20449 26376 20449 26376 0 _0525_
rlabel metal2 21336 27384 21336 27384 0 _0526_
rlabel metal3 22876 28840 22876 28840 0 _0527_
rlabel metal2 15232 25088 15232 25088 0 _0528_
rlabel metal2 23352 31640 23352 31640 0 _0529_
rlabel metal2 15540 30184 15540 30184 0 _0530_
rlabel metal2 16314 30408 16314 30408 0 _0531_
rlabel metal2 21756 31080 21756 31080 0 _0532_
rlabel metal2 22204 30408 22204 30408 0 _0533_
rlabel metal2 22624 32564 22624 32564 0 _0534_
rlabel metal2 15960 25900 15960 25900 0 _0535_
rlabel metal2 24892 21000 24892 21000 0 _0536_
rlabel metal3 25228 27048 25228 27048 0 _0537_
rlabel metal2 25928 30688 25928 30688 0 _0538_
rlabel metal2 25704 30408 25704 30408 0 _0539_
rlabel metal2 25704 32158 25704 32158 0 _0540_
rlabel metal2 8344 9856 8344 9856 0 _0541_
rlabel metal3 13104 12152 13104 12152 0 _0542_
rlabel metal2 11350 12096 11350 12096 0 _0543_
rlabel metal2 11144 13832 11144 13832 0 _0544_
rlabel metal2 10528 13412 10528 13412 0 _0545_
rlabel metal2 8904 13216 8904 13216 0 _0546_
rlabel metal2 8624 13440 8624 13440 0 _0547_
rlabel metal2 7336 7896 7336 7896 0 _0548_
rlabel metal3 8848 12152 8848 12152 0 _0549_
rlabel metal2 8008 7980 8008 7980 0 _0550_
rlabel metal3 9081 11368 9081 11368 0 _0551_
rlabel metal2 8008 10920 8008 10920 0 _0552_
rlabel metal2 8960 9240 8960 9240 0 _0553_
rlabel metal2 8120 9352 8120 9352 0 _0554_
rlabel metal2 7476 9016 7476 9016 0 _0555_
rlabel metal2 7728 7560 7728 7560 0 _0556_
rlabel metal2 9352 8288 9352 8288 0 _0557_
rlabel metal2 8344 7112 8344 7112 0 _0558_
rlabel metal3 9072 7448 9072 7448 0 _0559_
rlabel metal3 9809 6664 9809 6664 0 _0560_
rlabel metal2 10276 6664 10276 6664 0 _0561_
rlabel metal2 24248 5460 24248 5460 0 clk_i
rlabel metal2 22008 11144 22008 11144 0 clknet_0_clk_i
rlabel metal2 5712 5880 5712 5880 0 clknet_3_0__leaf_clk_i
rlabel metal2 18452 4312 18452 4312 0 clknet_3_1__leaf_clk_i
rlabel metal2 2128 21560 2128 21560 0 clknet_3_2__leaf_clk_i
rlabel metal2 10164 24024 10164 24024 0 clknet_3_3__leaf_clk_i
rlabel metal2 24864 5096 24864 5096 0 clknet_3_4__leaf_clk_i
rlabel metal2 37184 19376 37184 19376 0 clknet_3_5__leaf_clk_i
rlabel metal2 24640 24976 24640 24976 0 clknet_3_6__leaf_clk_i
rlabel metal2 34328 29400 34328 29400 0 clknet_3_7__leaf_clk_i
rlabel metal2 38360 36960 38360 36960 0 custom_setting
rlabel metal3 10472 23128 10472 23128 0 dest\[0\]
rlabel metal2 8008 19712 8008 19712 0 dest\[10\]
rlabel metal2 11872 18424 11872 18424 0 dest\[11\]
rlabel metal2 13048 16912 13048 16912 0 dest\[12\]
rlabel metal2 14336 20440 14336 20440 0 dest\[13\]
rlabel metal2 12768 24052 12768 24052 0 dest\[14\]
rlabel metal2 13664 24220 13664 24220 0 dest\[15\]
rlabel metal2 24808 25424 24808 25424 0 dest\[16\]
rlabel metal3 7532 25480 7532 25480 0 dest\[1\]
rlabel metal2 7112 26376 7112 26376 0 dest\[2\]
rlabel metal2 2016 31052 2016 31052 0 dest\[3\]
rlabel metal2 2520 31416 2520 31416 0 dest\[4\]
rlabel metal2 3136 26348 3136 26348 0 dest\[5\]
rlabel metal2 4760 24920 4760 24920 0 dest\[6\]
rlabel metal2 5544 21280 5544 21280 0 dest\[7\]
rlabel metal2 7336 20888 7336 20888 0 dest\[8\]
rlabel metal3 6720 20776 6720 20776 0 dest\[9\]
rlabel metal3 25144 7448 25144 7448 0 dia\[0\]
rlabel metal2 28392 5544 28392 5544 0 dia\[1\]
rlabel metal3 29288 6664 29288 6664 0 dia\[2\]
rlabel metal2 32648 5320 32648 5320 0 dia\[3\]
rlabel metal2 35672 5936 35672 5936 0 dia\[4\]
rlabel metal2 37688 6608 37688 6608 0 dia\[5\]
rlabel metal3 36736 8232 36736 8232 0 dia\[6\]
rlabel metal2 36512 17752 36512 17752 0 dia\[7\]
rlabel metal3 25648 9800 25648 9800 0 dib\[0\]
rlabel metal2 27832 9828 27832 9828 0 dib\[1\]
rlabel metal2 29288 10136 29288 10136 0 dib\[2\]
rlabel metal2 32760 12488 32760 12488 0 dib\[3\]
rlabel metal3 35784 13888 35784 13888 0 dib\[4\]
rlabel metal2 36568 13216 36568 13216 0 dib\[5\]
rlabel metal3 36288 15288 36288 15288 0 dib\[6\]
rlabel metal2 36344 17416 36344 17416 0 dib\[7\]
rlabel metal2 38360 7896 38360 7896 0 io_in[0]
rlabel metal2 38360 11312 38360 11312 0 io_in[1]
rlabel metal2 38360 14392 38360 14392 0 io_in[2]
rlabel metal2 38360 17360 38360 17360 0 io_in[3]
rlabel metal2 38416 19208 38416 19208 0 io_in[4]
rlabel metal2 38360 23016 38360 23016 0 io_in[5]
rlabel metal3 38794 25816 38794 25816 0 io_in[6]
rlabel metal2 38360 31752 38360 31752 0 io_in[7]
rlabel metal2 15736 34720 15736 34720 0 io_out[10]
rlabel metal2 16184 34832 16184 34832 0 io_out[11]
rlabel metal2 16184 37128 16184 37128 0 io_out[12]
rlabel metal3 18984 33600 18984 33600 0 io_out[13]
rlabel metal2 18872 37842 18872 37842 0 io_out[14]
rlabel metal3 19600 36680 19600 36680 0 io_out[15]
rlabel metal2 22344 35168 22344 35168 0 io_out[16]
rlabel metal2 25928 35616 25928 35616 0 io_out[17]
rlabel metal2 26264 35392 26264 35392 0 io_out[18]
rlabel metal2 24360 36904 24360 36904 0 io_out[19]
rlabel metal2 25592 37170 25592 37170 0 io_out[20]
rlabel metal2 26712 37282 26712 37282 0 io_out[21]
rlabel metal2 27832 37226 27832 37226 0 io_out[22]
rlabel metal2 28952 36834 28952 36834 0 io_out[23]
rlabel metal2 34216 32816 34216 32816 0 io_out[24]
rlabel metal2 31192 37170 31192 37170 0 io_out[25]
rlabel metal3 33152 29960 33152 29960 0 io_out[26]
rlabel metal2 33880 29792 33880 29792 0 io_out[27]
rlabel metal2 34720 28840 34720 28840 0 io_out[28]
rlabel metal2 31528 31808 31528 31808 0 io_out[29]
rlabel metal2 36792 26516 36792 26516 0 io_out[30]
rlabel metal2 12376 37352 12376 37352 0 io_out[8]
rlabel metal3 12824 36456 12824 36456 0 io_out[9]
rlabel metal3 11256 12936 11256 12936 0 mar\[0\]
rlabel metal2 10024 12936 10024 12936 0 mar\[1\]
rlabel metal2 8008 6160 8008 6160 0 mar\[2\]
rlabel metal2 7000 7448 7000 7448 0 mar\[3\]
rlabel metal2 6552 5936 6552 5936 0 mar\[4\]
rlabel metal3 7280 5208 7280 5208 0 mar\[5\]
rlabel metal2 3528 4648 3528 4648 0 mar\[6\]
rlabel metal2 9744 6104 9744 6104 0 mar\[7\]
rlabel metal2 14616 12432 14616 12432 0 mc14500.DATA_OUT
rlabel metal2 31024 35896 31024 35896 0 mc14500.FLAG_O
rlabel metal2 28616 16296 28616 16296 0 mc14500.IEN_l
rlabel metal2 26432 14364 26432 14364 0 mc14500.OEN_l
rlabel metal3 31612 17752 31612 17752 0 mc14500.RR
rlabel via2 20216 12936 20216 12936 0 mc14500.X1
rlabel metal2 22344 12824 22344 12824 0 mc14500.instr_l\[0\]
rlabel metal2 21000 11368 21000 11368 0 mc14500.instr_l\[1\]
rlabel metal2 21504 15932 21504 15932 0 mc14500.instr_l\[2\]
rlabel metal2 20328 14784 20328 14784 0 mc14500.instr_l\[3\]
rlabel metal2 19992 19152 19992 19152 0 mc14500.skip
rlabel metal2 32928 25032 32928 25032 0 net1
rlabel metal3 38668 24584 38668 24584 0 net10
rlabel metal2 19824 8008 19824 8008 0 net11
rlabel metal2 26600 11088 26600 11088 0 net12
rlabel metal2 26796 8680 26796 8680 0 net13
rlabel metal2 30240 6020 30240 6020 0 net14
rlabel metal2 29708 6664 29708 6664 0 net15
rlabel metal2 33936 6188 33936 6188 0 net16
rlabel metal2 35280 4620 35280 4620 0 net17
rlabel metal2 34496 7364 34496 7364 0 net18
rlabel metal2 36064 15176 36064 15176 0 net19
rlabel metal3 25172 25480 25172 25480 0 net2
rlabel via2 7672 30072 7672 30072 0 net20
rlabel metal2 15792 35672 15792 35672 0 net21
rlabel metal2 8904 36008 8904 36008 0 net22
rlabel metal2 17976 33586 17976 33586 0 net23
rlabel metal2 16632 35000 16632 35000 0 net24
rlabel metal3 21280 34888 21280 34888 0 net25
rlabel metal3 19992 31920 19992 31920 0 net26
rlabel metal2 21000 35840 21000 35840 0 net27
rlabel metal2 20888 35840 20888 35840 0 net28
rlabel metal2 23912 24080 23912 24080 0 net29
rlabel metal2 22212 12852 22212 12852 0 net3
rlabel metal3 22708 25256 22708 25256 0 net30
rlabel metal2 26488 30240 26488 30240 0 net31
rlabel metal2 24360 32088 24360 32088 0 net32
rlabel metal2 24136 20888 24136 20888 0 net33
rlabel metal2 28504 28896 28504 28896 0 net34
rlabel metal2 33096 35965 33096 35965 0 net35
rlabel via1 35336 30170 35336 30170 0 net36
rlabel metal2 36120 29581 36120 29581 0 net37
rlabel metal2 36456 30338 36456 30338 0 net38
rlabel metal2 32312 32018 32312 32018 0 net39
rlabel metal2 24528 13552 24528 13552 0 net4
rlabel metal2 35560 30632 35560 30632 0 net40
rlabel metal2 11928 28616 11928 28616 0 net41
rlabel metal2 10360 31136 10360 31136 0 net42
rlabel via2 4200 5082 4200 5082 0 net43
rlabel metal2 2856 3626 2856 3626 0 net44
rlabel metal2 5768 3920 5768 3920 0 net45
rlabel metal2 6552 4605 6552 4605 0 net46
rlabel metal2 6664 4186 6664 4186 0 net47
rlabel metal3 8036 4872 8036 4872 0 net48
rlabel metal2 26320 23688 26320 23688 0 net49
rlabel metal2 18004 13944 18004 13944 0 net5
rlabel metal2 12488 7896 12488 7896 0 net50
rlabel metal3 12096 5992 12096 5992 0 net51
rlabel metal2 13944 3738 13944 3738 0 net52
rlabel metal2 17528 6005 17528 6005 0 net53
rlabel metal2 19040 6748 19040 6748 0 net54
rlabel metal2 21112 5026 21112 5026 0 net55
rlabel metal2 21224 3976 21224 3976 0 net56
rlabel metal2 22120 5936 22120 5936 0 net57
rlabel metal2 20104 27888 20104 27888 0 net58
rlabel metal3 19880 30968 19880 30968 0 net59
rlabel metal2 21784 16990 21784 16990 0 net6
rlabel metal2 17528 32928 17528 32928 0 net60
rlabel via2 16296 35691 16296 35691 0 net61
rlabel metal2 16072 34272 16072 34272 0 net62
rlabel metal2 10920 29960 10920 29960 0 net63
rlabel metal2 12208 28840 12208 28840 0 net64
rlabel metal2 18200 13552 18200 13552 0 net65
rlabel metal2 19432 13832 19432 13832 0 net66
rlabel metal2 23576 13496 23576 13496 0 net67
rlabel metal2 3192 38010 3192 38010 0 net68
rlabel metal2 4592 36596 4592 36596 0 net69
rlabel metal2 37016 20832 37016 20832 0 net7
rlabel metal2 5712 36596 5712 36596 0 net70
rlabel metal2 6832 36596 6832 36596 0 net71
rlabel metal2 7952 36596 7952 36596 0 net72
rlabel metal2 8736 36596 8736 36596 0 net73
rlabel metal2 9744 36372 9744 36372 0 net74
rlabel metal2 11284 35896 11284 35896 0 net75
rlabel metal2 35224 24752 35224 24752 0 net8
rlabel metal2 37912 24752 37912 24752 0 net9
rlabel metal2 33712 34776 33712 34776 0 out_1
rlabel metal2 29848 33544 29848 33544 0 out_2
rlabel metal2 25144 33376 25144 33376 0 rst_latency\[0\]
rlabel metal2 26600 32424 26600 32424 0 rst_latency\[1\]
rlabel metal2 38360 5264 38360 5264 0 rst_n
rlabel metal3 35224 30968 35224 30968 0 scratch\[0\]
rlabel metal2 37464 29624 37464 29624 0 scratch\[1\]
rlabel metal2 35672 20608 35672 20608 0 scratch\[2\]
rlabel metal3 35532 20776 35532 20776 0 scratch\[3\]
rlabel metal2 37688 31416 37688 31416 0 scratch\[4\]
rlabel metal2 32088 29568 32088 29568 0 scratch\[5\]
rlabel metal2 1176 2086 1176 2086 0 sram_addr[0]
rlabel metal2 2968 2086 2968 2086 0 sram_addr[1]
rlabel metal2 4760 2422 4760 2422 0 sram_addr[2]
rlabel metal2 6552 2422 6552 2422 0 sram_addr[3]
rlabel metal2 8344 2142 8344 2142 0 sram_addr[4]
rlabel metal2 10136 798 10136 798 0 sram_addr[5]
rlabel metal3 31472 33320 31472 33320 0 sram_gwe
rlabel metal2 11928 2030 11928 2030 0 sram_in[0]
rlabel metal2 13720 2254 13720 2254 0 sram_in[1]
rlabel metal2 15512 2030 15512 2030 0 sram_in[2]
rlabel metal2 17304 2702 17304 2702 0 sram_in[3]
rlabel metal2 19096 2030 19096 2030 0 sram_in[4]
rlabel metal2 20888 2198 20888 2198 0 sram_in[5]
rlabel metal2 22680 2198 22680 2198 0 sram_in[6]
rlabel metal2 24472 1806 24472 1806 0 sram_in[7]
rlabel metal2 26264 2142 26264 2142 0 sram_out[0]
rlabel metal3 29260 3528 29260 3528 0 sram_out[1]
rlabel metal3 30184 3528 30184 3528 0 sram_out[2]
rlabel metal2 31696 3304 31696 3304 0 sram_out[3]
rlabel metal2 33432 2058 33432 2058 0 sram_out[4]
rlabel metal2 35224 2058 35224 2058 0 sram_out[5]
rlabel metal2 37016 2058 37016 2058 0 sram_out[6]
rlabel metal2 38584 2632 38584 2632 0 sram_out[7]
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
