magic
tech gf180mcuD
magscale 1 5
timestamp 1754054935
<< nwell >>
rect 629 77793 114339 78223
rect 629 77009 114339 77439
rect 629 76225 114339 76655
rect 629 75441 114339 75871
rect 629 74657 114339 75087
rect 629 73873 114339 74303
rect 629 73089 114339 73519
rect 629 72305 114339 72735
rect 629 71521 114339 71951
rect 629 70737 114339 71167
rect 629 69953 114339 70383
rect 629 69169 114339 69599
rect 629 68385 114339 68815
rect 629 67601 114339 68031
rect 629 66817 114339 67247
rect 629 66033 114339 66463
rect 629 65249 114339 65679
rect 629 64465 114339 64895
rect 629 63681 114339 64111
rect 629 62897 114339 63327
rect 629 62113 114339 62543
rect 629 61329 114339 61759
rect 629 60545 114339 60975
rect 629 59761 114339 60191
rect 629 58977 114339 59407
rect 629 58193 114339 58623
rect 629 57409 114339 57839
rect 629 56625 114339 57055
rect 629 55841 114339 56271
rect 629 55057 114339 55487
rect 629 54273 114339 54703
rect 629 53489 114339 53919
rect 629 52705 114339 53135
rect 629 51921 114339 52351
rect 629 51137 114339 51567
rect 629 50353 114339 50783
rect 629 49569 114339 49999
rect 629 48785 114339 49215
rect 629 48001 114339 48431
rect 629 47217 114339 47647
rect 629 46433 114339 46863
rect 629 45649 114339 46079
rect 629 44865 114339 45295
rect 629 44081 114339 44511
rect 629 43297 114339 43727
rect 629 42513 114339 42943
rect 629 41729 114339 42159
rect 629 40945 114339 41375
rect 629 40161 114339 40591
rect 629 39377 114339 39807
rect 629 38593 114339 39023
rect 629 37809 114339 38239
rect 629 37025 114339 37455
rect 629 36241 114339 36671
rect 629 35457 114339 35887
rect 629 34673 114339 35103
rect 629 33889 114339 34319
rect 629 33105 114339 33535
rect 629 32321 114339 32751
rect 629 31537 114339 31967
rect 629 30753 114339 31183
rect 629 29969 114339 30399
rect 629 29185 114339 29615
rect 629 28401 114339 28831
rect 629 27617 114339 28047
rect 629 26833 114339 27263
rect 629 26049 114339 26479
rect 629 25265 114339 25695
rect 629 24481 114339 24911
rect 629 23697 114339 24127
rect 629 22913 114339 23343
rect 629 22129 114339 22559
rect 629 21345 114339 21775
rect 629 20561 114339 20991
rect 629 19777 114339 20207
rect 629 18993 114339 19423
rect 629 18209 114339 18639
rect 629 17425 114339 17855
rect 629 16641 114339 17071
rect 629 15857 114339 16287
rect 629 15073 114339 15503
rect 629 14289 114339 14719
rect 629 13505 114339 13935
rect 629 12721 114339 13151
rect 629 11937 114339 12367
rect 629 11153 114339 11583
rect 629 10369 114339 10799
rect 629 9585 114339 10015
rect 629 8801 114339 9231
rect 629 8017 114339 8447
rect 629 7233 114339 7663
rect 629 6449 114339 6879
rect 629 5665 114339 6095
rect 629 4881 114339 5311
rect 629 4097 114339 4527
rect 629 3313 114339 3743
rect 629 2529 114339 2959
rect 629 1745 114339 2175
<< pwell >>
rect 629 78223 114339 78443
rect 629 77439 114339 77793
rect 629 76655 114339 77009
rect 629 75871 114339 76225
rect 629 75087 114339 75441
rect 629 74303 114339 74657
rect 629 73519 114339 73873
rect 629 72735 114339 73089
rect 629 71951 114339 72305
rect 629 71167 114339 71521
rect 629 70383 114339 70737
rect 629 69599 114339 69953
rect 629 68815 114339 69169
rect 629 68031 114339 68385
rect 629 67247 114339 67601
rect 629 66463 114339 66817
rect 629 65679 114339 66033
rect 629 64895 114339 65249
rect 629 64111 114339 64465
rect 629 63327 114339 63681
rect 629 62543 114339 62897
rect 629 61759 114339 62113
rect 629 60975 114339 61329
rect 629 60191 114339 60545
rect 629 59407 114339 59761
rect 629 58623 114339 58977
rect 629 57839 114339 58193
rect 629 57055 114339 57409
rect 629 56271 114339 56625
rect 629 55487 114339 55841
rect 629 54703 114339 55057
rect 629 53919 114339 54273
rect 629 53135 114339 53489
rect 629 52351 114339 52705
rect 629 51567 114339 51921
rect 629 50783 114339 51137
rect 629 49999 114339 50353
rect 629 49215 114339 49569
rect 629 48431 114339 48785
rect 629 47647 114339 48001
rect 629 46863 114339 47217
rect 629 46079 114339 46433
rect 629 45295 114339 45649
rect 629 44511 114339 44865
rect 629 43727 114339 44081
rect 629 42943 114339 43297
rect 629 42159 114339 42513
rect 629 41375 114339 41729
rect 629 40591 114339 40945
rect 629 39807 114339 40161
rect 629 39023 114339 39377
rect 629 38239 114339 38593
rect 629 37455 114339 37809
rect 629 36671 114339 37025
rect 629 35887 114339 36241
rect 629 35103 114339 35457
rect 629 34319 114339 34673
rect 629 33535 114339 33889
rect 629 32751 114339 33105
rect 629 31967 114339 32321
rect 629 31183 114339 31537
rect 629 30399 114339 30753
rect 629 29615 114339 29969
rect 629 28831 114339 29185
rect 629 28047 114339 28401
rect 629 27263 114339 27617
rect 629 26479 114339 26833
rect 629 25695 114339 26049
rect 629 24911 114339 25265
rect 629 24127 114339 24481
rect 629 23343 114339 23697
rect 629 22559 114339 22913
rect 629 21775 114339 22129
rect 629 20991 114339 21345
rect 629 20207 114339 20561
rect 629 19423 114339 19777
rect 629 18639 114339 18993
rect 629 17855 114339 18209
rect 629 17071 114339 17425
rect 629 16287 114339 16641
rect 629 15503 114339 15857
rect 629 14719 114339 15073
rect 629 13935 114339 14289
rect 629 13151 114339 13505
rect 629 12367 114339 12721
rect 629 11583 114339 11937
rect 629 10799 114339 11153
rect 629 10015 114339 10369
rect 629 9231 114339 9585
rect 629 8447 114339 8801
rect 629 7663 114339 8017
rect 629 6879 114339 7233
rect 629 6095 114339 6449
rect 629 5311 114339 5665
rect 629 4527 114339 4881
rect 629 3743 114339 4097
rect 629 2959 114339 3313
rect 629 2175 114339 2529
rect 629 1525 114339 1745
<< obsm1 >>
rect 672 1538 114296 78497
<< metal2 >>
rect 57456 79600 57512 80000
rect 28672 0 28728 400
rect 86128 0 86184 400
<< obsm2 >>
rect 798 79570 57426 79600
rect 57542 79570 114226 79600
rect 798 430 114226 79570
rect 798 400 28642 430
rect 28758 400 86098 430
rect 86214 400 114226 430
<< metal3 >>
rect 114600 78512 115000 78568
rect 114600 77056 115000 77112
rect 114600 75600 115000 75656
rect 114600 74144 115000 74200
rect 114600 72688 115000 72744
rect 114600 71232 115000 71288
rect 114600 69776 115000 69832
rect 114600 68320 115000 68376
rect 114600 66864 115000 66920
rect 114600 65408 115000 65464
rect 114600 63952 115000 64008
rect 114600 62496 115000 62552
rect 114600 61040 115000 61096
rect 114600 59584 115000 59640
rect 114600 58128 115000 58184
rect 114600 56672 115000 56728
rect 114600 55216 115000 55272
rect 114600 53760 115000 53816
rect 114600 52304 115000 52360
rect 114600 50848 115000 50904
rect 114600 49392 115000 49448
rect 114600 47936 115000 47992
rect 114600 46480 115000 46536
rect 114600 45024 115000 45080
rect 114600 43568 115000 43624
rect 114600 42112 115000 42168
rect 114600 40656 115000 40712
rect 114600 39200 115000 39256
rect 114600 37744 115000 37800
rect 114600 36288 115000 36344
rect 114600 34832 115000 34888
rect 114600 33376 115000 33432
rect 114600 31920 115000 31976
rect 114600 30464 115000 30520
rect 114600 29008 115000 29064
rect 114600 27552 115000 27608
rect 114600 26096 115000 26152
rect 114600 24640 115000 24696
rect 114600 23184 115000 23240
rect 114600 21728 115000 21784
rect 114600 20272 115000 20328
rect 114600 18816 115000 18872
rect 114600 17360 115000 17416
rect 114600 15904 115000 15960
rect 114600 14448 115000 14504
rect 114600 12992 115000 13048
rect 114600 11536 115000 11592
rect 114600 10080 115000 10136
rect 114600 8624 115000 8680
rect 114600 7168 115000 7224
rect 114600 5712 115000 5768
rect 114600 4256 115000 4312
rect 114600 2800 115000 2856
rect 114600 1344 115000 1400
<< obsm3 >>
rect 793 78598 114674 79226
rect 793 78482 114570 78598
rect 793 77142 114674 78482
rect 793 77026 114570 77142
rect 793 75686 114674 77026
rect 793 75570 114570 75686
rect 793 74230 114674 75570
rect 793 74114 114570 74230
rect 793 72774 114674 74114
rect 793 72658 114570 72774
rect 793 71318 114674 72658
rect 793 71202 114570 71318
rect 793 69862 114674 71202
rect 793 69746 114570 69862
rect 793 68406 114674 69746
rect 793 68290 114570 68406
rect 793 66950 114674 68290
rect 793 66834 114570 66950
rect 793 65494 114674 66834
rect 793 65378 114570 65494
rect 793 64038 114674 65378
rect 793 63922 114570 64038
rect 793 62582 114674 63922
rect 793 62466 114570 62582
rect 793 61126 114674 62466
rect 793 61010 114570 61126
rect 793 59670 114674 61010
rect 793 59554 114570 59670
rect 793 58214 114674 59554
rect 793 58098 114570 58214
rect 793 56758 114674 58098
rect 793 56642 114570 56758
rect 793 55302 114674 56642
rect 793 55186 114570 55302
rect 793 53846 114674 55186
rect 793 53730 114570 53846
rect 793 52390 114674 53730
rect 793 52274 114570 52390
rect 793 50934 114674 52274
rect 793 50818 114570 50934
rect 793 49478 114674 50818
rect 793 49362 114570 49478
rect 793 48022 114674 49362
rect 793 47906 114570 48022
rect 793 46566 114674 47906
rect 793 46450 114570 46566
rect 793 45110 114674 46450
rect 793 44994 114570 45110
rect 793 43654 114674 44994
rect 793 43538 114570 43654
rect 793 42198 114674 43538
rect 793 42082 114570 42198
rect 793 40742 114674 42082
rect 793 40626 114570 40742
rect 793 39286 114674 40626
rect 793 39170 114570 39286
rect 793 37830 114674 39170
rect 793 37714 114570 37830
rect 793 36374 114674 37714
rect 793 36258 114570 36374
rect 793 34918 114674 36258
rect 793 34802 114570 34918
rect 793 33462 114674 34802
rect 793 33346 114570 33462
rect 793 32006 114674 33346
rect 793 31890 114570 32006
rect 793 30550 114674 31890
rect 793 30434 114570 30550
rect 793 29094 114674 30434
rect 793 28978 114570 29094
rect 793 27638 114674 28978
rect 793 27522 114570 27638
rect 793 26182 114674 27522
rect 793 26066 114570 26182
rect 793 24726 114674 26066
rect 793 24610 114570 24726
rect 793 23270 114674 24610
rect 793 23154 114570 23270
rect 793 21814 114674 23154
rect 793 21698 114570 21814
rect 793 20358 114674 21698
rect 793 20242 114570 20358
rect 793 18902 114674 20242
rect 793 18786 114570 18902
rect 793 17446 114674 18786
rect 793 17330 114570 17446
rect 793 15990 114674 17330
rect 793 15874 114570 15990
rect 793 14534 114674 15874
rect 793 14418 114570 14534
rect 793 13078 114674 14418
rect 793 12962 114570 13078
rect 793 11622 114674 12962
rect 793 11506 114570 11622
rect 793 10166 114674 11506
rect 793 10050 114570 10166
rect 793 8710 114674 10050
rect 793 8594 114570 8710
rect 793 7254 114674 8594
rect 793 7138 114570 7254
rect 793 5798 114674 7138
rect 793 5682 114570 5798
rect 793 4342 114674 5682
rect 793 4226 114570 4342
rect 793 2886 114674 4226
rect 793 2770 114570 2886
rect 793 1430 114674 2770
rect 793 1358 114570 1430
<< metal4 >>
rect 2224 1538 2384 78430
rect 9904 1538 10064 78430
rect 17584 1538 17744 78430
rect 25264 1538 25424 78430
rect 32944 1538 33104 78430
rect 40624 1538 40784 78430
rect 48304 1538 48464 78430
rect 55984 1538 56144 78430
rect 63664 1538 63824 78430
rect 71344 1538 71504 78430
rect 79024 1538 79184 78430
rect 86704 1538 86864 78430
rect 94384 1538 94544 78430
rect 102064 1538 102224 78430
rect 109744 1538 109904 78430
<< obsm4 >>
rect 1358 2529 2194 76767
rect 2414 2529 9874 76767
rect 10094 2529 17554 76767
rect 17774 2529 25234 76767
rect 25454 2529 32914 76767
rect 33134 2529 40594 76767
rect 40814 2529 48274 76767
rect 48494 2529 55954 76767
rect 56174 2529 63634 76767
rect 63854 2529 71314 76767
rect 71534 2529 78994 76767
rect 79214 2529 86674 76767
rect 86894 2529 94354 76767
rect 94574 2529 102034 76767
rect 102254 2529 109714 76767
rect 109934 2529 113386 76767
<< labels >>
rlabel metal3 s 114600 1344 115000 1400 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 114600 15904 115000 15960 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 114600 17360 115000 17416 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 114600 18816 115000 18872 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 114600 20272 115000 20328 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 114600 21728 115000 21784 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 114600 23184 115000 23240 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 114600 24640 115000 24696 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 114600 26096 115000 26152 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 114600 27552 115000 27608 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 114600 29008 115000 29064 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 114600 2800 115000 2856 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 114600 30464 115000 30520 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 114600 31920 115000 31976 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 114600 33376 115000 33432 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 114600 34832 115000 34888 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 114600 36288 115000 36344 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 114600 37744 115000 37800 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 114600 39200 115000 39256 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 114600 40656 115000 40712 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 114600 42112 115000 42168 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 114600 43568 115000 43624 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 114600 4256 115000 4312 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 114600 45024 115000 45080 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 114600 46480 115000 46536 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 114600 47936 115000 47992 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 114600 5712 115000 5768 6 io_in[3]
port 27 nsew signal input
rlabel metal3 s 114600 7168 115000 7224 6 io_in[4]
port 28 nsew signal input
rlabel metal3 s 114600 8624 115000 8680 6 io_in[5]
port 29 nsew signal input
rlabel metal3 s 114600 10080 115000 10136 6 io_in[6]
port 30 nsew signal input
rlabel metal3 s 114600 11536 115000 11592 6 io_in[7]
port 31 nsew signal input
rlabel metal3 s 114600 12992 115000 13048 6 io_in[8]
port 32 nsew signal input
rlabel metal3 s 114600 14448 115000 14504 6 io_in[9]
port 33 nsew signal input
rlabel metal2 s 57456 79600 57512 80000 6 io_oeb
port 34 nsew signal output
rlabel metal3 s 114600 49392 115000 49448 6 io_out[0]
port 35 nsew signal output
rlabel metal3 s 114600 63952 115000 64008 6 io_out[10]
port 36 nsew signal output
rlabel metal3 s 114600 65408 115000 65464 6 io_out[11]
port 37 nsew signal output
rlabel metal3 s 114600 66864 115000 66920 6 io_out[12]
port 38 nsew signal output
rlabel metal3 s 114600 68320 115000 68376 6 io_out[13]
port 39 nsew signal output
rlabel metal3 s 114600 69776 115000 69832 6 io_out[14]
port 40 nsew signal output
rlabel metal3 s 114600 71232 115000 71288 6 io_out[15]
port 41 nsew signal output
rlabel metal3 s 114600 72688 115000 72744 6 io_out[16]
port 42 nsew signal output
rlabel metal3 s 114600 74144 115000 74200 6 io_out[17]
port 43 nsew signal output
rlabel metal3 s 114600 75600 115000 75656 6 io_out[18]
port 44 nsew signal output
rlabel metal3 s 114600 77056 115000 77112 6 io_out[19]
port 45 nsew signal output
rlabel metal3 s 114600 50848 115000 50904 6 io_out[1]
port 46 nsew signal output
rlabel metal3 s 114600 78512 115000 78568 6 io_out[20]
port 47 nsew signal output
rlabel metal3 s 114600 52304 115000 52360 6 io_out[2]
port 48 nsew signal output
rlabel metal3 s 114600 53760 115000 53816 6 io_out[3]
port 49 nsew signal output
rlabel metal3 s 114600 55216 115000 55272 6 io_out[4]
port 50 nsew signal output
rlabel metal3 s 114600 56672 115000 56728 6 io_out[5]
port 51 nsew signal output
rlabel metal3 s 114600 58128 115000 58184 6 io_out[6]
port 52 nsew signal output
rlabel metal3 s 114600 59584 115000 59640 6 io_out[7]
port 53 nsew signal output
rlabel metal3 s 114600 61040 115000 61096 6 io_out[8]
port 54 nsew signal output
rlabel metal3 s 114600 62496 115000 62552 6 io_out[9]
port 55 nsew signal output
rlabel metal2 s 86128 0 86184 400 6 rst_n
port 56 nsew signal input
rlabel metal4 s 2224 1538 2384 78430 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 78430 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 78430 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 78430 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 78430 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 78430 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 78430 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 78430 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 78430 6 vss
port 58 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 78430 6 vss
port 58 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 78430 6 vss
port 58 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 78430 6 vss
port 58 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 78430 6 vss
port 58 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 78430 6 vss
port 58 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 78430 6 vss
port 58 nsew ground bidirectional
rlabel metal2 s 28672 0 28728 400 6 wb_clk_i
port 59 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 115000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 30428416
string GDS_FILE /home/lucah/gfmpw1-multi/openlane/wrapped_sid/runs/25_08_01_15_03/results/signoff/wrapped_sid.magic.gds
string GDS_START 297614
<< end >>

