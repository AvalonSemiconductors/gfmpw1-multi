magic
tech gf180mcuD
magscale 1 10
timestamp 1712524553
<< metal1 >>
rect 1344 42362 44576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 44576 42362
rect 1344 42276 44576 42310
rect 18286 42194 18338 42206
rect 18286 42130 18338 42142
rect 33518 42194 33570 42206
rect 33518 42130 33570 42142
rect 6178 42030 6190 42082
rect 6242 42030 6254 42082
rect 9986 42030 9998 42082
rect 10050 42030 10062 42082
rect 5070 41970 5122 41982
rect 5070 41906 5122 41918
rect 5854 41970 5906 41982
rect 5854 41906 5906 41918
rect 8878 41970 8930 41982
rect 8878 41906 8930 41918
rect 9662 41970 9714 41982
rect 13458 41918 13470 41970
rect 13522 41918 13534 41970
rect 17266 41918 17278 41970
rect 17330 41918 17342 41970
rect 21074 41918 21086 41970
rect 21138 41918 21150 41970
rect 24882 41918 24894 41970
rect 24946 41918 24958 41970
rect 28690 41918 28702 41970
rect 28754 41918 28766 41970
rect 30370 41918 30382 41970
rect 30434 41918 30446 41970
rect 32498 41918 32510 41970
rect 32562 41918 32574 41970
rect 36306 41918 36318 41970
rect 36370 41918 36382 41970
rect 40114 41918 40126 41970
rect 40178 41918 40190 41970
rect 9662 41906 9714 41918
rect 14478 41858 14530 41870
rect 14478 41794 14530 41806
rect 22094 41858 22146 41870
rect 22094 41794 22146 41806
rect 25902 41858 25954 41870
rect 25902 41794 25954 41806
rect 37326 41858 37378 41870
rect 37326 41794 37378 41806
rect 41134 41858 41186 41870
rect 41134 41794 41186 41806
rect 1344 41578 44576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 44576 41578
rect 1344 41492 44576 41526
rect 43150 41410 43202 41422
rect 43150 41346 43202 41358
rect 43922 41134 43934 41186
rect 43986 41134 43998 41186
rect 39790 40962 39842 40974
rect 39790 40898 39842 40910
rect 1344 40794 44576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 44576 40794
rect 1344 40708 44576 40742
rect 15710 40626 15762 40638
rect 15710 40562 15762 40574
rect 16718 40626 16770 40638
rect 16718 40562 16770 40574
rect 11566 40514 11618 40526
rect 11566 40450 11618 40462
rect 12126 40514 12178 40526
rect 12126 40450 12178 40462
rect 12350 40514 12402 40526
rect 15486 40514 15538 40526
rect 14690 40462 14702 40514
rect 14754 40462 14766 40514
rect 12350 40450 12402 40462
rect 15486 40450 15538 40462
rect 16942 40514 16994 40526
rect 16942 40450 16994 40462
rect 5630 40402 5682 40414
rect 9774 40402 9826 40414
rect 2258 40350 2270 40402
rect 2322 40350 2334 40402
rect 2930 40350 2942 40402
rect 2994 40350 3006 40402
rect 6178 40350 6190 40402
rect 6242 40350 6254 40402
rect 5630 40338 5682 40350
rect 9774 40338 9826 40350
rect 11342 40402 11394 40414
rect 11342 40338 11394 40350
rect 11678 40402 11730 40414
rect 11678 40338 11730 40350
rect 12574 40402 12626 40414
rect 12574 40338 12626 40350
rect 14366 40402 14418 40414
rect 14366 40338 14418 40350
rect 15374 40402 15426 40414
rect 15374 40338 15426 40350
rect 16606 40402 16658 40414
rect 16606 40338 16658 40350
rect 20078 40402 20130 40414
rect 31950 40402 32002 40414
rect 40462 40402 40514 40414
rect 20290 40350 20302 40402
rect 20354 40350 20366 40402
rect 25330 40350 25342 40402
rect 25394 40350 25406 40402
rect 28578 40350 28590 40402
rect 28642 40350 28654 40402
rect 37426 40350 37438 40402
rect 37490 40350 37502 40402
rect 41010 40350 41022 40402
rect 41074 40350 41086 40402
rect 20078 40338 20130 40350
rect 31950 40338 32002 40350
rect 40462 40338 40514 40350
rect 12462 40290 12514 40302
rect 38110 40290 38162 40302
rect 5058 40238 5070 40290
rect 5122 40238 5134 40290
rect 6850 40238 6862 40290
rect 6914 40238 6926 40290
rect 8978 40238 8990 40290
rect 9042 40238 9054 40290
rect 21074 40238 21086 40290
rect 21138 40238 21150 40290
rect 23202 40238 23214 40290
rect 23266 40238 23278 40290
rect 26002 40238 26014 40290
rect 26066 40238 26078 40290
rect 28130 40238 28142 40290
rect 28194 40238 28206 40290
rect 29250 40238 29262 40290
rect 29314 40238 29326 40290
rect 31378 40238 31390 40290
rect 31442 40238 31454 40290
rect 34626 40238 34638 40290
rect 34690 40238 34702 40290
rect 36754 40238 36766 40290
rect 36818 40238 36830 40290
rect 41794 40238 41806 40290
rect 41858 40238 41870 40290
rect 43922 40238 43934 40290
rect 43986 40238 43998 40290
rect 12462 40226 12514 40238
rect 38110 40226 38162 40238
rect 1344 40010 44576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 44576 40010
rect 1344 39924 44576 39958
rect 11230 39730 11282 39742
rect 11230 39666 11282 39678
rect 12014 39730 12066 39742
rect 12014 39666 12066 39678
rect 16046 39730 16098 39742
rect 21422 39730 21474 39742
rect 41246 39730 41298 39742
rect 20738 39678 20750 39730
rect 20802 39678 20814 39730
rect 31602 39678 31614 39730
rect 31666 39678 31678 39730
rect 33730 39678 33742 39730
rect 33794 39678 33806 39730
rect 40786 39678 40798 39730
rect 40850 39678 40862 39730
rect 16046 39666 16098 39678
rect 21422 39666 21474 39678
rect 41246 39666 41298 39678
rect 42702 39730 42754 39742
rect 42702 39666 42754 39678
rect 11006 39618 11058 39630
rect 11006 39554 11058 39566
rect 14254 39618 14306 39630
rect 14254 39554 14306 39566
rect 14926 39618 14978 39630
rect 15598 39618 15650 39630
rect 28366 39618 28418 39630
rect 34190 39618 34242 39630
rect 15250 39566 15262 39618
rect 15314 39566 15326 39618
rect 17826 39566 17838 39618
rect 17890 39566 17902 39618
rect 18610 39566 18622 39618
rect 18674 39566 18686 39618
rect 30930 39566 30942 39618
rect 30994 39566 31006 39618
rect 37874 39566 37886 39618
rect 37938 39566 37950 39618
rect 14926 39554 14978 39566
rect 15598 39554 15650 39566
rect 28366 39554 28418 39566
rect 34190 39554 34242 39566
rect 7982 39506 8034 39518
rect 7982 39442 8034 39454
rect 8318 39506 8370 39518
rect 8318 39442 8370 39454
rect 14030 39506 14082 39518
rect 14030 39442 14082 39454
rect 16830 39506 16882 39518
rect 38658 39454 38670 39506
rect 38722 39454 38734 39506
rect 16830 39442 16882 39454
rect 11678 39394 11730 39406
rect 10658 39342 10670 39394
rect 10722 39342 10734 39394
rect 11678 39330 11730 39342
rect 11902 39394 11954 39406
rect 11902 39330 11954 39342
rect 12126 39394 12178 39406
rect 15486 39394 15538 39406
rect 14578 39342 14590 39394
rect 14642 39342 14654 39394
rect 12126 39330 12178 39342
rect 15486 39330 15538 39342
rect 15934 39394 15986 39406
rect 15934 39330 15986 39342
rect 16158 39394 16210 39406
rect 16158 39330 16210 39342
rect 16382 39394 16434 39406
rect 16382 39330 16434 39342
rect 16942 39394 16994 39406
rect 16942 39330 16994 39342
rect 17054 39394 17106 39406
rect 17054 39330 17106 39342
rect 37550 39394 37602 39406
rect 37550 39330 37602 39342
rect 41134 39394 41186 39406
rect 41134 39330 41186 39342
rect 42590 39394 42642 39406
rect 42590 39330 42642 39342
rect 1344 39226 44576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 44576 39226
rect 1344 39140 44576 39174
rect 13918 39058 13970 39070
rect 13918 38994 13970 39006
rect 15150 39058 15202 39070
rect 15150 38994 15202 39006
rect 15710 39058 15762 39070
rect 15710 38994 15762 39006
rect 12574 38946 12626 38958
rect 12574 38882 12626 38894
rect 12686 38946 12738 38958
rect 12686 38882 12738 38894
rect 15486 38946 15538 38958
rect 15486 38882 15538 38894
rect 13806 38834 13858 38846
rect 13806 38770 13858 38782
rect 14030 38834 14082 38846
rect 14030 38770 14082 38782
rect 14478 38834 14530 38846
rect 14478 38770 14530 38782
rect 15038 38834 15090 38846
rect 15038 38770 15090 38782
rect 15810 38670 15822 38722
rect 15874 38670 15886 38722
rect 1344 38442 44576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 44576 38442
rect 1344 38356 44576 38390
rect 26014 38162 26066 38174
rect 37102 38162 37154 38174
rect 2706 38110 2718 38162
rect 2770 38110 2782 38162
rect 4834 38110 4846 38162
rect 4898 38110 4910 38162
rect 7186 38110 7198 38162
rect 7250 38110 7262 38162
rect 9314 38110 9326 38162
rect 9378 38110 9390 38162
rect 25554 38110 25566 38162
rect 25618 38110 25630 38162
rect 31938 38110 31950 38162
rect 32002 38110 32014 38162
rect 26014 38098 26066 38110
rect 37102 38098 37154 38110
rect 12014 38050 12066 38062
rect 39454 38050 39506 38062
rect 2034 37998 2046 38050
rect 2098 37998 2110 38050
rect 6402 37998 6414 38050
rect 6466 37998 6478 38050
rect 22754 37998 22766 38050
rect 22818 37998 22830 38050
rect 34850 37998 34862 38050
rect 34914 37998 34926 38050
rect 12014 37986 12066 37998
rect 39454 37986 39506 37998
rect 39566 38050 39618 38062
rect 39566 37986 39618 37998
rect 11678 37938 11730 37950
rect 36990 37938 37042 37950
rect 23426 37886 23438 37938
rect 23490 37886 23502 37938
rect 34066 37886 34078 37938
rect 34130 37886 34142 37938
rect 11678 37874 11730 37886
rect 36990 37874 37042 37886
rect 37326 37938 37378 37950
rect 37326 37874 37378 37886
rect 37550 37938 37602 37950
rect 37550 37874 37602 37886
rect 39902 37938 39954 37950
rect 39902 37874 39954 37886
rect 5742 37826 5794 37838
rect 5742 37762 5794 37774
rect 9774 37826 9826 37838
rect 9774 37762 9826 37774
rect 11790 37826 11842 37838
rect 11790 37762 11842 37774
rect 12462 37826 12514 37838
rect 12462 37762 12514 37774
rect 35310 37826 35362 37838
rect 35310 37762 35362 37774
rect 39790 37826 39842 37838
rect 39790 37762 39842 37774
rect 40798 37826 40850 37838
rect 40798 37762 40850 37774
rect 1344 37658 44576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 44576 37658
rect 1344 37572 44576 37606
rect 10670 37490 10722 37502
rect 10670 37426 10722 37438
rect 11118 37490 11170 37502
rect 11118 37426 11170 37438
rect 39006 37490 39058 37502
rect 39006 37426 39058 37438
rect 39790 37490 39842 37502
rect 39790 37426 39842 37438
rect 9886 37378 9938 37390
rect 39902 37378 39954 37390
rect 3714 37326 3726 37378
rect 3778 37326 3790 37378
rect 10322 37326 10334 37378
rect 10386 37326 10398 37378
rect 12226 37326 12238 37378
rect 12290 37326 12302 37378
rect 14242 37326 14254 37378
rect 14306 37326 14318 37378
rect 16258 37326 16270 37378
rect 16322 37326 16334 37378
rect 25554 37326 25566 37378
rect 25618 37326 25630 37378
rect 41906 37326 41918 37378
rect 41970 37326 41982 37378
rect 9886 37314 9938 37326
rect 39902 37314 39954 37326
rect 11006 37266 11058 37278
rect 3042 37214 3054 37266
rect 3106 37214 3118 37266
rect 11006 37202 11058 37214
rect 11230 37266 11282 37278
rect 11230 37202 11282 37214
rect 11566 37266 11618 37278
rect 25230 37266 25282 37278
rect 32062 37266 32114 37278
rect 39230 37266 39282 37278
rect 12338 37214 12350 37266
rect 12402 37214 12414 37266
rect 14466 37214 14478 37266
rect 14530 37214 14542 37266
rect 15586 37214 15598 37266
rect 15650 37214 15662 37266
rect 31602 37214 31614 37266
rect 31666 37214 31678 37266
rect 38546 37214 38558 37266
rect 38610 37214 38622 37266
rect 38770 37214 38782 37266
rect 38834 37214 38846 37266
rect 11566 37202 11618 37214
rect 25230 37202 25282 37214
rect 32062 37202 32114 37214
rect 39230 37202 39282 37214
rect 39566 37266 39618 37278
rect 40226 37214 40238 37266
rect 40290 37214 40302 37266
rect 41234 37214 41246 37266
rect 41298 37214 41310 37266
rect 39566 37202 39618 37214
rect 6302 37154 6354 37166
rect 5842 37102 5854 37154
rect 5906 37102 5918 37154
rect 6302 37090 6354 37102
rect 16718 37154 16770 37166
rect 16718 37090 16770 37102
rect 19630 37154 19682 37166
rect 34414 37154 34466 37166
rect 28690 37102 28702 37154
rect 28754 37102 28766 37154
rect 30818 37102 30830 37154
rect 30882 37102 30894 37154
rect 38434 37102 38446 37154
rect 38498 37102 38510 37154
rect 40338 37102 40350 37154
rect 40402 37102 40414 37154
rect 44034 37102 44046 37154
rect 44098 37102 44110 37154
rect 19630 37090 19682 37102
rect 34414 37090 34466 37102
rect 9998 37042 10050 37054
rect 9998 36978 10050 36990
rect 1344 36874 44576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 44576 36874
rect 1344 36788 44576 36822
rect 25566 36706 25618 36718
rect 14242 36654 14254 36706
rect 14306 36654 14318 36706
rect 25566 36642 25618 36654
rect 6974 36594 7026 36606
rect 6974 36530 7026 36542
rect 12014 36594 12066 36606
rect 12014 36530 12066 36542
rect 12350 36594 12402 36606
rect 12350 36530 12402 36542
rect 12910 36594 12962 36606
rect 32286 36594 32338 36606
rect 34526 36594 34578 36606
rect 14802 36542 14814 36594
rect 14866 36542 14878 36594
rect 24546 36542 24558 36594
rect 24610 36542 24622 36594
rect 33842 36542 33854 36594
rect 33906 36542 33918 36594
rect 12910 36530 12962 36542
rect 32286 36530 32338 36542
rect 34526 36530 34578 36542
rect 35422 36594 35474 36606
rect 35422 36530 35474 36542
rect 37438 36594 37490 36606
rect 37438 36530 37490 36542
rect 39454 36594 39506 36606
rect 39454 36530 39506 36542
rect 12574 36482 12626 36494
rect 13806 36482 13858 36494
rect 13458 36430 13470 36482
rect 13522 36430 13534 36482
rect 12574 36418 12626 36430
rect 13806 36418 13858 36430
rect 14478 36482 14530 36494
rect 14478 36418 14530 36430
rect 15486 36482 15538 36494
rect 15486 36418 15538 36430
rect 18398 36482 18450 36494
rect 18398 36418 18450 36430
rect 19070 36482 19122 36494
rect 19070 36418 19122 36430
rect 19294 36482 19346 36494
rect 26462 36482 26514 36494
rect 24770 36430 24782 36482
rect 24834 36430 24846 36482
rect 19294 36418 19346 36430
rect 26462 36418 26514 36430
rect 34078 36482 34130 36494
rect 34078 36418 34130 36430
rect 34414 36482 34466 36494
rect 34414 36418 34466 36430
rect 34638 36482 34690 36494
rect 34638 36418 34690 36430
rect 39342 36482 39394 36494
rect 39342 36418 39394 36430
rect 13694 36370 13746 36382
rect 13694 36306 13746 36318
rect 15038 36370 15090 36382
rect 15038 36306 15090 36318
rect 19966 36370 20018 36382
rect 24110 36370 24162 36382
rect 20290 36318 20302 36370
rect 20354 36318 20366 36370
rect 19966 36306 20018 36318
rect 24110 36306 24162 36318
rect 25790 36370 25842 36382
rect 25790 36306 25842 36318
rect 26350 36370 26402 36382
rect 33742 36370 33794 36382
rect 33506 36318 33518 36370
rect 33570 36318 33582 36370
rect 26350 36306 26402 36318
rect 33742 36306 33794 36318
rect 34974 36370 35026 36382
rect 34974 36306 35026 36318
rect 7086 36258 7138 36270
rect 7086 36194 7138 36206
rect 14814 36258 14866 36270
rect 14814 36194 14866 36206
rect 18062 36258 18114 36270
rect 18062 36194 18114 36206
rect 18286 36258 18338 36270
rect 25678 36258 25730 36270
rect 18722 36206 18734 36258
rect 18786 36206 18798 36258
rect 18286 36194 18338 36206
rect 25678 36194 25730 36206
rect 26126 36258 26178 36270
rect 26126 36194 26178 36206
rect 32398 36258 32450 36270
rect 32398 36194 32450 36206
rect 33854 36258 33906 36270
rect 33854 36194 33906 36206
rect 37102 36258 37154 36270
rect 37102 36194 37154 36206
rect 37326 36258 37378 36270
rect 37326 36194 37378 36206
rect 37550 36258 37602 36270
rect 37550 36194 37602 36206
rect 39118 36258 39170 36270
rect 39118 36194 39170 36206
rect 39566 36258 39618 36270
rect 39566 36194 39618 36206
rect 40014 36258 40066 36270
rect 40014 36194 40066 36206
rect 40574 36258 40626 36270
rect 40574 36194 40626 36206
rect 1344 36090 44576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 44576 36090
rect 1344 36004 44576 36038
rect 34414 35922 34466 35934
rect 10770 35870 10782 35922
rect 10834 35870 10846 35922
rect 13570 35870 13582 35922
rect 13634 35870 13646 35922
rect 14578 35870 14590 35922
rect 14642 35870 14654 35922
rect 34414 35858 34466 35870
rect 36654 35922 36706 35934
rect 36654 35858 36706 35870
rect 10222 35810 10274 35822
rect 10222 35746 10274 35758
rect 13022 35810 13074 35822
rect 17726 35810 17778 35822
rect 14690 35758 14702 35810
rect 14754 35758 14766 35810
rect 15474 35758 15486 35810
rect 15538 35758 15550 35810
rect 13022 35746 13074 35758
rect 17726 35746 17778 35758
rect 20974 35810 21026 35822
rect 34638 35810 34690 35822
rect 26898 35758 26910 35810
rect 26962 35758 26974 35810
rect 20974 35746 21026 35758
rect 34638 35746 34690 35758
rect 13246 35698 13298 35710
rect 13246 35634 13298 35646
rect 14590 35698 14642 35710
rect 14590 35634 14642 35646
rect 17278 35698 17330 35710
rect 19182 35698 19234 35710
rect 19966 35698 20018 35710
rect 18162 35646 18174 35698
rect 18226 35646 18238 35698
rect 19506 35646 19518 35698
rect 19570 35646 19582 35698
rect 17278 35634 17330 35646
rect 19182 35634 19234 35646
rect 19966 35634 20018 35646
rect 20078 35698 20130 35710
rect 25230 35698 25282 35710
rect 34750 35698 34802 35710
rect 20290 35646 20302 35698
rect 20354 35646 20366 35698
rect 21634 35646 21646 35698
rect 21698 35646 21710 35698
rect 25890 35646 25902 35698
rect 25954 35646 25966 35698
rect 20078 35634 20130 35646
rect 25230 35634 25282 35646
rect 34750 35634 34802 35646
rect 36542 35698 36594 35710
rect 36542 35634 36594 35646
rect 36766 35698 36818 35710
rect 36766 35634 36818 35646
rect 37214 35698 37266 35710
rect 37214 35634 37266 35646
rect 36206 35586 36258 35598
rect 21746 35534 21758 35586
rect 21810 35534 21822 35586
rect 27346 35534 27358 35586
rect 27410 35534 27422 35586
rect 36206 35522 36258 35534
rect 10446 35474 10498 35486
rect 18834 35422 18846 35474
rect 18898 35422 18910 35474
rect 10446 35410 10498 35422
rect 1344 35306 44576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 44576 35306
rect 1344 35220 44576 35254
rect 16606 35138 16658 35150
rect 16606 35074 16658 35086
rect 18286 35138 18338 35150
rect 18286 35074 18338 35086
rect 18622 35138 18674 35150
rect 18622 35074 18674 35086
rect 37438 35138 37490 35150
rect 37438 35074 37490 35086
rect 40910 35138 40962 35150
rect 40910 35074 40962 35086
rect 16718 35026 16770 35038
rect 14802 34974 14814 35026
rect 14866 34974 14878 35026
rect 16718 34962 16770 34974
rect 19294 35026 19346 35038
rect 19294 34962 19346 34974
rect 20750 35026 20802 35038
rect 20750 34962 20802 34974
rect 25902 35026 25954 35038
rect 25902 34962 25954 34974
rect 19742 34914 19794 34926
rect 15026 34862 15038 34914
rect 15090 34862 15102 34914
rect 19742 34850 19794 34862
rect 21310 34914 21362 34926
rect 21310 34850 21362 34862
rect 25790 34914 25842 34926
rect 25790 34850 25842 34862
rect 26014 34914 26066 34926
rect 28366 34914 28418 34926
rect 28130 34862 28142 34914
rect 28194 34862 28206 34914
rect 26014 34850 26066 34862
rect 28366 34850 28418 34862
rect 29038 34914 29090 34926
rect 29038 34850 29090 34862
rect 29374 34914 29426 34926
rect 29374 34850 29426 34862
rect 35086 34914 35138 34926
rect 35086 34850 35138 34862
rect 35646 34914 35698 34926
rect 35646 34850 35698 34862
rect 14814 34802 14866 34814
rect 14814 34738 14866 34750
rect 18398 34802 18450 34814
rect 18398 34738 18450 34750
rect 19518 34802 19570 34814
rect 19518 34738 19570 34750
rect 19966 34802 20018 34814
rect 19966 34738 20018 34750
rect 20078 34802 20130 34814
rect 20078 34738 20130 34750
rect 26238 34802 26290 34814
rect 26238 34738 26290 34750
rect 27470 34802 27522 34814
rect 27470 34738 27522 34750
rect 37326 34802 37378 34814
rect 37326 34738 37378 34750
rect 40238 34802 40290 34814
rect 40238 34738 40290 34750
rect 40350 34802 40402 34814
rect 40350 34738 40402 34750
rect 40798 34802 40850 34814
rect 40798 34738 40850 34750
rect 14590 34690 14642 34702
rect 29262 34690 29314 34702
rect 18946 34638 18958 34690
rect 19010 34638 19022 34690
rect 21634 34638 21646 34690
rect 21698 34638 21710 34690
rect 14590 34626 14642 34638
rect 29262 34626 29314 34638
rect 37438 34690 37490 34702
rect 37438 34626 37490 34638
rect 40574 34690 40626 34702
rect 40574 34626 40626 34638
rect 40910 34690 40962 34702
rect 40910 34626 40962 34638
rect 1344 34522 44576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 44576 34522
rect 1344 34436 44576 34470
rect 13918 34354 13970 34366
rect 19070 34354 19122 34366
rect 14242 34302 14254 34354
rect 14306 34302 14318 34354
rect 13918 34290 13970 34302
rect 19070 34290 19122 34302
rect 19182 34242 19234 34254
rect 37426 34190 37438 34242
rect 37490 34190 37502 34242
rect 19182 34178 19234 34190
rect 37102 34130 37154 34142
rect 41234 34078 41246 34130
rect 41298 34078 41310 34130
rect 37102 34066 37154 34078
rect 36766 34018 36818 34030
rect 36766 33954 36818 33966
rect 40350 34018 40402 34030
rect 41906 33966 41918 34018
rect 41970 33966 41982 34018
rect 44034 33966 44046 34018
rect 44098 33966 44110 34018
rect 40350 33954 40402 33966
rect 1344 33738 44576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 44576 33738
rect 1344 33652 44576 33686
rect 41246 33570 41298 33582
rect 41246 33506 41298 33518
rect 6626 33406 6638 33458
rect 6690 33406 6702 33458
rect 33618 33406 33630 33458
rect 33682 33406 33694 33458
rect 10334 33346 10386 33358
rect 9538 33294 9550 33346
rect 9602 33294 9614 33346
rect 10334 33282 10386 33294
rect 11006 33346 11058 33358
rect 33182 33346 33234 33358
rect 29362 33294 29374 33346
rect 29426 33294 29438 33346
rect 11006 33282 11058 33294
rect 33182 33282 33234 33294
rect 34078 33346 34130 33358
rect 34078 33282 34130 33294
rect 40574 33346 40626 33358
rect 41358 33346 41410 33358
rect 40898 33294 40910 33346
rect 40962 33294 40974 33346
rect 40574 33282 40626 33294
rect 41358 33282 41410 33294
rect 41582 33234 41634 33246
rect 8754 33182 8766 33234
rect 8818 33182 8830 33234
rect 34402 33182 34414 33234
rect 34466 33182 34478 33234
rect 41582 33170 41634 33182
rect 41694 33234 41746 33246
rect 41694 33170 41746 33182
rect 42142 33234 42194 33246
rect 42142 33170 42194 33182
rect 9998 33122 10050 33134
rect 9998 33058 10050 33070
rect 10446 33122 10498 33134
rect 10446 33058 10498 33070
rect 10558 33122 10610 33134
rect 10558 33058 10610 33070
rect 11454 33122 11506 33134
rect 40462 33122 40514 33134
rect 29138 33070 29150 33122
rect 29202 33070 29214 33122
rect 11454 33058 11506 33070
rect 40462 33058 40514 33070
rect 41134 33122 41186 33134
rect 41134 33058 41186 33070
rect 1344 32954 44576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 44576 32954
rect 1344 32868 44576 32902
rect 8318 32786 8370 32798
rect 8318 32722 8370 32734
rect 9774 32786 9826 32798
rect 9774 32722 9826 32734
rect 24334 32786 24386 32798
rect 24334 32722 24386 32734
rect 8430 32674 8482 32686
rect 8430 32610 8482 32622
rect 8990 32674 9042 32686
rect 8990 32610 9042 32622
rect 24222 32674 24274 32686
rect 24222 32610 24274 32622
rect 25230 32674 25282 32686
rect 32498 32622 32510 32674
rect 32562 32622 32574 32674
rect 25230 32610 25282 32622
rect 25342 32562 25394 32574
rect 2706 32510 2718 32562
rect 2770 32510 2782 32562
rect 8082 32510 8094 32562
rect 8146 32510 8158 32562
rect 25342 32498 25394 32510
rect 25454 32562 25506 32574
rect 25454 32498 25506 32510
rect 25678 32562 25730 32574
rect 36430 32562 36482 32574
rect 32274 32510 32286 32562
rect 32338 32510 32350 32562
rect 33170 32510 33182 32562
rect 33234 32510 33246 32562
rect 25678 32498 25730 32510
rect 36430 32498 36482 32510
rect 5966 32450 6018 32462
rect 3378 32398 3390 32450
rect 3442 32398 3454 32450
rect 5506 32398 5518 32450
rect 5570 32398 5582 32450
rect 5966 32386 6018 32398
rect 10334 32450 10386 32462
rect 33842 32398 33854 32450
rect 33906 32398 33918 32450
rect 35970 32398 35982 32450
rect 36034 32398 36046 32450
rect 10334 32386 10386 32398
rect 8878 32338 8930 32350
rect 8878 32274 8930 32286
rect 24446 32338 24498 32350
rect 24446 32274 24498 32286
rect 1344 32170 44576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 44576 32170
rect 1344 32084 44576 32118
rect 16830 31890 16882 31902
rect 5058 31838 5070 31890
rect 5122 31838 5134 31890
rect 13458 31838 13470 31890
rect 13522 31838 13534 31890
rect 16830 31826 16882 31838
rect 24894 31890 24946 31902
rect 33394 31838 33406 31890
rect 33458 31838 33470 31890
rect 24894 31826 24946 31838
rect 33854 31778 33906 31790
rect 2258 31726 2270 31778
rect 2322 31726 2334 31778
rect 16370 31726 16382 31778
rect 16434 31726 16446 31778
rect 24994 31726 25006 31778
rect 25058 31726 25070 31778
rect 33854 31714 33906 31726
rect 34302 31778 34354 31790
rect 34302 31714 34354 31726
rect 39342 31778 39394 31790
rect 39342 31714 39394 31726
rect 24110 31666 24162 31678
rect 2930 31614 2942 31666
rect 2994 31614 3006 31666
rect 15586 31614 15598 31666
rect 15650 31614 15662 31666
rect 24110 31602 24162 31614
rect 24446 31666 24498 31678
rect 24446 31602 24498 31614
rect 24782 31666 24834 31678
rect 24782 31602 24834 31614
rect 25230 31666 25282 31678
rect 25230 31602 25282 31614
rect 32958 31666 33010 31678
rect 32958 31602 33010 31614
rect 33294 31666 33346 31678
rect 33294 31602 33346 31614
rect 33966 31666 34018 31678
rect 33966 31602 34018 31614
rect 34638 31666 34690 31678
rect 34638 31602 34690 31614
rect 34750 31666 34802 31678
rect 38782 31666 38834 31678
rect 37314 31614 37326 31666
rect 37378 31614 37390 31666
rect 34750 31602 34802 31614
rect 38782 31602 38834 31614
rect 39006 31666 39058 31678
rect 39006 31602 39058 31614
rect 5742 31554 5794 31566
rect 5742 31490 5794 31502
rect 33518 31554 33570 31566
rect 33518 31490 33570 31502
rect 34190 31554 34242 31566
rect 34190 31490 34242 31502
rect 34974 31554 35026 31566
rect 34974 31490 35026 31502
rect 36542 31554 36594 31566
rect 36542 31490 36594 31502
rect 36990 31554 37042 31566
rect 36990 31490 37042 31502
rect 39230 31554 39282 31566
rect 39230 31490 39282 31502
rect 1344 31386 44576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 44576 31386
rect 1344 31300 44576 31334
rect 15822 31218 15874 31230
rect 15822 31154 15874 31166
rect 24222 31218 24274 31230
rect 24222 31154 24274 31166
rect 24446 31106 24498 31118
rect 10434 31054 10446 31106
rect 10498 31054 10510 31106
rect 24446 31042 24498 31054
rect 24558 31106 24610 31118
rect 24558 31042 24610 31054
rect 32622 30994 32674 31006
rect 15474 30942 15486 30994
rect 15538 30942 15550 30994
rect 21410 30942 21422 30994
rect 21474 30942 21486 30994
rect 30258 30942 30270 30994
rect 30322 30942 30334 30994
rect 33170 30942 33182 30994
rect 33234 30942 33246 30994
rect 32622 30930 32674 30942
rect 15934 30882 15986 30894
rect 15934 30818 15986 30830
rect 16494 30882 16546 30894
rect 16494 30818 16546 30830
rect 18286 30882 18338 30894
rect 23998 30882 24050 30894
rect 30718 30882 30770 30894
rect 18610 30830 18622 30882
rect 18674 30830 18686 30882
rect 20738 30830 20750 30882
rect 20802 30830 20814 30882
rect 27346 30830 27358 30882
rect 27410 30830 27422 30882
rect 29474 30830 29486 30882
rect 29538 30830 29550 30882
rect 36866 30830 36878 30882
rect 36930 30830 36942 30882
rect 18286 30818 18338 30830
rect 23998 30818 24050 30830
rect 30718 30818 30770 30830
rect 1344 30602 44576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 44576 30602
rect 1344 30516 44576 30550
rect 8766 30434 8818 30446
rect 8766 30370 8818 30382
rect 9102 30322 9154 30334
rect 16818 30270 16830 30322
rect 16882 30270 16894 30322
rect 24546 30270 24558 30322
rect 24610 30270 24622 30322
rect 37426 30270 37438 30322
rect 37490 30270 37502 30322
rect 39554 30270 39566 30322
rect 39618 30270 39630 30322
rect 9102 30258 9154 30270
rect 9662 30210 9714 30222
rect 10670 30210 10722 30222
rect 37102 30210 37154 30222
rect 8754 30158 8766 30210
rect 8818 30158 8830 30210
rect 10098 30158 10110 30210
rect 10162 30158 10174 30210
rect 13570 30158 13582 30210
rect 13634 30158 13646 30210
rect 16034 30158 16046 30210
rect 16098 30158 16110 30210
rect 24882 30158 24894 30210
rect 24946 30158 24958 30210
rect 28130 30158 28142 30210
rect 28194 30158 28206 30210
rect 28354 30158 28366 30210
rect 28418 30158 28430 30210
rect 29362 30158 29374 30210
rect 29426 30158 29438 30210
rect 40338 30158 40350 30210
rect 40402 30158 40414 30210
rect 9662 30146 9714 30158
rect 10670 30146 10722 30158
rect 37102 30146 37154 30158
rect 14030 30098 14082 30110
rect 14030 30034 14082 30046
rect 25342 30098 25394 30110
rect 25342 30034 25394 30046
rect 28590 30098 28642 30110
rect 42702 30098 42754 30110
rect 31378 30046 31390 30098
rect 31442 30046 31454 30098
rect 28590 30034 28642 30046
rect 42702 30034 42754 30046
rect 20302 29986 20354 29998
rect 20302 29922 20354 29934
rect 42590 29986 42642 29998
rect 42590 29922 42642 29934
rect 1344 29818 44576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 44576 29818
rect 1344 29732 44576 29766
rect 5070 29650 5122 29662
rect 5070 29586 5122 29598
rect 17502 29650 17554 29662
rect 17502 29586 17554 29598
rect 18622 29650 18674 29662
rect 18622 29586 18674 29598
rect 18958 29650 19010 29662
rect 18958 29586 19010 29598
rect 19630 29650 19682 29662
rect 19630 29586 19682 29598
rect 28366 29650 28418 29662
rect 28366 29586 28418 29598
rect 29934 29650 29986 29662
rect 29934 29586 29986 29598
rect 33182 29650 33234 29662
rect 33182 29586 33234 29598
rect 37550 29650 37602 29662
rect 37550 29586 37602 29598
rect 38782 29650 38834 29662
rect 38782 29586 38834 29598
rect 38894 29650 38946 29662
rect 38894 29586 38946 29598
rect 39118 29650 39170 29662
rect 39118 29586 39170 29598
rect 40350 29650 40402 29662
rect 40350 29586 40402 29598
rect 5630 29538 5682 29550
rect 5630 29474 5682 29486
rect 8654 29538 8706 29550
rect 14478 29538 14530 29550
rect 10770 29486 10782 29538
rect 10834 29486 10846 29538
rect 8654 29474 8706 29486
rect 14478 29474 14530 29486
rect 15486 29538 15538 29550
rect 15486 29474 15538 29486
rect 16158 29538 16210 29550
rect 16158 29474 16210 29486
rect 17614 29538 17666 29550
rect 17614 29474 17666 29486
rect 19854 29538 19906 29550
rect 19854 29474 19906 29486
rect 25230 29538 25282 29550
rect 25230 29474 25282 29486
rect 29150 29538 29202 29550
rect 29150 29474 29202 29486
rect 29374 29538 29426 29550
rect 29374 29474 29426 29486
rect 33070 29538 33122 29550
rect 37662 29538 37714 29550
rect 36642 29486 36654 29538
rect 36706 29486 36718 29538
rect 33070 29474 33122 29486
rect 37662 29474 37714 29486
rect 38670 29538 38722 29550
rect 38670 29474 38722 29486
rect 3726 29426 3778 29438
rect 3726 29362 3778 29374
rect 3950 29426 4002 29438
rect 3950 29362 4002 29374
rect 4398 29426 4450 29438
rect 4398 29362 4450 29374
rect 4622 29426 4674 29438
rect 4622 29362 4674 29374
rect 4846 29426 4898 29438
rect 4846 29362 4898 29374
rect 5182 29426 5234 29438
rect 5182 29362 5234 29374
rect 8990 29426 9042 29438
rect 11454 29426 11506 29438
rect 9986 29374 9998 29426
rect 10050 29374 10062 29426
rect 10546 29374 10558 29426
rect 10610 29374 10622 29426
rect 8990 29362 9042 29374
rect 11454 29362 11506 29374
rect 11902 29426 11954 29438
rect 11902 29362 11954 29374
rect 12126 29426 12178 29438
rect 12126 29362 12178 29374
rect 14366 29426 14418 29438
rect 14366 29362 14418 29374
rect 16270 29426 16322 29438
rect 16270 29362 16322 29374
rect 16382 29426 16434 29438
rect 16382 29362 16434 29374
rect 17390 29426 17442 29438
rect 18846 29426 18898 29438
rect 17826 29374 17838 29426
rect 17890 29374 17902 29426
rect 18050 29374 18062 29426
rect 18114 29374 18126 29426
rect 17390 29362 17442 29374
rect 18846 29362 18898 29374
rect 19070 29426 19122 29438
rect 19070 29362 19122 29374
rect 19294 29426 19346 29438
rect 36318 29426 36370 29438
rect 25554 29374 25566 29426
rect 25618 29374 25630 29426
rect 41122 29374 41134 29426
rect 41186 29374 41198 29426
rect 19294 29362 19346 29374
rect 36318 29362 36370 29374
rect 3838 29314 3890 29326
rect 3838 29250 3890 29262
rect 6078 29314 6130 29326
rect 15598 29314 15650 29326
rect 19966 29314 20018 29326
rect 9650 29262 9662 29314
rect 9714 29262 9726 29314
rect 12674 29262 12686 29314
rect 12738 29262 12750 29314
rect 16818 29262 16830 29314
rect 16882 29262 16894 29314
rect 6078 29250 6130 29262
rect 15598 29250 15650 29262
rect 19966 29250 20018 29262
rect 20302 29314 20354 29326
rect 20302 29250 20354 29262
rect 25342 29314 25394 29326
rect 25342 29250 25394 29262
rect 26014 29314 26066 29326
rect 26014 29250 26066 29262
rect 28814 29314 28866 29326
rect 35982 29314 36034 29326
rect 29474 29262 29486 29314
rect 29538 29262 29550 29314
rect 41906 29262 41918 29314
rect 41970 29262 41982 29314
rect 44034 29262 44046 29314
rect 44098 29262 44110 29314
rect 28814 29250 28866 29262
rect 35982 29250 36034 29262
rect 5518 29202 5570 29214
rect 5518 29138 5570 29150
rect 11678 29202 11730 29214
rect 11678 29138 11730 29150
rect 15710 29202 15762 29214
rect 15710 29138 15762 29150
rect 33182 29202 33234 29214
rect 33182 29138 33234 29150
rect 37550 29202 37602 29214
rect 37550 29138 37602 29150
rect 1344 29034 44576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 44576 29034
rect 1344 28948 44576 28982
rect 3278 28866 3330 28878
rect 3278 28802 3330 28814
rect 4286 28866 4338 28878
rect 4286 28802 4338 28814
rect 5182 28866 5234 28878
rect 5182 28802 5234 28814
rect 6414 28866 6466 28878
rect 6414 28802 6466 28814
rect 9662 28866 9714 28878
rect 41234 28814 41246 28866
rect 41298 28814 41310 28866
rect 9662 28802 9714 28814
rect 6974 28754 7026 28766
rect 6974 28690 7026 28702
rect 17278 28754 17330 28766
rect 17278 28690 17330 28702
rect 18398 28754 18450 28766
rect 35086 28754 35138 28766
rect 23538 28702 23550 28754
rect 23602 28702 23614 28754
rect 25666 28702 25678 28754
rect 25730 28702 25742 28754
rect 31042 28702 31054 28754
rect 31106 28702 31118 28754
rect 33170 28702 33182 28754
rect 33234 28702 33246 28754
rect 18398 28690 18450 28702
rect 35086 28690 35138 28702
rect 40014 28754 40066 28766
rect 40014 28690 40066 28702
rect 40462 28754 40514 28766
rect 40462 28690 40514 28702
rect 41694 28754 41746 28766
rect 41694 28690 41746 28702
rect 4510 28642 4562 28654
rect 3154 28590 3166 28642
rect 3218 28590 3230 28642
rect 4510 28578 4562 28590
rect 4734 28642 4786 28654
rect 4734 28578 4786 28590
rect 5966 28642 6018 28654
rect 5966 28578 6018 28590
rect 7982 28642 8034 28654
rect 7982 28578 8034 28590
rect 8766 28642 8818 28654
rect 8766 28578 8818 28590
rect 8878 28642 8930 28654
rect 12574 28642 12626 28654
rect 9202 28590 9214 28642
rect 9266 28590 9278 28642
rect 9874 28590 9886 28642
rect 9938 28590 9950 28642
rect 10434 28590 10446 28642
rect 10498 28590 10510 28642
rect 11218 28590 11230 28642
rect 11282 28590 11294 28642
rect 11554 28590 11566 28642
rect 11618 28590 11630 28642
rect 8878 28578 8930 28590
rect 12574 28578 12626 28590
rect 13470 28642 13522 28654
rect 16270 28642 16322 28654
rect 13906 28590 13918 28642
rect 13970 28590 13982 28642
rect 16034 28590 16046 28642
rect 16098 28590 16110 28642
rect 13470 28578 13522 28590
rect 16270 28578 16322 28590
rect 16382 28642 16434 28654
rect 26126 28642 26178 28654
rect 33742 28642 33794 28654
rect 22866 28590 22878 28642
rect 22930 28590 22942 28642
rect 30258 28590 30270 28642
rect 30322 28590 30334 28642
rect 16382 28578 16434 28590
rect 26126 28578 26178 28590
rect 33742 28578 33794 28590
rect 33966 28642 34018 28654
rect 33966 28578 34018 28590
rect 34190 28642 34242 28654
rect 34190 28578 34242 28590
rect 35422 28642 35474 28654
rect 41470 28642 41522 28654
rect 41122 28590 41134 28642
rect 41186 28590 41198 28642
rect 35422 28578 35474 28590
rect 41470 28578 41522 28590
rect 3726 28530 3778 28542
rect 3490 28478 3502 28530
rect 3554 28478 3566 28530
rect 3726 28466 3778 28478
rect 4062 28530 4114 28542
rect 4062 28466 4114 28478
rect 6414 28530 6466 28542
rect 6414 28466 6466 28478
rect 6526 28530 6578 28542
rect 6526 28466 6578 28478
rect 8318 28530 8370 28542
rect 10782 28530 10834 28542
rect 33518 28530 33570 28542
rect 41806 28530 41858 28542
rect 9090 28478 9102 28530
rect 9154 28478 9166 28530
rect 12002 28478 12014 28530
rect 12066 28478 12078 28530
rect 35746 28478 35758 28530
rect 35810 28478 35822 28530
rect 8318 28466 8370 28478
rect 10782 28466 10834 28478
rect 33518 28466 33570 28478
rect 41806 28466 41858 28478
rect 2942 28418 2994 28430
rect 7870 28418 7922 28430
rect 5618 28366 5630 28418
rect 5682 28366 5694 28418
rect 2942 28354 2994 28366
rect 7870 28354 7922 28366
rect 8206 28418 8258 28430
rect 16818 28366 16830 28418
rect 16882 28366 16894 28418
rect 8206 28354 8258 28366
rect 1344 28250 44576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 44576 28250
rect 1344 28164 44576 28198
rect 3614 28082 3666 28094
rect 3614 28018 3666 28030
rect 4510 28082 4562 28094
rect 4510 28018 4562 28030
rect 4622 28082 4674 28094
rect 4622 28018 4674 28030
rect 5070 28082 5122 28094
rect 5070 28018 5122 28030
rect 10558 28082 10610 28094
rect 10558 28018 10610 28030
rect 10894 28082 10946 28094
rect 10894 28018 10946 28030
rect 18174 28082 18226 28094
rect 18174 28018 18226 28030
rect 41358 28082 41410 28094
rect 41358 28018 41410 28030
rect 5406 27970 5458 27982
rect 17390 27970 17442 27982
rect 4162 27918 4174 27970
rect 4226 27918 4238 27970
rect 9986 27918 9998 27970
rect 10050 27918 10062 27970
rect 5406 27906 5458 27918
rect 17390 27906 17442 27918
rect 18062 27970 18114 27982
rect 18062 27906 18114 27918
rect 4734 27858 4786 27870
rect 4274 27806 4286 27858
rect 4338 27806 4350 27858
rect 4734 27794 4786 27806
rect 9550 27858 9602 27870
rect 9550 27794 9602 27806
rect 9774 27858 9826 27870
rect 17614 27858 17666 27870
rect 10098 27806 10110 27858
rect 10162 27806 10174 27858
rect 9774 27794 9826 27806
rect 17614 27794 17666 27806
rect 17838 27858 17890 27870
rect 17838 27794 17890 27806
rect 40350 27858 40402 27870
rect 41122 27806 41134 27858
rect 41186 27806 41198 27858
rect 40350 27794 40402 27806
rect 15486 27746 15538 27758
rect 15486 27682 15538 27694
rect 21870 27746 21922 27758
rect 21870 27682 21922 27694
rect 33182 27746 33234 27758
rect 33182 27682 33234 27694
rect 33630 27746 33682 27758
rect 33630 27682 33682 27694
rect 41470 27634 41522 27646
rect 41470 27570 41522 27582
rect 1344 27466 44576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 44576 27466
rect 1344 27380 44576 27414
rect 14142 27186 14194 27198
rect 15822 27186 15874 27198
rect 20302 27186 20354 27198
rect 25454 27186 25506 27198
rect 15026 27134 15038 27186
rect 15090 27134 15102 27186
rect 16146 27134 16158 27186
rect 16210 27134 16222 27186
rect 21746 27134 21758 27186
rect 21810 27134 21822 27186
rect 14142 27122 14194 27134
rect 15822 27122 15874 27134
rect 20302 27122 20354 27134
rect 25454 27122 25506 27134
rect 26350 27186 26402 27198
rect 26350 27122 26402 27134
rect 36430 27186 36482 27198
rect 41470 27186 41522 27198
rect 39890 27134 39902 27186
rect 39954 27134 39966 27186
rect 41010 27134 41022 27186
rect 41074 27134 41086 27186
rect 36430 27122 36482 27134
rect 41470 27122 41522 27134
rect 17166 27074 17218 27086
rect 22542 27074 22594 27086
rect 35422 27074 35474 27086
rect 14914 27022 14926 27074
rect 14978 27022 14990 27074
rect 15250 27022 15262 27074
rect 15314 27022 15326 27074
rect 17714 27022 17726 27074
rect 17778 27022 17790 27074
rect 25890 27022 25902 27074
rect 25954 27022 25966 27074
rect 17166 27010 17218 27022
rect 22542 27010 22594 27022
rect 35422 27010 35474 27022
rect 37102 27074 37154 27086
rect 40786 27022 40798 27074
rect 40850 27022 40862 27074
rect 37102 27010 37154 27022
rect 20526 26962 20578 26974
rect 14466 26910 14478 26962
rect 14530 26910 14542 26962
rect 20526 26898 20578 26910
rect 20638 26962 20690 26974
rect 20638 26898 20690 26910
rect 21310 26962 21362 26974
rect 29710 26962 29762 26974
rect 22194 26910 22206 26962
rect 22258 26910 22270 26962
rect 29362 26910 29374 26962
rect 29426 26910 29438 26962
rect 21310 26898 21362 26910
rect 29710 26898 29762 26910
rect 30270 26962 30322 26974
rect 30270 26898 30322 26910
rect 39454 26962 39506 26974
rect 39454 26898 39506 26910
rect 17278 26850 17330 26862
rect 17278 26786 17330 26798
rect 17390 26850 17442 26862
rect 17390 26786 17442 26798
rect 20862 26850 20914 26862
rect 20862 26786 20914 26798
rect 35086 26850 35138 26862
rect 35086 26786 35138 26798
rect 35310 26850 35362 26862
rect 37426 26798 37438 26850
rect 37490 26798 37502 26850
rect 35310 26786 35362 26798
rect 1344 26682 44576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 44576 26682
rect 1344 26596 44576 26630
rect 6638 26514 6690 26526
rect 18846 26514 18898 26526
rect 14354 26462 14366 26514
rect 14418 26462 14430 26514
rect 6638 26450 6690 26462
rect 18846 26450 18898 26462
rect 19854 26514 19906 26526
rect 19854 26450 19906 26462
rect 37214 26514 37266 26526
rect 37214 26450 37266 26462
rect 37662 26514 37714 26526
rect 37662 26450 37714 26462
rect 3838 26402 3890 26414
rect 3838 26338 3890 26350
rect 6414 26402 6466 26414
rect 17726 26402 17778 26414
rect 10770 26350 10782 26402
rect 10834 26350 10846 26402
rect 14466 26350 14478 26402
rect 14530 26350 14542 26402
rect 15250 26350 15262 26402
rect 15314 26350 15326 26402
rect 15810 26350 15822 26402
rect 15874 26350 15886 26402
rect 20962 26350 20974 26402
rect 21026 26350 21038 26402
rect 6414 26338 6466 26350
rect 17726 26338 17778 26350
rect 5966 26290 6018 26302
rect 16046 26290 16098 26302
rect 17614 26290 17666 26302
rect 18734 26290 18786 26302
rect 12226 26238 12238 26290
rect 12290 26238 12302 26290
rect 12674 26238 12686 26290
rect 12738 26238 12750 26290
rect 17378 26238 17390 26290
rect 17442 26238 17454 26290
rect 18162 26238 18174 26290
rect 18226 26238 18238 26290
rect 18498 26238 18510 26290
rect 18562 26238 18574 26290
rect 5966 26226 6018 26238
rect 16046 26226 16098 26238
rect 17614 26226 17666 26238
rect 18734 26226 18786 26238
rect 18958 26290 19010 26302
rect 37438 26290 37490 26302
rect 19170 26238 19182 26290
rect 19234 26238 19246 26290
rect 20178 26238 20190 26290
rect 20242 26238 20254 26290
rect 26786 26238 26798 26290
rect 26850 26238 26862 26290
rect 33954 26238 33966 26290
rect 34018 26238 34030 26290
rect 18958 26226 19010 26238
rect 37438 26226 37490 26238
rect 6526 26178 6578 26190
rect 6526 26114 6578 26126
rect 16158 26178 16210 26190
rect 30046 26178 30098 26190
rect 37326 26178 37378 26190
rect 23090 26126 23102 26178
rect 23154 26126 23166 26178
rect 27458 26126 27470 26178
rect 27522 26126 27534 26178
rect 29586 26126 29598 26178
rect 29650 26126 29662 26178
rect 34738 26126 34750 26178
rect 34802 26126 34814 26178
rect 36866 26126 36878 26178
rect 36930 26126 36942 26178
rect 16158 26114 16210 26126
rect 30046 26114 30098 26126
rect 37326 26114 37378 26126
rect 40126 26178 40178 26190
rect 40126 26114 40178 26126
rect 3726 26066 3778 26078
rect 3726 26002 3778 26014
rect 1344 25898 44576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 44576 25898
rect 1344 25812 44576 25846
rect 12238 25730 12290 25742
rect 6290 25678 6302 25730
rect 6354 25727 6366 25730
rect 6514 25727 6526 25730
rect 6354 25681 6526 25727
rect 6354 25678 6366 25681
rect 6514 25678 6526 25681
rect 6578 25678 6590 25730
rect 12238 25666 12290 25678
rect 12462 25730 12514 25742
rect 17602 25678 17614 25730
rect 17666 25678 17678 25730
rect 12462 25666 12514 25678
rect 8878 25618 8930 25630
rect 8878 25554 8930 25566
rect 27134 25618 27186 25630
rect 27134 25554 27186 25566
rect 27582 25618 27634 25630
rect 27582 25554 27634 25566
rect 34974 25618 35026 25630
rect 34974 25554 35026 25566
rect 35422 25618 35474 25630
rect 35422 25554 35474 25566
rect 37214 25618 37266 25630
rect 37214 25554 37266 25566
rect 39902 25618 39954 25630
rect 44034 25566 44046 25618
rect 44098 25566 44110 25618
rect 39902 25554 39954 25566
rect 5518 25506 5570 25518
rect 5518 25442 5570 25454
rect 5966 25506 6018 25518
rect 11790 25506 11842 25518
rect 8642 25454 8654 25506
rect 8706 25454 8718 25506
rect 5966 25442 6018 25454
rect 11790 25442 11842 25454
rect 12686 25506 12738 25518
rect 24894 25506 24946 25518
rect 29374 25506 29426 25518
rect 35198 25506 35250 25518
rect 14354 25454 14366 25506
rect 14418 25454 14430 25506
rect 15586 25454 15598 25506
rect 15650 25454 15662 25506
rect 17490 25454 17502 25506
rect 17554 25454 17566 25506
rect 24210 25454 24222 25506
rect 24274 25454 24286 25506
rect 28242 25454 28254 25506
rect 28306 25454 28318 25506
rect 29698 25454 29710 25506
rect 29762 25454 29774 25506
rect 12686 25442 12738 25454
rect 24894 25442 24946 25454
rect 29374 25442 29426 25454
rect 35198 25442 35250 25454
rect 35870 25506 35922 25518
rect 35870 25442 35922 25454
rect 40014 25506 40066 25518
rect 40014 25442 40066 25454
rect 40462 25506 40514 25518
rect 41122 25454 41134 25506
rect 41186 25454 41198 25506
rect 40462 25442 40514 25454
rect 6190 25394 6242 25406
rect 6190 25330 6242 25342
rect 8990 25394 9042 25406
rect 8990 25330 9042 25342
rect 12910 25394 12962 25406
rect 18174 25394 18226 25406
rect 17154 25342 17166 25394
rect 17218 25342 17230 25394
rect 12910 25330 12962 25342
rect 18174 25330 18226 25342
rect 24446 25394 24498 25406
rect 24446 25330 24498 25342
rect 27806 25394 27858 25406
rect 27806 25330 27858 25342
rect 29262 25394 29314 25406
rect 29262 25330 29314 25342
rect 35646 25394 35698 25406
rect 35646 25330 35698 25342
rect 40686 25394 40738 25406
rect 41906 25342 41918 25394
rect 41970 25342 41982 25394
rect 40686 25330 40738 25342
rect 5742 25282 5794 25294
rect 5742 25218 5794 25230
rect 6750 25282 6802 25294
rect 6750 25218 6802 25230
rect 27470 25282 27522 25294
rect 27470 25218 27522 25230
rect 27694 25282 27746 25294
rect 27694 25218 27746 25230
rect 29150 25282 29202 25294
rect 29150 25218 29202 25230
rect 30158 25282 30210 25294
rect 30158 25218 30210 25230
rect 40574 25282 40626 25294
rect 40574 25218 40626 25230
rect 1344 25114 44576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 44576 25114
rect 1344 25028 44576 25062
rect 18958 24946 19010 24958
rect 16034 24894 16046 24946
rect 16098 24894 16110 24946
rect 18958 24882 19010 24894
rect 28926 24946 28978 24958
rect 28926 24882 28978 24894
rect 38222 24946 38274 24958
rect 38222 24882 38274 24894
rect 41358 24946 41410 24958
rect 41358 24882 41410 24894
rect 40910 24834 40962 24846
rect 12450 24782 12462 24834
rect 12514 24782 12526 24834
rect 16146 24782 16158 24834
rect 16210 24782 16222 24834
rect 40910 24770 40962 24782
rect 7646 24722 7698 24734
rect 7646 24658 7698 24670
rect 8206 24722 8258 24734
rect 14478 24722 14530 24734
rect 12338 24670 12350 24722
rect 12402 24670 12414 24722
rect 8206 24658 8258 24670
rect 14478 24658 14530 24670
rect 32510 24722 32562 24734
rect 32510 24658 32562 24670
rect 33182 24722 33234 24734
rect 33182 24658 33234 24670
rect 33406 24722 33458 24734
rect 33406 24658 33458 24670
rect 33742 24722 33794 24734
rect 33742 24658 33794 24670
rect 38446 24722 38498 24734
rect 41246 24722 41298 24734
rect 38770 24670 38782 24722
rect 38834 24670 38846 24722
rect 38446 24658 38498 24670
rect 41246 24658 41298 24670
rect 41582 24722 41634 24734
rect 41582 24658 41634 24670
rect 28478 24610 28530 24622
rect 28478 24546 28530 24558
rect 33518 24610 33570 24622
rect 33518 24546 33570 24558
rect 38334 24610 38386 24622
rect 38334 24546 38386 24558
rect 40350 24610 40402 24622
rect 40350 24546 40402 24558
rect 1344 24330 44576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 44576 24330
rect 1344 24244 44576 24278
rect 35758 24162 35810 24174
rect 29698 24110 29710 24162
rect 29762 24159 29774 24162
rect 29922 24159 29934 24162
rect 29762 24113 29934 24159
rect 29762 24110 29774 24113
rect 29922 24110 29934 24113
rect 29986 24110 29998 24162
rect 35758 24098 35810 24110
rect 6414 24050 6466 24062
rect 2930 23998 2942 24050
rect 2994 23998 3006 24050
rect 5058 23998 5070 24050
rect 5122 23998 5134 24050
rect 6414 23986 6466 23998
rect 7310 24050 7362 24062
rect 7310 23986 7362 23998
rect 16942 24050 16994 24062
rect 16942 23986 16994 23998
rect 23438 24050 23490 24062
rect 23438 23986 23490 23998
rect 23886 24050 23938 24062
rect 23886 23986 23938 23998
rect 29934 24050 29986 24062
rect 34302 24050 34354 24062
rect 31714 23998 31726 24050
rect 31778 23998 31790 24050
rect 33842 23998 33854 24050
rect 33906 23998 33918 24050
rect 29934 23986 29986 23998
rect 34302 23986 34354 23998
rect 35534 24050 35586 24062
rect 35534 23986 35586 23998
rect 35870 24050 35922 24062
rect 35870 23986 35922 23998
rect 5854 23938 5906 23950
rect 19294 23938 19346 23950
rect 2258 23886 2270 23938
rect 2322 23886 2334 23938
rect 6850 23886 6862 23938
rect 6914 23886 6926 23938
rect 10770 23886 10782 23938
rect 10834 23886 10846 23938
rect 11106 23886 11118 23938
rect 11170 23886 11182 23938
rect 15138 23886 15150 23938
rect 15202 23886 15214 23938
rect 17154 23886 17166 23938
rect 17218 23886 17230 23938
rect 5854 23874 5906 23886
rect 19294 23874 19346 23886
rect 22878 23938 22930 23950
rect 24894 23938 24946 23950
rect 24322 23886 24334 23938
rect 24386 23886 24398 23938
rect 29250 23886 29262 23938
rect 29314 23886 29326 23938
rect 31042 23886 31054 23938
rect 31106 23886 31118 23938
rect 22878 23874 22930 23886
rect 24894 23874 24946 23886
rect 16270 23826 16322 23838
rect 11666 23774 11678 23826
rect 11730 23774 11742 23826
rect 16270 23762 16322 23774
rect 17726 23826 17778 23838
rect 17726 23762 17778 23774
rect 22766 23826 22818 23838
rect 22766 23762 22818 23774
rect 7422 23714 7474 23726
rect 7422 23650 7474 23662
rect 10446 23714 10498 23726
rect 22542 23714 22594 23726
rect 11330 23662 11342 23714
rect 11394 23662 11406 23714
rect 19618 23662 19630 23714
rect 19682 23662 19694 23714
rect 10446 23650 10498 23662
rect 22542 23650 22594 23662
rect 24558 23714 24610 23726
rect 40686 23714 40738 23726
rect 25218 23662 25230 23714
rect 25282 23662 25294 23714
rect 29474 23662 29486 23714
rect 29538 23662 29550 23714
rect 24558 23650 24610 23662
rect 40686 23650 40738 23662
rect 1344 23546 44576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 44576 23546
rect 1344 23460 44576 23494
rect 15934 23378 15986 23390
rect 21534 23378 21586 23390
rect 19058 23326 19070 23378
rect 19122 23326 19134 23378
rect 15934 23314 15986 23326
rect 21534 23314 21586 23326
rect 22654 23378 22706 23390
rect 33406 23378 33458 23390
rect 26674 23326 26686 23378
rect 26738 23326 26750 23378
rect 22654 23314 22706 23326
rect 33406 23314 33458 23326
rect 39118 23378 39170 23390
rect 41458 23326 41470 23378
rect 41522 23326 41534 23378
rect 39118 23314 39170 23326
rect 33070 23266 33122 23278
rect 3154 23214 3166 23266
rect 3218 23214 3230 23266
rect 19170 23214 19182 23266
rect 19234 23214 19246 23266
rect 21074 23214 21086 23266
rect 21138 23214 21150 23266
rect 29138 23214 29150 23266
rect 29202 23214 29214 23266
rect 33070 23202 33122 23214
rect 33182 23266 33234 23278
rect 33182 23202 33234 23214
rect 35870 23266 35922 23278
rect 35870 23202 35922 23214
rect 37326 23266 37378 23278
rect 37326 23202 37378 23214
rect 41806 23266 41858 23278
rect 41806 23202 41858 23214
rect 20190 23154 20242 23166
rect 2482 23102 2494 23154
rect 2546 23102 2558 23154
rect 10770 23102 10782 23154
rect 10834 23102 10846 23154
rect 11666 23102 11678 23154
rect 11730 23102 11742 23154
rect 12674 23102 12686 23154
rect 12738 23102 12750 23154
rect 13794 23102 13806 23154
rect 13858 23102 13870 23154
rect 17490 23102 17502 23154
rect 17554 23102 17566 23154
rect 19394 23102 19406 23154
rect 19458 23102 19470 23154
rect 19842 23102 19854 23154
rect 19906 23102 19918 23154
rect 20190 23090 20242 23102
rect 20414 23154 20466 23166
rect 20414 23090 20466 23102
rect 20750 23154 20802 23166
rect 20750 23090 20802 23102
rect 23326 23154 23378 23166
rect 23326 23090 23378 23102
rect 23550 23154 23602 23166
rect 23550 23090 23602 23102
rect 24446 23154 24498 23166
rect 26014 23154 26066 23166
rect 25554 23102 25566 23154
rect 25618 23102 25630 23154
rect 24446 23090 24498 23102
rect 26014 23090 26066 23102
rect 26350 23154 26402 23166
rect 29486 23154 29538 23166
rect 28914 23102 28926 23154
rect 28978 23102 28990 23154
rect 26350 23090 26402 23102
rect 29486 23090 29538 23102
rect 34974 23154 35026 23166
rect 36654 23154 36706 23166
rect 35410 23102 35422 23154
rect 35474 23102 35486 23154
rect 34974 23090 35026 23102
rect 36654 23090 36706 23102
rect 36990 23154 37042 23166
rect 36990 23090 37042 23102
rect 39454 23154 39506 23166
rect 39666 23102 39678 23154
rect 39730 23102 39742 23154
rect 41122 23102 41134 23154
rect 41186 23102 41198 23154
rect 41570 23102 41582 23154
rect 41634 23102 41646 23154
rect 39454 23090 39506 23102
rect 5854 23042 5906 23054
rect 16046 23042 16098 23054
rect 5282 22990 5294 23042
rect 5346 22990 5358 23042
rect 14466 22990 14478 23042
rect 14530 22990 14542 23042
rect 5854 22978 5906 22990
rect 16046 22978 16098 22990
rect 17950 23042 18002 23054
rect 17950 22978 18002 22990
rect 23886 23042 23938 23054
rect 36542 23042 36594 23054
rect 29922 22990 29934 23042
rect 29986 22990 29998 23042
rect 23886 22978 23938 22990
rect 36542 22978 36594 22990
rect 36878 23042 36930 23054
rect 36878 22978 36930 22990
rect 40350 23042 40402 23054
rect 40350 22978 40402 22990
rect 14690 22878 14702 22930
rect 14754 22878 14766 22930
rect 22978 22878 22990 22930
rect 23042 22878 23054 22930
rect 41234 22878 41246 22930
rect 41298 22878 41310 22930
rect 1344 22762 44576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 44576 22762
rect 1344 22676 44576 22710
rect 19406 22594 19458 22606
rect 16146 22542 16158 22594
rect 16210 22542 16222 22594
rect 19406 22530 19458 22542
rect 40798 22594 40850 22606
rect 40798 22530 40850 22542
rect 41134 22594 41186 22606
rect 41134 22530 41186 22542
rect 19630 22482 19682 22494
rect 40014 22482 40066 22494
rect 15922 22430 15934 22482
rect 15986 22430 15998 22482
rect 26226 22430 26238 22482
rect 26290 22430 26302 22482
rect 19630 22418 19682 22430
rect 40014 22418 40066 22430
rect 17166 22370 17218 22382
rect 21534 22370 21586 22382
rect 40574 22370 40626 22382
rect 13458 22318 13470 22370
rect 13522 22318 13534 22370
rect 14354 22318 14366 22370
rect 14418 22318 14430 22370
rect 19058 22318 19070 22370
rect 19122 22318 19134 22370
rect 21746 22318 21758 22370
rect 21810 22318 21822 22370
rect 17166 22306 17218 22318
rect 21534 22306 21586 22318
rect 40574 22306 40626 22318
rect 17054 22258 17106 22270
rect 14466 22206 14478 22258
rect 14530 22206 14542 22258
rect 15698 22206 15710 22258
rect 15762 22206 15774 22258
rect 17054 22194 17106 22206
rect 41022 22258 41074 22270
rect 41022 22194 41074 22206
rect 13694 22146 13746 22158
rect 13794 22094 13806 22146
rect 13858 22094 13870 22146
rect 13694 22082 13746 22094
rect 1344 21978 44576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 44576 21978
rect 1344 21892 44576 21926
rect 15374 21810 15426 21822
rect 13570 21758 13582 21810
rect 13634 21758 13646 21810
rect 15374 21746 15426 21758
rect 24670 21810 24722 21822
rect 24670 21746 24722 21758
rect 25790 21810 25842 21822
rect 25790 21746 25842 21758
rect 42590 21810 42642 21822
rect 42590 21746 42642 21758
rect 18846 21698 18898 21710
rect 10322 21646 10334 21698
rect 10386 21646 10398 21698
rect 12898 21646 12910 21698
rect 12962 21646 12974 21698
rect 18846 21634 18898 21646
rect 19070 21698 19122 21710
rect 19070 21634 19122 21646
rect 26686 21698 26738 21710
rect 26686 21634 26738 21646
rect 28926 21698 28978 21710
rect 29586 21646 29598 21698
rect 29650 21646 29662 21698
rect 30034 21646 30046 21698
rect 30098 21646 30110 21698
rect 37090 21646 37102 21698
rect 37154 21646 37166 21698
rect 28926 21634 28978 21646
rect 7310 21586 7362 21598
rect 6850 21534 6862 21586
rect 6914 21534 6926 21586
rect 7310 21522 7362 21534
rect 7422 21586 7474 21598
rect 9986 21534 9998 21586
rect 10050 21534 10062 21586
rect 11330 21534 11342 21586
rect 11394 21534 11406 21586
rect 13346 21534 13358 21586
rect 13410 21534 13422 21586
rect 30146 21534 30158 21586
rect 30210 21534 30222 21586
rect 36418 21534 36430 21586
rect 36482 21534 36494 21586
rect 7422 21522 7474 21534
rect 18958 21474 19010 21486
rect 18958 21410 19010 21422
rect 25230 21474 25282 21486
rect 25230 21410 25282 21422
rect 26126 21474 26178 21486
rect 39790 21474 39842 21486
rect 39218 21422 39230 21474
rect 39282 21422 39294 21474
rect 26126 21410 26178 21422
rect 39790 21410 39842 21422
rect 42702 21474 42754 21486
rect 42702 21410 42754 21422
rect 1344 21194 44576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 44576 21194
rect 1344 21108 44576 21142
rect 29810 20974 29822 21026
rect 29874 20974 29886 21026
rect 16942 20914 16994 20926
rect 11330 20862 11342 20914
rect 11394 20862 11406 20914
rect 16146 20862 16158 20914
rect 16210 20862 16222 20914
rect 16942 20850 16994 20862
rect 26238 20914 26290 20926
rect 41458 20862 41470 20914
rect 41522 20862 41534 20914
rect 43586 20862 43598 20914
rect 43650 20862 43662 20914
rect 26238 20850 26290 20862
rect 17054 20802 17106 20814
rect 8418 20750 8430 20802
rect 8482 20750 8494 20802
rect 9426 20750 9438 20802
rect 9490 20750 9502 20802
rect 10546 20750 10558 20802
rect 10610 20750 10622 20802
rect 10882 20750 10894 20802
rect 10946 20750 10958 20802
rect 13794 20750 13806 20802
rect 13858 20750 13870 20802
rect 15138 20750 15150 20802
rect 15202 20750 15214 20802
rect 17054 20738 17106 20750
rect 25230 20802 25282 20814
rect 30158 20802 30210 20814
rect 25666 20750 25678 20802
rect 25730 20750 25742 20802
rect 25230 20738 25282 20750
rect 30158 20738 30210 20750
rect 30382 20802 30434 20814
rect 30382 20738 30434 20750
rect 30606 20802 30658 20814
rect 40674 20750 40686 20802
rect 40738 20750 40750 20802
rect 30606 20738 30658 20750
rect 9202 20638 9214 20690
rect 9266 20638 9278 20690
rect 11218 20638 11230 20690
rect 11282 20638 11294 20690
rect 14018 20638 14030 20690
rect 14082 20638 14094 20690
rect 15026 20638 15038 20690
rect 15090 20638 15102 20690
rect 17266 20638 17278 20690
rect 17330 20638 17342 20690
rect 18050 20638 18062 20690
rect 18114 20638 18126 20690
rect 8430 20578 8482 20590
rect 40350 20578 40402 20590
rect 9314 20526 9326 20578
rect 9378 20526 9390 20578
rect 10098 20526 10110 20578
rect 10162 20526 10174 20578
rect 8430 20514 8482 20526
rect 40350 20514 40402 20526
rect 1344 20410 44576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 44576 20410
rect 1344 20324 44576 20358
rect 8990 20242 9042 20254
rect 8990 20178 9042 20190
rect 10222 20242 10274 20254
rect 15474 20190 15486 20242
rect 15538 20190 15550 20242
rect 10222 20178 10274 20190
rect 8542 20130 8594 20142
rect 8542 20066 8594 20078
rect 9998 20130 10050 20142
rect 9998 20066 10050 20078
rect 10446 20130 10498 20142
rect 10446 20066 10498 20078
rect 14814 20130 14866 20142
rect 16034 20078 16046 20130
rect 16098 20078 16110 20130
rect 14814 20066 14866 20078
rect 8430 20018 8482 20030
rect 8430 19954 8482 19966
rect 8878 20018 8930 20030
rect 8878 19954 8930 19966
rect 10782 20018 10834 20030
rect 19742 20018 19794 20030
rect 14578 19966 14590 20018
rect 14642 19966 14654 20018
rect 15810 19966 15822 20018
rect 15874 19966 15886 20018
rect 10782 19954 10834 19966
rect 19742 19954 19794 19966
rect 19966 20018 20018 20030
rect 19966 19954 20018 19966
rect 20414 20018 20466 20030
rect 29474 19966 29486 20018
rect 29538 19966 29550 20018
rect 20414 19954 20466 19966
rect 4958 19906 5010 19918
rect 4958 19842 5010 19854
rect 10334 19906 10386 19918
rect 10334 19842 10386 19854
rect 10894 19906 10946 19918
rect 10894 19842 10946 19854
rect 19854 19906 19906 19918
rect 33182 19906 33234 19918
rect 30146 19854 30158 19906
rect 30210 19854 30222 19906
rect 32274 19854 32286 19906
rect 32338 19854 32350 19906
rect 19854 19842 19906 19854
rect 33182 19842 33234 19854
rect 1344 19626 44576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 44576 19626
rect 1344 19540 44576 19574
rect 9886 19458 9938 19470
rect 9886 19394 9938 19406
rect 15150 19458 15202 19470
rect 15150 19394 15202 19406
rect 30158 19458 30210 19470
rect 30158 19394 30210 19406
rect 30494 19458 30546 19470
rect 31266 19406 31278 19458
rect 31330 19406 31342 19458
rect 30494 19394 30546 19406
rect 28030 19346 28082 19358
rect 4722 19294 4734 19346
rect 4786 19294 4798 19346
rect 5730 19294 5742 19346
rect 5794 19294 5806 19346
rect 17826 19294 17838 19346
rect 17890 19294 17902 19346
rect 27570 19294 27582 19346
rect 27634 19294 27646 19346
rect 33506 19294 33518 19346
rect 33570 19294 33582 19346
rect 28030 19282 28082 19294
rect 30270 19234 30322 19246
rect 1810 19182 1822 19234
rect 1874 19182 1886 19234
rect 6066 19182 6078 19234
rect 6130 19182 6142 19234
rect 20626 19182 20638 19234
rect 20690 19182 20702 19234
rect 24098 19182 24110 19234
rect 24162 19182 24174 19234
rect 24770 19182 24782 19234
rect 24834 19182 24846 19234
rect 30270 19170 30322 19182
rect 30606 19234 30658 19246
rect 31950 19234 32002 19246
rect 31714 19182 31726 19234
rect 31778 19182 31790 19234
rect 36418 19182 36430 19234
rect 36482 19182 36494 19234
rect 30606 19170 30658 19182
rect 31950 19170 32002 19182
rect 9774 19122 9826 19134
rect 2594 19070 2606 19122
rect 2658 19070 2670 19122
rect 9774 19058 9826 19070
rect 15038 19122 15090 19134
rect 24334 19122 24386 19134
rect 19954 19070 19966 19122
rect 20018 19070 20030 19122
rect 25442 19070 25454 19122
rect 25506 19070 25518 19122
rect 35634 19070 35646 19122
rect 35698 19070 35710 19122
rect 15038 19058 15090 19070
rect 24334 19058 24386 19070
rect 21422 19010 21474 19022
rect 21422 18946 21474 18958
rect 29822 19010 29874 19022
rect 29822 18946 29874 18958
rect 37102 19010 37154 19022
rect 37102 18946 37154 18958
rect 1344 18842 44576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 44576 18842
rect 1344 18756 44576 18790
rect 14254 18674 14306 18686
rect 10546 18622 10558 18674
rect 10610 18622 10622 18674
rect 14254 18610 14306 18622
rect 14702 18674 14754 18686
rect 20190 18674 20242 18686
rect 19506 18622 19518 18674
rect 19570 18622 19582 18674
rect 24546 18622 24558 18674
rect 24610 18622 24622 18674
rect 31826 18622 31838 18674
rect 31890 18622 31902 18674
rect 14702 18610 14754 18622
rect 20190 18610 20242 18622
rect 4062 18562 4114 18574
rect 14478 18562 14530 18574
rect 10098 18510 10110 18562
rect 10162 18510 10174 18562
rect 10658 18510 10670 18562
rect 10722 18510 10734 18562
rect 4062 18498 4114 18510
rect 14478 18498 14530 18510
rect 14814 18562 14866 18574
rect 14814 18498 14866 18510
rect 19070 18562 19122 18574
rect 19070 18498 19122 18510
rect 23214 18562 23266 18574
rect 23214 18498 23266 18510
rect 23438 18562 23490 18574
rect 23438 18498 23490 18510
rect 34526 18562 34578 18574
rect 34526 18498 34578 18510
rect 11006 18450 11058 18462
rect 5170 18398 5182 18450
rect 5234 18398 5246 18450
rect 11006 18386 11058 18398
rect 13806 18450 13858 18462
rect 13806 18386 13858 18398
rect 14366 18450 14418 18462
rect 14366 18386 14418 18398
rect 15038 18450 15090 18462
rect 20750 18450 20802 18462
rect 23550 18450 23602 18462
rect 15474 18398 15486 18450
rect 15538 18398 15550 18450
rect 15698 18398 15710 18450
rect 15762 18398 15774 18450
rect 19282 18398 19294 18450
rect 19346 18398 19358 18450
rect 19618 18398 19630 18450
rect 19682 18398 19694 18450
rect 22978 18398 22990 18450
rect 23042 18398 23054 18450
rect 15038 18386 15090 18398
rect 20750 18386 20802 18398
rect 23550 18386 23602 18398
rect 23886 18450 23938 18462
rect 23886 18386 23938 18398
rect 23998 18450 24050 18462
rect 23998 18386 24050 18398
rect 24110 18450 24162 18462
rect 24110 18386 24162 18398
rect 32174 18450 32226 18462
rect 32174 18386 32226 18398
rect 33966 18450 34018 18462
rect 33966 18386 34018 18398
rect 34302 18450 34354 18462
rect 34302 18386 34354 18398
rect 5630 18338 5682 18350
rect 3938 18286 3950 18338
rect 4002 18286 4014 18338
rect 4834 18286 4846 18338
rect 4898 18286 4910 18338
rect 5630 18274 5682 18286
rect 16158 18338 16210 18350
rect 16158 18274 16210 18286
rect 22654 18338 22706 18350
rect 22654 18274 22706 18286
rect 32398 18338 32450 18350
rect 34626 18286 34638 18338
rect 34690 18286 34702 18338
rect 32398 18274 32450 18286
rect 4286 18226 4338 18238
rect 4286 18162 4338 18174
rect 15262 18226 15314 18238
rect 15262 18162 15314 18174
rect 19518 18226 19570 18238
rect 19518 18162 19570 18174
rect 1344 18058 44576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 44576 18058
rect 1344 17972 44576 18006
rect 4510 17778 4562 17790
rect 4510 17714 4562 17726
rect 5966 17778 6018 17790
rect 5966 17714 6018 17726
rect 12014 17778 12066 17790
rect 22878 17778 22930 17790
rect 14690 17726 14702 17778
rect 14754 17726 14766 17778
rect 16818 17726 16830 17778
rect 16882 17726 16894 17778
rect 12014 17714 12066 17726
rect 22878 17714 22930 17726
rect 23326 17778 23378 17790
rect 23326 17714 23378 17726
rect 24446 17778 24498 17790
rect 24446 17714 24498 17726
rect 6078 17666 6130 17678
rect 5618 17614 5630 17666
rect 5682 17614 5694 17666
rect 6078 17602 6130 17614
rect 9886 17666 9938 17678
rect 9886 17602 9938 17614
rect 10110 17666 10162 17678
rect 10110 17602 10162 17614
rect 10222 17666 10274 17678
rect 10222 17602 10274 17614
rect 10446 17666 10498 17678
rect 10446 17602 10498 17614
rect 11230 17666 11282 17678
rect 11230 17602 11282 17614
rect 11454 17666 11506 17678
rect 23438 17666 23490 17678
rect 14018 17614 14030 17666
rect 14082 17614 14094 17666
rect 11454 17602 11506 17614
rect 23438 17602 23490 17614
rect 23886 17666 23938 17678
rect 23886 17602 23938 17614
rect 24334 17666 24386 17678
rect 35758 17666 35810 17678
rect 32946 17614 32958 17666
rect 33010 17614 33022 17666
rect 24334 17602 24386 17614
rect 35758 17602 35810 17614
rect 11006 17554 11058 17566
rect 11006 17490 11058 17502
rect 23214 17554 23266 17566
rect 35198 17554 35250 17566
rect 32386 17502 32398 17554
rect 32450 17502 32462 17554
rect 32834 17502 32846 17554
rect 32898 17502 32910 17554
rect 23214 17490 23266 17502
rect 35198 17490 35250 17502
rect 35310 17554 35362 17566
rect 35310 17490 35362 17502
rect 35870 17554 35922 17566
rect 35870 17490 35922 17502
rect 36990 17554 37042 17566
rect 36990 17490 37042 17502
rect 5854 17442 5906 17454
rect 5854 17378 5906 17390
rect 6190 17442 6242 17454
rect 11118 17442 11170 17454
rect 9426 17390 9438 17442
rect 9490 17390 9502 17442
rect 6190 17378 6242 17390
rect 11118 17378 11170 17390
rect 17278 17442 17330 17454
rect 35534 17442 35586 17454
rect 32274 17390 32286 17442
rect 32338 17390 32350 17442
rect 17278 17378 17330 17390
rect 35534 17378 35586 17390
rect 37326 17442 37378 17454
rect 37326 17378 37378 17390
rect 1344 17274 44576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 44576 17274
rect 1344 17188 44576 17222
rect 17502 17106 17554 17118
rect 17502 17042 17554 17054
rect 30494 17106 30546 17118
rect 30494 17042 30546 17054
rect 30942 17106 30994 17118
rect 30942 17042 30994 17054
rect 9662 16994 9714 17006
rect 31054 16994 31106 17006
rect 6738 16942 6750 16994
rect 6802 16942 6814 16994
rect 10210 16942 10222 16994
rect 10274 16942 10286 16994
rect 9662 16930 9714 16942
rect 31054 16930 31106 16942
rect 15710 16882 15762 16894
rect 6066 16830 6078 16882
rect 6130 16830 6142 16882
rect 15250 16830 15262 16882
rect 15314 16830 15326 16882
rect 15710 16818 15762 16830
rect 17614 16882 17666 16894
rect 17614 16818 17666 16830
rect 20190 16882 20242 16894
rect 20190 16818 20242 16830
rect 20750 16882 20802 16894
rect 32510 16882 32562 16894
rect 31602 16830 31614 16882
rect 31666 16830 31678 16882
rect 33058 16830 33070 16882
rect 33122 16830 33134 16882
rect 20750 16818 20802 16830
rect 32510 16818 32562 16830
rect 31950 16770 32002 16782
rect 8866 16718 8878 16770
rect 8930 16718 8942 16770
rect 37090 16718 37102 16770
rect 37154 16718 37166 16770
rect 31950 16706 32002 16718
rect 17502 16658 17554 16670
rect 17502 16594 17554 16606
rect 30942 16658 30994 16670
rect 30942 16594 30994 16606
rect 31614 16658 31666 16670
rect 31614 16594 31666 16606
rect 1344 16490 44576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 44576 16490
rect 1344 16404 44576 16438
rect 23438 16322 23490 16334
rect 23438 16258 23490 16270
rect 31054 16322 31106 16334
rect 31054 16258 31106 16270
rect 34862 16322 34914 16334
rect 36418 16270 36430 16322
rect 36482 16270 36494 16322
rect 34862 16258 34914 16270
rect 10222 16210 10274 16222
rect 35870 16210 35922 16222
rect 10994 16158 11006 16210
rect 11058 16158 11070 16210
rect 31266 16158 31278 16210
rect 31330 16158 31342 16210
rect 37426 16158 37438 16210
rect 37490 16158 37502 16210
rect 39554 16158 39566 16210
rect 39618 16158 39630 16210
rect 10222 16146 10274 16158
rect 35870 16146 35922 16158
rect 9662 16098 9714 16110
rect 11230 16098 11282 16110
rect 10546 16046 10558 16098
rect 10610 16046 10622 16098
rect 10770 16046 10782 16098
rect 10834 16046 10846 16098
rect 9662 16034 9714 16046
rect 11230 16034 11282 16046
rect 11566 16098 11618 16110
rect 11566 16034 11618 16046
rect 12910 16098 12962 16110
rect 12910 16034 12962 16046
rect 13806 16098 13858 16110
rect 23326 16098 23378 16110
rect 34414 16098 34466 16110
rect 15698 16046 15710 16098
rect 15762 16046 15774 16098
rect 31378 16046 31390 16098
rect 31442 16046 31454 16098
rect 13806 16034 13858 16046
rect 23326 16034 23378 16046
rect 34414 16034 34466 16046
rect 36094 16098 36146 16110
rect 40338 16046 40350 16098
rect 40402 16046 40414 16098
rect 36094 16034 36146 16046
rect 11006 15986 11058 15998
rect 11006 15922 11058 15934
rect 11454 15986 11506 15998
rect 33854 15986 33906 15998
rect 12562 15934 12574 15986
rect 12626 15934 12638 15986
rect 13458 15934 13470 15986
rect 13522 15934 13534 15986
rect 18386 15934 18398 15986
rect 18450 15934 18462 15986
rect 11454 15922 11506 15934
rect 33854 15922 33906 15934
rect 34302 15986 34354 15998
rect 34302 15922 34354 15934
rect 34526 15986 34578 15998
rect 34526 15922 34578 15934
rect 34974 15986 35026 15998
rect 34974 15922 35026 15934
rect 35086 15986 35138 15998
rect 35086 15922 35138 15934
rect 19966 15874 20018 15886
rect 19966 15810 20018 15822
rect 22990 15874 23042 15886
rect 22990 15810 23042 15822
rect 23438 15874 23490 15886
rect 23438 15810 23490 15822
rect 37102 15874 37154 15886
rect 37102 15810 37154 15822
rect 1344 15706 44576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 44576 15706
rect 1344 15620 44576 15654
rect 33182 15538 33234 15550
rect 19842 15486 19854 15538
rect 19906 15486 19918 15538
rect 25330 15486 25342 15538
rect 25394 15486 25406 15538
rect 35970 15486 35982 15538
rect 36034 15486 36046 15538
rect 33182 15474 33234 15486
rect 23214 15426 23266 15438
rect 23214 15362 23266 15374
rect 23326 15426 23378 15438
rect 23326 15362 23378 15374
rect 23550 15426 23602 15438
rect 25790 15426 25842 15438
rect 23986 15374 23998 15426
rect 24050 15374 24062 15426
rect 23550 15362 23602 15374
rect 25790 15362 25842 15374
rect 27806 15426 27858 15438
rect 35422 15426 35474 15438
rect 31714 15374 31726 15426
rect 31778 15374 31790 15426
rect 27806 15362 27858 15374
rect 35422 15362 35474 15374
rect 36878 15426 36930 15438
rect 36878 15362 36930 15374
rect 23662 15314 23714 15326
rect 19618 15262 19630 15314
rect 19682 15262 19694 15314
rect 20738 15262 20750 15314
rect 20802 15262 20814 15314
rect 23662 15250 23714 15262
rect 24222 15314 24274 15326
rect 24222 15250 24274 15262
rect 24670 15314 24722 15326
rect 25218 15262 25230 15314
rect 25282 15262 25294 15314
rect 29026 15262 29038 15314
rect 29090 15262 29102 15314
rect 32498 15262 32510 15314
rect 32562 15262 32574 15314
rect 34178 15262 34190 15314
rect 34242 15262 34254 15314
rect 37986 15262 37998 15314
rect 38050 15262 38062 15314
rect 24670 15250 24722 15262
rect 24446 15202 24498 15214
rect 20402 15150 20414 15202
rect 20466 15150 20478 15202
rect 24446 15138 24498 15150
rect 24558 15202 24610 15214
rect 29586 15150 29598 15202
rect 29650 15150 29662 15202
rect 24558 15138 24610 15150
rect 1344 14922 44576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 44576 14922
rect 1344 14836 44576 14870
rect 25454 14754 25506 14766
rect 23314 14702 23326 14754
rect 23378 14702 23390 14754
rect 25454 14690 25506 14702
rect 15150 14642 15202 14654
rect 5730 14590 5742 14642
rect 5794 14590 5806 14642
rect 15150 14578 15202 14590
rect 20078 14642 20130 14654
rect 20078 14578 20130 14590
rect 25006 14642 25058 14654
rect 25006 14578 25058 14590
rect 25566 14642 25618 14654
rect 25566 14578 25618 14590
rect 28702 14642 28754 14654
rect 31938 14590 31950 14642
rect 32002 14590 32014 14642
rect 28702 14578 28754 14590
rect 22990 14530 23042 14542
rect 1922 14478 1934 14530
rect 1986 14478 1998 14530
rect 23650 14478 23662 14530
rect 23714 14478 23726 14530
rect 24434 14478 24446 14530
rect 24498 14478 24510 14530
rect 29138 14478 29150 14530
rect 29202 14478 29214 14530
rect 22990 14466 23042 14478
rect 14254 14418 14306 14430
rect 2594 14366 2606 14418
rect 2658 14366 2670 14418
rect 14254 14354 14306 14366
rect 14366 14418 14418 14430
rect 24222 14418 24274 14430
rect 15474 14366 15486 14418
rect 15538 14366 15550 14418
rect 14366 14354 14418 14366
rect 24222 14354 24274 14366
rect 6190 14306 6242 14318
rect 4834 14254 4846 14306
rect 4898 14254 4910 14306
rect 6190 14242 6242 14254
rect 14590 14306 14642 14318
rect 14590 14242 14642 14254
rect 1344 14138 44576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 44576 14138
rect 1344 14052 44576 14086
rect 9998 13970 10050 13982
rect 12014 13970 12066 13982
rect 11666 13918 11678 13970
rect 11730 13918 11742 13970
rect 9998 13906 10050 13918
rect 12014 13906 12066 13918
rect 12462 13970 12514 13982
rect 12462 13906 12514 13918
rect 14254 13970 14306 13982
rect 14254 13906 14306 13918
rect 16046 13970 16098 13982
rect 16046 13906 16098 13918
rect 30046 13970 30098 13982
rect 30046 13906 30098 13918
rect 35422 13970 35474 13982
rect 35422 13906 35474 13918
rect 35646 13970 35698 13982
rect 35646 13906 35698 13918
rect 15598 13858 15650 13870
rect 14914 13806 14926 13858
rect 14978 13806 14990 13858
rect 27234 13806 27246 13858
rect 27298 13806 27310 13858
rect 15598 13794 15650 13806
rect 9774 13746 9826 13758
rect 13694 13746 13746 13758
rect 9538 13694 9550 13746
rect 9602 13694 9614 13746
rect 10210 13694 10222 13746
rect 10274 13694 10286 13746
rect 9774 13682 9826 13694
rect 13694 13682 13746 13694
rect 14142 13746 14194 13758
rect 14142 13682 14194 13694
rect 14366 13746 14418 13758
rect 14366 13682 14418 13694
rect 14590 13746 14642 13758
rect 14590 13682 14642 13694
rect 15374 13746 15426 13758
rect 34974 13746 35026 13758
rect 26562 13694 26574 13746
rect 26626 13694 26638 13746
rect 15374 13682 15426 13694
rect 34974 13682 35026 13694
rect 36318 13746 36370 13758
rect 36318 13682 36370 13694
rect 36542 13746 36594 13758
rect 36542 13682 36594 13694
rect 5182 13634 5234 13646
rect 5182 13570 5234 13582
rect 9886 13634 9938 13646
rect 9886 13570 9938 13582
rect 15486 13634 15538 13646
rect 15486 13570 15538 13582
rect 29374 13634 29426 13646
rect 29374 13570 29426 13582
rect 34750 13634 34802 13646
rect 34750 13570 34802 13582
rect 35534 13634 35586 13646
rect 35534 13570 35586 13582
rect 15150 13522 15202 13534
rect 35970 13470 35982 13522
rect 36034 13470 36046 13522
rect 15150 13458 15202 13470
rect 1344 13354 44576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 44576 13354
rect 1344 13268 44576 13302
rect 24110 13186 24162 13198
rect 24110 13122 24162 13134
rect 35870 13186 35922 13198
rect 35870 13122 35922 13134
rect 5742 13074 5794 13086
rect 12910 13074 12962 13086
rect 21870 13074 21922 13086
rect 10210 13022 10222 13074
rect 10274 13022 10286 13074
rect 15026 13022 15038 13074
rect 15090 13022 15102 13074
rect 15698 13022 15710 13074
rect 15762 13022 15774 13074
rect 17826 13022 17838 13074
rect 17890 13022 17902 13074
rect 36082 13022 36094 13074
rect 36146 13022 36158 13074
rect 36978 13022 36990 13074
rect 37042 13022 37054 13074
rect 39106 13022 39118 13074
rect 39170 13022 39182 13074
rect 5742 13010 5794 13022
rect 12910 13010 12962 13022
rect 21870 13010 21922 13022
rect 6078 12962 6130 12974
rect 14926 12962 14978 12974
rect 23438 12962 23490 12974
rect 6402 12910 6414 12962
rect 6466 12910 6478 12962
rect 6962 12910 6974 12962
rect 7026 12910 7038 12962
rect 8418 12910 8430 12962
rect 8482 12910 8494 12962
rect 9874 12910 9886 12962
rect 9938 12910 9950 12962
rect 12226 12910 12238 12962
rect 12290 12910 12302 12962
rect 18610 12910 18622 12962
rect 18674 12910 18686 12962
rect 25666 12910 25678 12962
rect 25730 12910 25742 12962
rect 39778 12910 39790 12962
rect 39842 12910 39854 12962
rect 6078 12898 6130 12910
rect 14926 12898 14978 12910
rect 23438 12898 23490 12910
rect 4958 12850 5010 12862
rect 4958 12786 5010 12798
rect 5070 12850 5122 12862
rect 5070 12786 5122 12798
rect 5630 12850 5682 12862
rect 7422 12850 7474 12862
rect 14590 12850 14642 12862
rect 5842 12798 5854 12850
rect 5906 12798 5918 12850
rect 8754 12798 8766 12850
rect 8818 12798 8830 12850
rect 9762 12798 9774 12850
rect 9826 12798 9838 12850
rect 12450 12798 12462 12850
rect 12514 12798 12526 12850
rect 5630 12786 5682 12798
rect 7422 12786 7474 12798
rect 14590 12786 14642 12798
rect 23998 12850 24050 12862
rect 23998 12786 24050 12798
rect 36094 12850 36146 12862
rect 36094 12786 36146 12798
rect 7198 12738 7250 12750
rect 7198 12674 7250 12686
rect 7534 12738 7586 12750
rect 7534 12674 7586 12686
rect 19070 12738 19122 12750
rect 19070 12674 19122 12686
rect 23774 12738 23826 12750
rect 23774 12674 23826 12686
rect 24446 12738 24498 12750
rect 25442 12686 25454 12738
rect 25506 12686 25518 12738
rect 24446 12674 24498 12686
rect 1344 12570 44576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 44576 12570
rect 1344 12484 44576 12518
rect 5294 12402 5346 12414
rect 5294 12338 5346 12350
rect 6638 12402 6690 12414
rect 6638 12338 6690 12350
rect 8542 12402 8594 12414
rect 8542 12338 8594 12350
rect 8654 12402 8706 12414
rect 8654 12338 8706 12350
rect 8766 12402 8818 12414
rect 11454 12402 11506 12414
rect 22206 12402 22258 12414
rect 9762 12350 9774 12402
rect 9826 12350 9838 12402
rect 20738 12350 20750 12402
rect 20802 12350 20814 12402
rect 8766 12338 8818 12350
rect 11454 12338 11506 12350
rect 22206 12338 22258 12350
rect 23438 12402 23490 12414
rect 23438 12338 23490 12350
rect 24558 12402 24610 12414
rect 24558 12338 24610 12350
rect 5518 12290 5570 12302
rect 5518 12226 5570 12238
rect 8318 12290 8370 12302
rect 8318 12226 8370 12238
rect 9550 12290 9602 12302
rect 9550 12226 9602 12238
rect 11006 12290 11058 12302
rect 11006 12226 11058 12238
rect 21086 12290 21138 12302
rect 21086 12226 21138 12238
rect 22654 12290 22706 12302
rect 22654 12226 22706 12238
rect 23662 12290 23714 12302
rect 23662 12226 23714 12238
rect 24110 12290 24162 12302
rect 24110 12226 24162 12238
rect 24670 12290 24722 12302
rect 24670 12226 24722 12238
rect 5630 12178 5682 12190
rect 9998 12178 10050 12190
rect 22094 12178 22146 12190
rect 8978 12126 8990 12178
rect 9042 12126 9054 12178
rect 9762 12126 9774 12178
rect 9826 12126 9838 12178
rect 10098 12126 10110 12178
rect 10162 12126 10174 12178
rect 10658 12126 10670 12178
rect 10722 12126 10734 12178
rect 20514 12126 20526 12178
rect 20578 12126 20590 12178
rect 5630 12114 5682 12126
rect 9998 12114 10050 12126
rect 22094 12114 22146 12126
rect 22430 12178 22482 12190
rect 22430 12114 22482 12126
rect 23102 12178 23154 12190
rect 23102 12114 23154 12126
rect 23214 12178 23266 12190
rect 23214 12114 23266 12126
rect 23998 12178 24050 12190
rect 23998 12114 24050 12126
rect 24334 12178 24386 12190
rect 24334 12114 24386 12126
rect 21646 12066 21698 12078
rect 21646 12002 21698 12014
rect 22318 12066 22370 12078
rect 22318 12002 22370 12014
rect 23774 12066 23826 12078
rect 23774 12002 23826 12014
rect 36654 12066 36706 12078
rect 36654 12002 36706 12014
rect 21310 11954 21362 11966
rect 21310 11890 21362 11902
rect 1344 11786 44576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 44576 11786
rect 1344 11700 44576 11734
rect 14926 11506 14978 11518
rect 13906 11454 13918 11506
rect 13970 11454 13982 11506
rect 14926 11442 14978 11454
rect 22206 11506 22258 11518
rect 34526 11506 34578 11518
rect 25218 11454 25230 11506
rect 25282 11454 25294 11506
rect 22206 11442 22258 11454
rect 34526 11442 34578 11454
rect 4398 11394 4450 11406
rect 5742 11394 5794 11406
rect 4834 11342 4846 11394
rect 4898 11342 4910 11394
rect 4398 11330 4450 11342
rect 5742 11330 5794 11342
rect 6078 11394 6130 11406
rect 6078 11330 6130 11342
rect 6638 11394 6690 11406
rect 6638 11330 6690 11342
rect 6750 11394 6802 11406
rect 6750 11330 6802 11342
rect 6862 11394 6914 11406
rect 6862 11330 6914 11342
rect 14030 11394 14082 11406
rect 14030 11330 14082 11342
rect 14254 11394 14306 11406
rect 14254 11330 14306 11342
rect 14366 11394 14418 11406
rect 14366 11330 14418 11342
rect 21758 11394 21810 11406
rect 21758 11330 21810 11342
rect 21982 11394 22034 11406
rect 21982 11330 22034 11342
rect 22430 11394 22482 11406
rect 22430 11330 22482 11342
rect 22654 11394 22706 11406
rect 23998 11394 24050 11406
rect 23650 11342 23662 11394
rect 23714 11342 23726 11394
rect 22654 11330 22706 11342
rect 23998 11330 24050 11342
rect 24334 11394 24386 11406
rect 24334 11330 24386 11342
rect 24670 11394 24722 11406
rect 34750 11394 34802 11406
rect 28130 11342 28142 11394
rect 28194 11342 28206 11394
rect 24670 11330 24722 11342
rect 34750 11330 34802 11342
rect 35422 11394 35474 11406
rect 35422 11330 35474 11342
rect 4174 11282 4226 11294
rect 5966 11282 6018 11294
rect 5058 11230 5070 11282
rect 5122 11230 5134 11282
rect 4174 11218 4226 11230
rect 5966 11218 6018 11230
rect 13918 11282 13970 11294
rect 13918 11218 13970 11230
rect 23438 11282 23490 11294
rect 23438 11218 23490 11230
rect 24222 11282 24274 11294
rect 27346 11230 27358 11282
rect 27410 11230 27422 11282
rect 24222 11218 24274 11230
rect 4286 11170 4338 11182
rect 4286 11106 4338 11118
rect 5854 11170 5906 11182
rect 5854 11106 5906 11118
rect 6190 11170 6242 11182
rect 6190 11106 6242 11118
rect 7086 11170 7138 11182
rect 7086 11106 7138 11118
rect 7646 11170 7698 11182
rect 7646 11106 7698 11118
rect 28590 11170 28642 11182
rect 28590 11106 28642 11118
rect 35198 11170 35250 11182
rect 35198 11106 35250 11118
rect 35310 11170 35362 11182
rect 35310 11106 35362 11118
rect 1344 11002 44576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 44576 11002
rect 1344 10916 44576 10950
rect 11678 10834 11730 10846
rect 11678 10770 11730 10782
rect 12014 10834 12066 10846
rect 12014 10770 12066 10782
rect 14366 10834 14418 10846
rect 14366 10770 14418 10782
rect 15262 10834 15314 10846
rect 15262 10770 15314 10782
rect 25342 10834 25394 10846
rect 25342 10770 25394 10782
rect 31726 10834 31778 10846
rect 31726 10770 31778 10782
rect 35422 10722 35474 10734
rect 2594 10670 2606 10722
rect 2658 10670 2670 10722
rect 13794 10670 13806 10722
rect 13858 10670 13870 10722
rect 35422 10658 35474 10670
rect 35646 10722 35698 10734
rect 35646 10658 35698 10670
rect 11790 10610 11842 10622
rect 1922 10558 1934 10610
rect 1986 10558 1998 10610
rect 11790 10546 11842 10558
rect 12126 10610 12178 10622
rect 13582 10610 13634 10622
rect 13234 10558 13246 10610
rect 13298 10558 13310 10610
rect 12126 10546 12178 10558
rect 13582 10546 13634 10558
rect 14030 10610 14082 10622
rect 14926 10610 14978 10622
rect 34862 10610 34914 10622
rect 14578 10558 14590 10610
rect 14642 10558 14654 10610
rect 28466 10558 28478 10610
rect 28530 10558 28542 10610
rect 14030 10546 14082 10558
rect 14926 10546 14978 10558
rect 34862 10546 34914 10558
rect 35086 10610 35138 10622
rect 35086 10546 35138 10558
rect 5182 10498 5234 10510
rect 4722 10446 4734 10498
rect 4786 10446 4798 10498
rect 5182 10434 5234 10446
rect 11902 10498 11954 10510
rect 11902 10434 11954 10446
rect 13918 10498 13970 10510
rect 18286 10498 18338 10510
rect 14466 10446 14478 10498
rect 14530 10446 14542 10498
rect 13918 10434 13970 10446
rect 18286 10434 18338 10446
rect 19742 10498 19794 10510
rect 35534 10498 35586 10510
rect 29138 10446 29150 10498
rect 29202 10446 29214 10498
rect 31266 10446 31278 10498
rect 31330 10446 31342 10498
rect 19742 10434 19794 10446
rect 35534 10434 35586 10446
rect 34514 10334 34526 10386
rect 34578 10334 34590 10386
rect 1344 10218 44576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 44576 10218
rect 1344 10132 44576 10166
rect 17278 10050 17330 10062
rect 17278 9986 17330 9998
rect 20414 10050 20466 10062
rect 20414 9986 20466 9998
rect 29598 10050 29650 10062
rect 29598 9986 29650 9998
rect 29710 10050 29762 10062
rect 31378 9998 31390 10050
rect 31442 9998 31454 10050
rect 29710 9986 29762 9998
rect 12910 9938 12962 9950
rect 11218 9886 11230 9938
rect 11282 9886 11294 9938
rect 12910 9874 12962 9886
rect 15038 9938 15090 9950
rect 18722 9886 18734 9938
rect 18786 9886 18798 9938
rect 15038 9874 15090 9886
rect 12238 9826 12290 9838
rect 12238 9762 12290 9774
rect 13806 9826 13858 9838
rect 14926 9826 14978 9838
rect 14130 9774 14142 9826
rect 14194 9774 14206 9826
rect 13806 9762 13858 9774
rect 14926 9762 14978 9774
rect 17502 9826 17554 9838
rect 17502 9762 17554 9774
rect 18286 9826 18338 9838
rect 29374 9826 29426 9838
rect 19170 9774 19182 9826
rect 19234 9774 19246 9826
rect 19618 9774 19630 9826
rect 19682 9774 19694 9826
rect 18286 9762 18338 9774
rect 29374 9762 29426 9774
rect 29934 9826 29986 9838
rect 30606 9826 30658 9838
rect 30146 9774 30158 9826
rect 30210 9774 30222 9826
rect 29934 9762 29986 9774
rect 30606 9762 30658 9774
rect 31054 9826 31106 9838
rect 31054 9762 31106 9774
rect 31838 9826 31890 9838
rect 31838 9762 31890 9774
rect 32062 9826 32114 9838
rect 33954 9774 33966 9826
rect 34018 9774 34030 9826
rect 32062 9762 32114 9774
rect 11342 9714 11394 9726
rect 11342 9650 11394 9662
rect 11566 9714 11618 9726
rect 11566 9650 11618 9662
rect 12014 9714 12066 9726
rect 12014 9650 12066 9662
rect 12350 9714 12402 9726
rect 12350 9650 12402 9662
rect 14590 9714 14642 9726
rect 30494 9714 30546 9726
rect 17826 9662 17838 9714
rect 17890 9662 17902 9714
rect 18162 9662 18174 9714
rect 18226 9662 18238 9714
rect 18834 9662 18846 9714
rect 18898 9662 18910 9714
rect 14590 9650 14642 9662
rect 30494 9650 30546 9662
rect 30830 9714 30882 9726
rect 30830 9650 30882 9662
rect 31950 9714 32002 9726
rect 33730 9662 33742 9714
rect 33794 9662 33806 9714
rect 31950 9650 32002 9662
rect 12462 9602 12514 9614
rect 12462 9538 12514 9550
rect 20190 9602 20242 9614
rect 20190 9538 20242 9550
rect 20302 9602 20354 9614
rect 20302 9538 20354 9550
rect 1344 9434 44576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 44576 9434
rect 1344 9348 44576 9382
rect 12462 9266 12514 9278
rect 12462 9202 12514 9214
rect 12686 9266 12738 9278
rect 12686 9202 12738 9214
rect 18622 9266 18674 9278
rect 18622 9202 18674 9214
rect 18846 9266 18898 9278
rect 18846 9202 18898 9214
rect 19854 9266 19906 9278
rect 19854 9202 19906 9214
rect 31390 9266 31442 9278
rect 31390 9202 31442 9214
rect 12798 9154 12850 9166
rect 12798 9090 12850 9102
rect 20078 9154 20130 9166
rect 20078 9090 20130 9102
rect 32062 9154 32114 9166
rect 32062 9090 32114 9102
rect 33294 9154 33346 9166
rect 35522 9102 35534 9154
rect 35586 9102 35598 9154
rect 33294 9090 33346 9102
rect 17614 9042 17666 9054
rect 17614 8978 17666 8990
rect 17838 9042 17890 9054
rect 17838 8978 17890 8990
rect 18062 9042 18114 9054
rect 18062 8978 18114 8990
rect 18398 9042 18450 9054
rect 18398 8978 18450 8990
rect 18510 9042 18562 9054
rect 18510 8978 18562 8990
rect 19630 9042 19682 9054
rect 19630 8978 19682 8990
rect 31614 9042 31666 9054
rect 31614 8978 31666 8990
rect 32286 9042 32338 9054
rect 32286 8978 32338 8990
rect 33070 9042 33122 9054
rect 33070 8978 33122 8990
rect 33742 9042 33794 9054
rect 34850 8990 34862 9042
rect 34914 8990 34926 9042
rect 33742 8978 33794 8990
rect 17950 8930 18002 8942
rect 17950 8866 18002 8878
rect 19742 8930 19794 8942
rect 19742 8866 19794 8878
rect 32174 8930 32226 8942
rect 32174 8866 32226 8878
rect 33518 8930 33570 8942
rect 38110 8930 38162 8942
rect 37650 8878 37662 8930
rect 37714 8878 37726 8930
rect 33518 8866 33570 8878
rect 38110 8866 38162 8878
rect 1344 8650 44576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 44576 8650
rect 1344 8564 44576 8598
rect 9886 8370 9938 8382
rect 7746 8318 7758 8370
rect 7810 8318 7822 8370
rect 9886 8306 9938 8318
rect 15262 8370 15314 8382
rect 21422 8370 21474 8382
rect 15810 8318 15822 8370
rect 15874 8318 15886 8370
rect 18946 8318 18958 8370
rect 19010 8318 19022 8370
rect 15262 8306 15314 8318
rect 21422 8306 21474 8318
rect 23102 8370 23154 8382
rect 23102 8306 23154 8318
rect 15486 8258 15538 8270
rect 7074 8206 7086 8258
rect 7138 8206 7150 8258
rect 15486 8194 15538 8206
rect 18062 8258 18114 8270
rect 18062 8194 18114 8206
rect 18398 8258 18450 8270
rect 18398 8194 18450 8206
rect 19294 8258 19346 8270
rect 19294 8194 19346 8206
rect 19854 8258 19906 8270
rect 19854 8194 19906 8206
rect 20078 8258 20130 8270
rect 20078 8194 20130 8206
rect 20414 8258 20466 8270
rect 23426 8206 23438 8258
rect 23490 8206 23502 8258
rect 20414 8194 20466 8206
rect 18286 8146 18338 8158
rect 13458 8094 13470 8146
rect 13522 8094 13534 8146
rect 18286 8082 18338 8094
rect 10558 8034 10610 8046
rect 10558 7970 10610 7982
rect 13806 8034 13858 8046
rect 13806 7970 13858 7982
rect 17838 8034 17890 8046
rect 17838 7970 17890 7982
rect 18734 8034 18786 8046
rect 18734 7970 18786 7982
rect 18958 8034 19010 8046
rect 18958 7970 19010 7982
rect 20078 8034 20130 8046
rect 20078 7970 20130 7982
rect 23214 8034 23266 8046
rect 23214 7970 23266 7982
rect 23886 8034 23938 8046
rect 23886 7970 23938 7982
rect 1344 7866 44576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 44576 7866
rect 1344 7780 44576 7814
rect 25342 7698 25394 7710
rect 25342 7634 25394 7646
rect 32062 7698 32114 7710
rect 32062 7634 32114 7646
rect 22530 7534 22542 7586
rect 22594 7534 22606 7586
rect 32398 7474 32450 7486
rect 21858 7422 21870 7474
rect 21922 7422 21934 7474
rect 32398 7410 32450 7422
rect 24658 7310 24670 7362
rect 24722 7310 24734 7362
rect 1344 7082 44576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 44576 7082
rect 1344 6996 44576 7030
rect 33518 6690 33570 6702
rect 29810 6638 29822 6690
rect 29874 6638 29886 6690
rect 33518 6626 33570 6638
rect 14814 6578 14866 6590
rect 14814 6514 14866 6526
rect 15150 6578 15202 6590
rect 30382 6578 30434 6590
rect 18274 6526 18286 6578
rect 18338 6526 18350 6578
rect 15150 6514 15202 6526
rect 30382 6514 30434 6526
rect 32398 6578 32450 6590
rect 32398 6514 32450 6526
rect 18622 6466 18674 6478
rect 30818 6414 30830 6466
rect 30882 6414 30894 6466
rect 18622 6402 18674 6414
rect 1344 6298 44576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 44576 6298
rect 1344 6212 44576 6246
rect 20750 6130 20802 6142
rect 20750 6066 20802 6078
rect 25454 6130 25506 6142
rect 25454 6066 25506 6078
rect 26238 6130 26290 6142
rect 26238 6066 26290 6078
rect 30046 6130 30098 6142
rect 30046 6066 30098 6078
rect 30270 6130 30322 6142
rect 30270 6066 30322 6078
rect 31166 6130 31218 6142
rect 31166 6066 31218 6078
rect 36430 6130 36482 6142
rect 36430 6066 36482 6078
rect 28702 6018 28754 6030
rect 10882 5966 10894 6018
rect 10946 5966 10958 6018
rect 18162 5966 18174 6018
rect 18226 5966 18238 6018
rect 28702 5954 28754 5966
rect 28814 6018 28866 6030
rect 28814 5954 28866 5966
rect 29150 6018 29202 6030
rect 35186 5966 35198 6018
rect 35250 5966 35262 6018
rect 29150 5954 29202 5966
rect 13470 5906 13522 5918
rect 28478 5906 28530 5918
rect 10210 5854 10222 5906
rect 10274 5854 10286 5906
rect 17378 5854 17390 5906
rect 17442 5854 17454 5906
rect 27458 5854 27470 5906
rect 27522 5854 27534 5906
rect 13470 5842 13522 5854
rect 28478 5842 28530 5854
rect 29374 5906 29426 5918
rect 29374 5842 29426 5854
rect 29598 5906 29650 5918
rect 29598 5842 29650 5854
rect 30158 5906 30210 5918
rect 30594 5854 30606 5906
rect 30658 5854 30670 5906
rect 35970 5854 35982 5906
rect 36034 5854 36046 5906
rect 30158 5842 30210 5854
rect 25678 5794 25730 5806
rect 13010 5742 13022 5794
rect 13074 5742 13086 5794
rect 20290 5742 20302 5794
rect 20354 5742 20366 5794
rect 25678 5730 25730 5742
rect 26798 5794 26850 5806
rect 29262 5794 29314 5806
rect 27682 5742 27694 5794
rect 27746 5742 27758 5794
rect 33058 5742 33070 5794
rect 33122 5742 33134 5794
rect 26798 5730 26850 5742
rect 29262 5730 29314 5742
rect 25342 5682 25394 5694
rect 25342 5618 25394 5630
rect 1344 5514 44576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 44576 5514
rect 1344 5428 44576 5462
rect 27806 5234 27858 5246
rect 32622 5234 32674 5246
rect 25218 5182 25230 5234
rect 25282 5182 25294 5234
rect 27346 5182 27358 5234
rect 27410 5182 27422 5234
rect 29138 5182 29150 5234
rect 29202 5182 29214 5234
rect 31266 5182 31278 5234
rect 31330 5182 31342 5234
rect 27806 5170 27858 5182
rect 32622 5170 32674 5182
rect 15922 5070 15934 5122
rect 15986 5070 15998 5122
rect 19730 5070 19742 5122
rect 19794 5070 19806 5122
rect 24546 5070 24558 5122
rect 24610 5070 24622 5122
rect 31938 5070 31950 5122
rect 32002 5070 32014 5122
rect 16034 4958 16046 5010
rect 16098 4958 16110 5010
rect 19618 4958 19630 5010
rect 19682 4958 19694 5010
rect 16930 4846 16942 4898
rect 16994 4846 17006 4898
rect 1344 4730 44576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 44576 4730
rect 1344 4644 44576 4678
rect 22990 4562 23042 4574
rect 22990 4498 23042 4510
rect 13122 4398 13134 4450
rect 13186 4398 13198 4450
rect 21746 4398 21758 4450
rect 21810 4398 21822 4450
rect 15710 4338 15762 4350
rect 12450 4286 12462 4338
rect 12514 4286 12526 4338
rect 22530 4286 22542 4338
rect 22594 4286 22606 4338
rect 15710 4274 15762 4286
rect 15250 4174 15262 4226
rect 15314 4174 15326 4226
rect 19618 4174 19630 4226
rect 19682 4174 19694 4226
rect 1344 3946 44576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 44576 3946
rect 1344 3860 44576 3894
rect 1344 3162 44576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 44576 3162
rect 1344 3076 44576 3110
<< via1 >>
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 18286 42142 18338 42194
rect 33518 42142 33570 42194
rect 6190 42030 6242 42082
rect 9998 42030 10050 42082
rect 5070 41918 5122 41970
rect 5854 41918 5906 41970
rect 8878 41918 8930 41970
rect 9662 41918 9714 41970
rect 13470 41918 13522 41970
rect 17278 41918 17330 41970
rect 21086 41918 21138 41970
rect 24894 41918 24946 41970
rect 28702 41918 28754 41970
rect 30382 41918 30434 41970
rect 32510 41918 32562 41970
rect 36318 41918 36370 41970
rect 40126 41918 40178 41970
rect 14478 41806 14530 41858
rect 22094 41806 22146 41858
rect 25902 41806 25954 41858
rect 37326 41806 37378 41858
rect 41134 41806 41186 41858
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 43150 41358 43202 41410
rect 43934 41134 43986 41186
rect 39790 40910 39842 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 15710 40574 15762 40626
rect 16718 40574 16770 40626
rect 11566 40462 11618 40514
rect 12126 40462 12178 40514
rect 12350 40462 12402 40514
rect 14702 40462 14754 40514
rect 15486 40462 15538 40514
rect 16942 40462 16994 40514
rect 2270 40350 2322 40402
rect 2942 40350 2994 40402
rect 5630 40350 5682 40402
rect 6190 40350 6242 40402
rect 9774 40350 9826 40402
rect 11342 40350 11394 40402
rect 11678 40350 11730 40402
rect 12574 40350 12626 40402
rect 14366 40350 14418 40402
rect 15374 40350 15426 40402
rect 16606 40350 16658 40402
rect 20078 40350 20130 40402
rect 20302 40350 20354 40402
rect 25342 40350 25394 40402
rect 28590 40350 28642 40402
rect 31950 40350 32002 40402
rect 37438 40350 37490 40402
rect 40462 40350 40514 40402
rect 41022 40350 41074 40402
rect 5070 40238 5122 40290
rect 6862 40238 6914 40290
rect 8990 40238 9042 40290
rect 12462 40238 12514 40290
rect 21086 40238 21138 40290
rect 23214 40238 23266 40290
rect 26014 40238 26066 40290
rect 28142 40238 28194 40290
rect 29262 40238 29314 40290
rect 31390 40238 31442 40290
rect 34638 40238 34690 40290
rect 36766 40238 36818 40290
rect 38110 40238 38162 40290
rect 41806 40238 41858 40290
rect 43934 40238 43986 40290
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 11230 39678 11282 39730
rect 12014 39678 12066 39730
rect 16046 39678 16098 39730
rect 20750 39678 20802 39730
rect 21422 39678 21474 39730
rect 31614 39678 31666 39730
rect 33742 39678 33794 39730
rect 40798 39678 40850 39730
rect 41246 39678 41298 39730
rect 42702 39678 42754 39730
rect 11006 39566 11058 39618
rect 14254 39566 14306 39618
rect 14926 39566 14978 39618
rect 15262 39566 15314 39618
rect 15598 39566 15650 39618
rect 17838 39566 17890 39618
rect 18622 39566 18674 39618
rect 28366 39566 28418 39618
rect 30942 39566 30994 39618
rect 34190 39566 34242 39618
rect 37886 39566 37938 39618
rect 7982 39454 8034 39506
rect 8318 39454 8370 39506
rect 14030 39454 14082 39506
rect 16830 39454 16882 39506
rect 38670 39454 38722 39506
rect 10670 39342 10722 39394
rect 11678 39342 11730 39394
rect 11902 39342 11954 39394
rect 12126 39342 12178 39394
rect 14590 39342 14642 39394
rect 15486 39342 15538 39394
rect 15934 39342 15986 39394
rect 16158 39342 16210 39394
rect 16382 39342 16434 39394
rect 16942 39342 16994 39394
rect 17054 39342 17106 39394
rect 37550 39342 37602 39394
rect 41134 39342 41186 39394
rect 42590 39342 42642 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 13918 39006 13970 39058
rect 15150 39006 15202 39058
rect 15710 39006 15762 39058
rect 12574 38894 12626 38946
rect 12686 38894 12738 38946
rect 15486 38894 15538 38946
rect 13806 38782 13858 38834
rect 14030 38782 14082 38834
rect 14478 38782 14530 38834
rect 15038 38782 15090 38834
rect 15822 38670 15874 38722
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 2718 38110 2770 38162
rect 4846 38110 4898 38162
rect 7198 38110 7250 38162
rect 9326 38110 9378 38162
rect 25566 38110 25618 38162
rect 26014 38110 26066 38162
rect 31950 38110 32002 38162
rect 37102 38110 37154 38162
rect 2046 37998 2098 38050
rect 6414 37998 6466 38050
rect 12014 37998 12066 38050
rect 22766 37998 22818 38050
rect 34862 37998 34914 38050
rect 39454 37998 39506 38050
rect 39566 37998 39618 38050
rect 11678 37886 11730 37938
rect 23438 37886 23490 37938
rect 34078 37886 34130 37938
rect 36990 37886 37042 37938
rect 37326 37886 37378 37938
rect 37550 37886 37602 37938
rect 39902 37886 39954 37938
rect 5742 37774 5794 37826
rect 9774 37774 9826 37826
rect 11790 37774 11842 37826
rect 12462 37774 12514 37826
rect 35310 37774 35362 37826
rect 39790 37774 39842 37826
rect 40798 37774 40850 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 10670 37438 10722 37490
rect 11118 37438 11170 37490
rect 39006 37438 39058 37490
rect 39790 37438 39842 37490
rect 3726 37326 3778 37378
rect 9886 37326 9938 37378
rect 10334 37326 10386 37378
rect 12238 37326 12290 37378
rect 14254 37326 14306 37378
rect 16270 37326 16322 37378
rect 25566 37326 25618 37378
rect 39902 37326 39954 37378
rect 41918 37326 41970 37378
rect 3054 37214 3106 37266
rect 11006 37214 11058 37266
rect 11230 37214 11282 37266
rect 11566 37214 11618 37266
rect 12350 37214 12402 37266
rect 14478 37214 14530 37266
rect 15598 37214 15650 37266
rect 25230 37214 25282 37266
rect 31614 37214 31666 37266
rect 32062 37214 32114 37266
rect 38558 37214 38610 37266
rect 38782 37214 38834 37266
rect 39230 37214 39282 37266
rect 39566 37214 39618 37266
rect 40238 37214 40290 37266
rect 41246 37214 41298 37266
rect 5854 37102 5906 37154
rect 6302 37102 6354 37154
rect 16718 37102 16770 37154
rect 19630 37102 19682 37154
rect 28702 37102 28754 37154
rect 30830 37102 30882 37154
rect 34414 37102 34466 37154
rect 38446 37102 38498 37154
rect 40350 37102 40402 37154
rect 44046 37102 44098 37154
rect 9998 36990 10050 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 14254 36654 14306 36706
rect 25566 36654 25618 36706
rect 6974 36542 7026 36594
rect 12014 36542 12066 36594
rect 12350 36542 12402 36594
rect 12910 36542 12962 36594
rect 14814 36542 14866 36594
rect 24558 36542 24610 36594
rect 32286 36542 32338 36594
rect 33854 36542 33906 36594
rect 34526 36542 34578 36594
rect 35422 36542 35474 36594
rect 37438 36542 37490 36594
rect 39454 36542 39506 36594
rect 12574 36430 12626 36482
rect 13470 36430 13522 36482
rect 13806 36430 13858 36482
rect 14478 36430 14530 36482
rect 15486 36430 15538 36482
rect 18398 36430 18450 36482
rect 19070 36430 19122 36482
rect 19294 36430 19346 36482
rect 24782 36430 24834 36482
rect 26462 36430 26514 36482
rect 34078 36430 34130 36482
rect 34414 36430 34466 36482
rect 34638 36430 34690 36482
rect 39342 36430 39394 36482
rect 13694 36318 13746 36370
rect 15038 36318 15090 36370
rect 19966 36318 20018 36370
rect 20302 36318 20354 36370
rect 24110 36318 24162 36370
rect 25790 36318 25842 36370
rect 26350 36318 26402 36370
rect 33518 36318 33570 36370
rect 33742 36318 33794 36370
rect 34974 36318 35026 36370
rect 7086 36206 7138 36258
rect 14814 36206 14866 36258
rect 18062 36206 18114 36258
rect 18286 36206 18338 36258
rect 18734 36206 18786 36258
rect 25678 36206 25730 36258
rect 26126 36206 26178 36258
rect 32398 36206 32450 36258
rect 33854 36206 33906 36258
rect 37102 36206 37154 36258
rect 37326 36206 37378 36258
rect 37550 36206 37602 36258
rect 39118 36206 39170 36258
rect 39566 36206 39618 36258
rect 40014 36206 40066 36258
rect 40574 36206 40626 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 10782 35870 10834 35922
rect 13582 35870 13634 35922
rect 14590 35870 14642 35922
rect 34414 35870 34466 35922
rect 36654 35870 36706 35922
rect 10222 35758 10274 35810
rect 13022 35758 13074 35810
rect 14702 35758 14754 35810
rect 15486 35758 15538 35810
rect 17726 35758 17778 35810
rect 20974 35758 21026 35810
rect 26910 35758 26962 35810
rect 34638 35758 34690 35810
rect 13246 35646 13298 35698
rect 14590 35646 14642 35698
rect 17278 35646 17330 35698
rect 18174 35646 18226 35698
rect 19182 35646 19234 35698
rect 19518 35646 19570 35698
rect 19966 35646 20018 35698
rect 20078 35646 20130 35698
rect 20302 35646 20354 35698
rect 21646 35646 21698 35698
rect 25230 35646 25282 35698
rect 25902 35646 25954 35698
rect 34750 35646 34802 35698
rect 36542 35646 36594 35698
rect 36766 35646 36818 35698
rect 37214 35646 37266 35698
rect 21758 35534 21810 35586
rect 27358 35534 27410 35586
rect 36206 35534 36258 35586
rect 10446 35422 10498 35474
rect 18846 35422 18898 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 16606 35086 16658 35138
rect 18286 35086 18338 35138
rect 18622 35086 18674 35138
rect 37438 35086 37490 35138
rect 40910 35086 40962 35138
rect 14814 34974 14866 35026
rect 16718 34974 16770 35026
rect 19294 34974 19346 35026
rect 20750 34974 20802 35026
rect 25902 34974 25954 35026
rect 15038 34862 15090 34914
rect 19742 34862 19794 34914
rect 21310 34862 21362 34914
rect 25790 34862 25842 34914
rect 26014 34862 26066 34914
rect 28142 34862 28194 34914
rect 28366 34862 28418 34914
rect 29038 34862 29090 34914
rect 29374 34862 29426 34914
rect 35086 34862 35138 34914
rect 35646 34862 35698 34914
rect 14814 34750 14866 34802
rect 18398 34750 18450 34802
rect 19518 34750 19570 34802
rect 19966 34750 20018 34802
rect 20078 34750 20130 34802
rect 26238 34750 26290 34802
rect 27470 34750 27522 34802
rect 37326 34750 37378 34802
rect 40238 34750 40290 34802
rect 40350 34750 40402 34802
rect 40798 34750 40850 34802
rect 14590 34638 14642 34690
rect 18958 34638 19010 34690
rect 21646 34638 21698 34690
rect 29262 34638 29314 34690
rect 37438 34638 37490 34690
rect 40574 34638 40626 34690
rect 40910 34638 40962 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 13918 34302 13970 34354
rect 14254 34302 14306 34354
rect 19070 34302 19122 34354
rect 19182 34190 19234 34242
rect 37438 34190 37490 34242
rect 37102 34078 37154 34130
rect 41246 34078 41298 34130
rect 36766 33966 36818 34018
rect 40350 33966 40402 34018
rect 41918 33966 41970 34018
rect 44046 33966 44098 34018
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 41246 33518 41298 33570
rect 6638 33406 6690 33458
rect 33630 33406 33682 33458
rect 9550 33294 9602 33346
rect 10334 33294 10386 33346
rect 11006 33294 11058 33346
rect 29374 33294 29426 33346
rect 33182 33294 33234 33346
rect 34078 33294 34130 33346
rect 40574 33294 40626 33346
rect 40910 33294 40962 33346
rect 41358 33294 41410 33346
rect 8766 33182 8818 33234
rect 34414 33182 34466 33234
rect 41582 33182 41634 33234
rect 41694 33182 41746 33234
rect 42142 33182 42194 33234
rect 9998 33070 10050 33122
rect 10446 33070 10498 33122
rect 10558 33070 10610 33122
rect 11454 33070 11506 33122
rect 29150 33070 29202 33122
rect 40462 33070 40514 33122
rect 41134 33070 41186 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 8318 32734 8370 32786
rect 9774 32734 9826 32786
rect 24334 32734 24386 32786
rect 8430 32622 8482 32674
rect 8990 32622 9042 32674
rect 24222 32622 24274 32674
rect 25230 32622 25282 32674
rect 32510 32622 32562 32674
rect 2718 32510 2770 32562
rect 8094 32510 8146 32562
rect 25342 32510 25394 32562
rect 25454 32510 25506 32562
rect 25678 32510 25730 32562
rect 32286 32510 32338 32562
rect 33182 32510 33234 32562
rect 36430 32510 36482 32562
rect 3390 32398 3442 32450
rect 5518 32398 5570 32450
rect 5966 32398 6018 32450
rect 10334 32398 10386 32450
rect 33854 32398 33906 32450
rect 35982 32398 36034 32450
rect 8878 32286 8930 32338
rect 24446 32286 24498 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 5070 31838 5122 31890
rect 13470 31838 13522 31890
rect 16830 31838 16882 31890
rect 24894 31838 24946 31890
rect 33406 31838 33458 31890
rect 2270 31726 2322 31778
rect 16382 31726 16434 31778
rect 25006 31726 25058 31778
rect 33854 31726 33906 31778
rect 34302 31726 34354 31778
rect 39342 31726 39394 31778
rect 2942 31614 2994 31666
rect 15598 31614 15650 31666
rect 24110 31614 24162 31666
rect 24446 31614 24498 31666
rect 24782 31614 24834 31666
rect 25230 31614 25282 31666
rect 32958 31614 33010 31666
rect 33294 31614 33346 31666
rect 33966 31614 34018 31666
rect 34638 31614 34690 31666
rect 34750 31614 34802 31666
rect 37326 31614 37378 31666
rect 38782 31614 38834 31666
rect 39006 31614 39058 31666
rect 5742 31502 5794 31554
rect 33518 31502 33570 31554
rect 34190 31502 34242 31554
rect 34974 31502 35026 31554
rect 36542 31502 36594 31554
rect 36990 31502 37042 31554
rect 39230 31502 39282 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 15822 31166 15874 31218
rect 24222 31166 24274 31218
rect 10446 31054 10498 31106
rect 24446 31054 24498 31106
rect 24558 31054 24610 31106
rect 15486 30942 15538 30994
rect 21422 30942 21474 30994
rect 30270 30942 30322 30994
rect 32622 30942 32674 30994
rect 33182 30942 33234 30994
rect 15934 30830 15986 30882
rect 16494 30830 16546 30882
rect 18286 30830 18338 30882
rect 18622 30830 18674 30882
rect 20750 30830 20802 30882
rect 23998 30830 24050 30882
rect 27358 30830 27410 30882
rect 29486 30830 29538 30882
rect 30718 30830 30770 30882
rect 36878 30830 36930 30882
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 8766 30382 8818 30434
rect 9102 30270 9154 30322
rect 16830 30270 16882 30322
rect 24558 30270 24610 30322
rect 37438 30270 37490 30322
rect 39566 30270 39618 30322
rect 8766 30158 8818 30210
rect 9662 30158 9714 30210
rect 10110 30158 10162 30210
rect 10670 30158 10722 30210
rect 13582 30158 13634 30210
rect 16046 30158 16098 30210
rect 24894 30158 24946 30210
rect 28142 30158 28194 30210
rect 28366 30158 28418 30210
rect 29374 30158 29426 30210
rect 37102 30158 37154 30210
rect 40350 30158 40402 30210
rect 14030 30046 14082 30098
rect 25342 30046 25394 30098
rect 28590 30046 28642 30098
rect 31390 30046 31442 30098
rect 42702 30046 42754 30098
rect 20302 29934 20354 29986
rect 42590 29934 42642 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 5070 29598 5122 29650
rect 17502 29598 17554 29650
rect 18622 29598 18674 29650
rect 18958 29598 19010 29650
rect 19630 29598 19682 29650
rect 28366 29598 28418 29650
rect 29934 29598 29986 29650
rect 33182 29598 33234 29650
rect 37550 29598 37602 29650
rect 38782 29598 38834 29650
rect 38894 29598 38946 29650
rect 39118 29598 39170 29650
rect 40350 29598 40402 29650
rect 5630 29486 5682 29538
rect 8654 29486 8706 29538
rect 10782 29486 10834 29538
rect 14478 29486 14530 29538
rect 15486 29486 15538 29538
rect 16158 29486 16210 29538
rect 17614 29486 17666 29538
rect 19854 29486 19906 29538
rect 25230 29486 25282 29538
rect 29150 29486 29202 29538
rect 29374 29486 29426 29538
rect 33070 29486 33122 29538
rect 36654 29486 36706 29538
rect 37662 29486 37714 29538
rect 38670 29486 38722 29538
rect 3726 29374 3778 29426
rect 3950 29374 4002 29426
rect 4398 29374 4450 29426
rect 4622 29374 4674 29426
rect 4846 29374 4898 29426
rect 5182 29374 5234 29426
rect 8990 29374 9042 29426
rect 9998 29374 10050 29426
rect 10558 29374 10610 29426
rect 11454 29374 11506 29426
rect 11902 29374 11954 29426
rect 12126 29374 12178 29426
rect 14366 29374 14418 29426
rect 16270 29374 16322 29426
rect 16382 29374 16434 29426
rect 17390 29374 17442 29426
rect 17838 29374 17890 29426
rect 18062 29374 18114 29426
rect 18846 29374 18898 29426
rect 19070 29374 19122 29426
rect 19294 29374 19346 29426
rect 25566 29374 25618 29426
rect 36318 29374 36370 29426
rect 41134 29374 41186 29426
rect 3838 29262 3890 29314
rect 6078 29262 6130 29314
rect 9662 29262 9714 29314
rect 12686 29262 12738 29314
rect 15598 29262 15650 29314
rect 16830 29262 16882 29314
rect 19966 29262 20018 29314
rect 20302 29262 20354 29314
rect 25342 29262 25394 29314
rect 26014 29262 26066 29314
rect 28814 29262 28866 29314
rect 29486 29262 29538 29314
rect 35982 29262 36034 29314
rect 41918 29262 41970 29314
rect 44046 29262 44098 29314
rect 5518 29150 5570 29202
rect 11678 29150 11730 29202
rect 15710 29150 15762 29202
rect 33182 29150 33234 29202
rect 37550 29150 37602 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 3278 28814 3330 28866
rect 4286 28814 4338 28866
rect 5182 28814 5234 28866
rect 6414 28814 6466 28866
rect 9662 28814 9714 28866
rect 41246 28814 41298 28866
rect 6974 28702 7026 28754
rect 17278 28702 17330 28754
rect 18398 28702 18450 28754
rect 23550 28702 23602 28754
rect 25678 28702 25730 28754
rect 31054 28702 31106 28754
rect 33182 28702 33234 28754
rect 35086 28702 35138 28754
rect 40014 28702 40066 28754
rect 40462 28702 40514 28754
rect 41694 28702 41746 28754
rect 3166 28590 3218 28642
rect 4510 28590 4562 28642
rect 4734 28590 4786 28642
rect 5966 28590 6018 28642
rect 7982 28590 8034 28642
rect 8766 28590 8818 28642
rect 8878 28590 8930 28642
rect 9214 28590 9266 28642
rect 9886 28590 9938 28642
rect 10446 28590 10498 28642
rect 11230 28590 11282 28642
rect 11566 28590 11618 28642
rect 12574 28590 12626 28642
rect 13470 28590 13522 28642
rect 13918 28590 13970 28642
rect 16046 28590 16098 28642
rect 16270 28590 16322 28642
rect 16382 28590 16434 28642
rect 22878 28590 22930 28642
rect 26126 28590 26178 28642
rect 30270 28590 30322 28642
rect 33742 28590 33794 28642
rect 33966 28590 34018 28642
rect 34190 28590 34242 28642
rect 35422 28590 35474 28642
rect 41134 28590 41186 28642
rect 41470 28590 41522 28642
rect 3502 28478 3554 28530
rect 3726 28478 3778 28530
rect 4062 28478 4114 28530
rect 6414 28478 6466 28530
rect 6526 28478 6578 28530
rect 8318 28478 8370 28530
rect 9102 28478 9154 28530
rect 10782 28478 10834 28530
rect 12014 28478 12066 28530
rect 33518 28478 33570 28530
rect 35758 28478 35810 28530
rect 41806 28478 41858 28530
rect 2942 28366 2994 28418
rect 5630 28366 5682 28418
rect 7870 28366 7922 28418
rect 8206 28366 8258 28418
rect 16830 28366 16882 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 3614 28030 3666 28082
rect 4510 28030 4562 28082
rect 4622 28030 4674 28082
rect 5070 28030 5122 28082
rect 10558 28030 10610 28082
rect 10894 28030 10946 28082
rect 18174 28030 18226 28082
rect 41358 28030 41410 28082
rect 4174 27918 4226 27970
rect 5406 27918 5458 27970
rect 9998 27918 10050 27970
rect 17390 27918 17442 27970
rect 18062 27918 18114 27970
rect 4286 27806 4338 27858
rect 4734 27806 4786 27858
rect 9550 27806 9602 27858
rect 9774 27806 9826 27858
rect 10110 27806 10162 27858
rect 17614 27806 17666 27858
rect 17838 27806 17890 27858
rect 40350 27806 40402 27858
rect 41134 27806 41186 27858
rect 15486 27694 15538 27746
rect 21870 27694 21922 27746
rect 33182 27694 33234 27746
rect 33630 27694 33682 27746
rect 41470 27582 41522 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 14142 27134 14194 27186
rect 15038 27134 15090 27186
rect 15822 27134 15874 27186
rect 16158 27134 16210 27186
rect 20302 27134 20354 27186
rect 21758 27134 21810 27186
rect 25454 27134 25506 27186
rect 26350 27134 26402 27186
rect 36430 27134 36482 27186
rect 39902 27134 39954 27186
rect 41022 27134 41074 27186
rect 41470 27134 41522 27186
rect 14926 27022 14978 27074
rect 15262 27022 15314 27074
rect 17166 27022 17218 27074
rect 17726 27022 17778 27074
rect 22542 27022 22594 27074
rect 25902 27022 25954 27074
rect 35422 27022 35474 27074
rect 37102 27022 37154 27074
rect 40798 27022 40850 27074
rect 14478 26910 14530 26962
rect 20526 26910 20578 26962
rect 20638 26910 20690 26962
rect 21310 26910 21362 26962
rect 22206 26910 22258 26962
rect 29374 26910 29426 26962
rect 29710 26910 29762 26962
rect 30270 26910 30322 26962
rect 39454 26910 39506 26962
rect 17278 26798 17330 26850
rect 17390 26798 17442 26850
rect 20862 26798 20914 26850
rect 35086 26798 35138 26850
rect 35310 26798 35362 26850
rect 37438 26798 37490 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 6638 26462 6690 26514
rect 14366 26462 14418 26514
rect 18846 26462 18898 26514
rect 19854 26462 19906 26514
rect 37214 26462 37266 26514
rect 37662 26462 37714 26514
rect 3838 26350 3890 26402
rect 6414 26350 6466 26402
rect 10782 26350 10834 26402
rect 14478 26350 14530 26402
rect 15262 26350 15314 26402
rect 15822 26350 15874 26402
rect 17726 26350 17778 26402
rect 20974 26350 21026 26402
rect 5966 26238 6018 26290
rect 12238 26238 12290 26290
rect 12686 26238 12738 26290
rect 16046 26238 16098 26290
rect 17390 26238 17442 26290
rect 17614 26238 17666 26290
rect 18174 26238 18226 26290
rect 18510 26238 18562 26290
rect 18734 26238 18786 26290
rect 18958 26238 19010 26290
rect 19182 26238 19234 26290
rect 20190 26238 20242 26290
rect 26798 26238 26850 26290
rect 33966 26238 34018 26290
rect 37438 26238 37490 26290
rect 6526 26126 6578 26178
rect 16158 26126 16210 26178
rect 23102 26126 23154 26178
rect 27470 26126 27522 26178
rect 29598 26126 29650 26178
rect 30046 26126 30098 26178
rect 34750 26126 34802 26178
rect 36878 26126 36930 26178
rect 37326 26126 37378 26178
rect 40126 26126 40178 26178
rect 3726 26014 3778 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 6302 25678 6354 25730
rect 6526 25678 6578 25730
rect 12238 25678 12290 25730
rect 12462 25678 12514 25730
rect 17614 25678 17666 25730
rect 8878 25566 8930 25618
rect 27134 25566 27186 25618
rect 27582 25566 27634 25618
rect 34974 25566 35026 25618
rect 35422 25566 35474 25618
rect 37214 25566 37266 25618
rect 39902 25566 39954 25618
rect 44046 25566 44098 25618
rect 5518 25454 5570 25506
rect 5966 25454 6018 25506
rect 8654 25454 8706 25506
rect 11790 25454 11842 25506
rect 12686 25454 12738 25506
rect 14366 25454 14418 25506
rect 15598 25454 15650 25506
rect 17502 25454 17554 25506
rect 24222 25454 24274 25506
rect 24894 25454 24946 25506
rect 28254 25454 28306 25506
rect 29374 25454 29426 25506
rect 29710 25454 29762 25506
rect 35198 25454 35250 25506
rect 35870 25454 35922 25506
rect 40014 25454 40066 25506
rect 40462 25454 40514 25506
rect 41134 25454 41186 25506
rect 6190 25342 6242 25394
rect 8990 25342 9042 25394
rect 12910 25342 12962 25394
rect 17166 25342 17218 25394
rect 18174 25342 18226 25394
rect 24446 25342 24498 25394
rect 27806 25342 27858 25394
rect 29262 25342 29314 25394
rect 35646 25342 35698 25394
rect 40686 25342 40738 25394
rect 41918 25342 41970 25394
rect 5742 25230 5794 25282
rect 6750 25230 6802 25282
rect 27470 25230 27522 25282
rect 27694 25230 27746 25282
rect 29150 25230 29202 25282
rect 30158 25230 30210 25282
rect 40574 25230 40626 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 16046 24894 16098 24946
rect 18958 24894 19010 24946
rect 28926 24894 28978 24946
rect 38222 24894 38274 24946
rect 41358 24894 41410 24946
rect 12462 24782 12514 24834
rect 16158 24782 16210 24834
rect 40910 24782 40962 24834
rect 7646 24670 7698 24722
rect 8206 24670 8258 24722
rect 12350 24670 12402 24722
rect 14478 24670 14530 24722
rect 32510 24670 32562 24722
rect 33182 24670 33234 24722
rect 33406 24670 33458 24722
rect 33742 24670 33794 24722
rect 38446 24670 38498 24722
rect 38782 24670 38834 24722
rect 41246 24670 41298 24722
rect 41582 24670 41634 24722
rect 28478 24558 28530 24610
rect 33518 24558 33570 24610
rect 38334 24558 38386 24610
rect 40350 24558 40402 24610
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 29710 24110 29762 24162
rect 29934 24110 29986 24162
rect 35758 24110 35810 24162
rect 2942 23998 2994 24050
rect 5070 23998 5122 24050
rect 6414 23998 6466 24050
rect 7310 23998 7362 24050
rect 16942 23998 16994 24050
rect 23438 23998 23490 24050
rect 23886 23998 23938 24050
rect 29934 23998 29986 24050
rect 31726 23998 31778 24050
rect 33854 23998 33906 24050
rect 34302 23998 34354 24050
rect 35534 23998 35586 24050
rect 35870 23998 35922 24050
rect 2270 23886 2322 23938
rect 5854 23886 5906 23938
rect 6862 23886 6914 23938
rect 10782 23886 10834 23938
rect 11118 23886 11170 23938
rect 15150 23886 15202 23938
rect 17166 23886 17218 23938
rect 19294 23886 19346 23938
rect 22878 23886 22930 23938
rect 24334 23886 24386 23938
rect 24894 23886 24946 23938
rect 29262 23886 29314 23938
rect 31054 23886 31106 23938
rect 11678 23774 11730 23826
rect 16270 23774 16322 23826
rect 17726 23774 17778 23826
rect 22766 23774 22818 23826
rect 7422 23662 7474 23714
rect 10446 23662 10498 23714
rect 11342 23662 11394 23714
rect 19630 23662 19682 23714
rect 22542 23662 22594 23714
rect 24558 23662 24610 23714
rect 25230 23662 25282 23714
rect 29486 23662 29538 23714
rect 40686 23662 40738 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 15934 23326 15986 23378
rect 19070 23326 19122 23378
rect 21534 23326 21586 23378
rect 22654 23326 22706 23378
rect 26686 23326 26738 23378
rect 33406 23326 33458 23378
rect 39118 23326 39170 23378
rect 41470 23326 41522 23378
rect 3166 23214 3218 23266
rect 19182 23214 19234 23266
rect 21086 23214 21138 23266
rect 29150 23214 29202 23266
rect 33070 23214 33122 23266
rect 33182 23214 33234 23266
rect 35870 23214 35922 23266
rect 37326 23214 37378 23266
rect 41806 23214 41858 23266
rect 2494 23102 2546 23154
rect 10782 23102 10834 23154
rect 11678 23102 11730 23154
rect 12686 23102 12738 23154
rect 13806 23102 13858 23154
rect 17502 23102 17554 23154
rect 19406 23102 19458 23154
rect 19854 23102 19906 23154
rect 20190 23102 20242 23154
rect 20414 23102 20466 23154
rect 20750 23102 20802 23154
rect 23326 23102 23378 23154
rect 23550 23102 23602 23154
rect 24446 23102 24498 23154
rect 25566 23102 25618 23154
rect 26014 23102 26066 23154
rect 26350 23102 26402 23154
rect 28926 23102 28978 23154
rect 29486 23102 29538 23154
rect 34974 23102 35026 23154
rect 35422 23102 35474 23154
rect 36654 23102 36706 23154
rect 36990 23102 37042 23154
rect 39454 23102 39506 23154
rect 39678 23102 39730 23154
rect 41134 23102 41186 23154
rect 41582 23102 41634 23154
rect 5294 22990 5346 23042
rect 5854 22990 5906 23042
rect 14478 22990 14530 23042
rect 16046 22990 16098 23042
rect 17950 22990 18002 23042
rect 23886 22990 23938 23042
rect 29934 22990 29986 23042
rect 36542 22990 36594 23042
rect 36878 22990 36930 23042
rect 40350 22990 40402 23042
rect 14702 22878 14754 22930
rect 22990 22878 23042 22930
rect 41246 22878 41298 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 16158 22542 16210 22594
rect 19406 22542 19458 22594
rect 40798 22542 40850 22594
rect 41134 22542 41186 22594
rect 15934 22430 15986 22482
rect 19630 22430 19682 22482
rect 26238 22430 26290 22482
rect 40014 22430 40066 22482
rect 13470 22318 13522 22370
rect 14366 22318 14418 22370
rect 17166 22318 17218 22370
rect 19070 22318 19122 22370
rect 21534 22318 21586 22370
rect 21758 22318 21810 22370
rect 40574 22318 40626 22370
rect 14478 22206 14530 22258
rect 15710 22206 15762 22258
rect 17054 22206 17106 22258
rect 41022 22206 41074 22258
rect 13694 22094 13746 22146
rect 13806 22094 13858 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 13582 21758 13634 21810
rect 15374 21758 15426 21810
rect 24670 21758 24722 21810
rect 25790 21758 25842 21810
rect 42590 21758 42642 21810
rect 10334 21646 10386 21698
rect 12910 21646 12962 21698
rect 18846 21646 18898 21698
rect 19070 21646 19122 21698
rect 26686 21646 26738 21698
rect 28926 21646 28978 21698
rect 29598 21646 29650 21698
rect 30046 21646 30098 21698
rect 37102 21646 37154 21698
rect 6862 21534 6914 21586
rect 7310 21534 7362 21586
rect 7422 21534 7474 21586
rect 9998 21534 10050 21586
rect 11342 21534 11394 21586
rect 13358 21534 13410 21586
rect 30158 21534 30210 21586
rect 36430 21534 36482 21586
rect 18958 21422 19010 21474
rect 25230 21422 25282 21474
rect 26126 21422 26178 21474
rect 39230 21422 39282 21474
rect 39790 21422 39842 21474
rect 42702 21422 42754 21474
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 29822 20974 29874 21026
rect 11342 20862 11394 20914
rect 16158 20862 16210 20914
rect 16942 20862 16994 20914
rect 26238 20862 26290 20914
rect 41470 20862 41522 20914
rect 43598 20862 43650 20914
rect 8430 20750 8482 20802
rect 9438 20750 9490 20802
rect 10558 20750 10610 20802
rect 10894 20750 10946 20802
rect 13806 20750 13858 20802
rect 15150 20750 15202 20802
rect 17054 20750 17106 20802
rect 25230 20750 25282 20802
rect 25678 20750 25730 20802
rect 30158 20750 30210 20802
rect 30382 20750 30434 20802
rect 30606 20750 30658 20802
rect 40686 20750 40738 20802
rect 9214 20638 9266 20690
rect 11230 20638 11282 20690
rect 14030 20638 14082 20690
rect 15038 20638 15090 20690
rect 17278 20638 17330 20690
rect 18062 20638 18114 20690
rect 8430 20526 8482 20578
rect 9326 20526 9378 20578
rect 10110 20526 10162 20578
rect 40350 20526 40402 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 8990 20190 9042 20242
rect 10222 20190 10274 20242
rect 15486 20190 15538 20242
rect 8542 20078 8594 20130
rect 9998 20078 10050 20130
rect 10446 20078 10498 20130
rect 14814 20078 14866 20130
rect 16046 20078 16098 20130
rect 8430 19966 8482 20018
rect 8878 19966 8930 20018
rect 10782 19966 10834 20018
rect 14590 19966 14642 20018
rect 15822 19966 15874 20018
rect 19742 19966 19794 20018
rect 19966 19966 20018 20018
rect 20414 19966 20466 20018
rect 29486 19966 29538 20018
rect 4958 19854 5010 19906
rect 10334 19854 10386 19906
rect 10894 19854 10946 19906
rect 19854 19854 19906 19906
rect 30158 19854 30210 19906
rect 32286 19854 32338 19906
rect 33182 19854 33234 19906
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 9886 19406 9938 19458
rect 15150 19406 15202 19458
rect 30158 19406 30210 19458
rect 30494 19406 30546 19458
rect 31278 19406 31330 19458
rect 4734 19294 4786 19346
rect 5742 19294 5794 19346
rect 17838 19294 17890 19346
rect 27582 19294 27634 19346
rect 28030 19294 28082 19346
rect 33518 19294 33570 19346
rect 1822 19182 1874 19234
rect 6078 19182 6130 19234
rect 20638 19182 20690 19234
rect 24110 19182 24162 19234
rect 24782 19182 24834 19234
rect 30270 19182 30322 19234
rect 30606 19182 30658 19234
rect 31726 19182 31778 19234
rect 31950 19182 32002 19234
rect 36430 19182 36482 19234
rect 2606 19070 2658 19122
rect 9774 19070 9826 19122
rect 15038 19070 15090 19122
rect 19966 19070 20018 19122
rect 24334 19070 24386 19122
rect 25454 19070 25506 19122
rect 35646 19070 35698 19122
rect 21422 18958 21474 19010
rect 29822 18958 29874 19010
rect 37102 18958 37154 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 10558 18622 10610 18674
rect 14254 18622 14306 18674
rect 14702 18622 14754 18674
rect 19518 18622 19570 18674
rect 20190 18622 20242 18674
rect 24558 18622 24610 18674
rect 31838 18622 31890 18674
rect 4062 18510 4114 18562
rect 10110 18510 10162 18562
rect 10670 18510 10722 18562
rect 14478 18510 14530 18562
rect 14814 18510 14866 18562
rect 19070 18510 19122 18562
rect 23214 18510 23266 18562
rect 23438 18510 23490 18562
rect 34526 18510 34578 18562
rect 5182 18398 5234 18450
rect 11006 18398 11058 18450
rect 13806 18398 13858 18450
rect 14366 18398 14418 18450
rect 15038 18398 15090 18450
rect 15486 18398 15538 18450
rect 15710 18398 15762 18450
rect 19294 18398 19346 18450
rect 19630 18398 19682 18450
rect 20750 18398 20802 18450
rect 22990 18398 23042 18450
rect 23550 18398 23602 18450
rect 23886 18398 23938 18450
rect 23998 18398 24050 18450
rect 24110 18398 24162 18450
rect 32174 18398 32226 18450
rect 33966 18398 34018 18450
rect 34302 18398 34354 18450
rect 3950 18286 4002 18338
rect 4846 18286 4898 18338
rect 5630 18286 5682 18338
rect 16158 18286 16210 18338
rect 22654 18286 22706 18338
rect 32398 18286 32450 18338
rect 34638 18286 34690 18338
rect 4286 18174 4338 18226
rect 15262 18174 15314 18226
rect 19518 18174 19570 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 4510 17726 4562 17778
rect 5966 17726 6018 17778
rect 12014 17726 12066 17778
rect 14702 17726 14754 17778
rect 16830 17726 16882 17778
rect 22878 17726 22930 17778
rect 23326 17726 23378 17778
rect 24446 17726 24498 17778
rect 5630 17614 5682 17666
rect 6078 17614 6130 17666
rect 9886 17614 9938 17666
rect 10110 17614 10162 17666
rect 10222 17614 10274 17666
rect 10446 17614 10498 17666
rect 11230 17614 11282 17666
rect 11454 17614 11506 17666
rect 14030 17614 14082 17666
rect 23438 17614 23490 17666
rect 23886 17614 23938 17666
rect 24334 17614 24386 17666
rect 32958 17614 33010 17666
rect 35758 17614 35810 17666
rect 11006 17502 11058 17554
rect 23214 17502 23266 17554
rect 32398 17502 32450 17554
rect 32846 17502 32898 17554
rect 35198 17502 35250 17554
rect 35310 17502 35362 17554
rect 35870 17502 35922 17554
rect 36990 17502 37042 17554
rect 5854 17390 5906 17442
rect 6190 17390 6242 17442
rect 9438 17390 9490 17442
rect 11118 17390 11170 17442
rect 17278 17390 17330 17442
rect 32286 17390 32338 17442
rect 35534 17390 35586 17442
rect 37326 17390 37378 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 17502 17054 17554 17106
rect 30494 17054 30546 17106
rect 30942 17054 30994 17106
rect 6750 16942 6802 16994
rect 9662 16942 9714 16994
rect 10222 16942 10274 16994
rect 31054 16942 31106 16994
rect 6078 16830 6130 16882
rect 15262 16830 15314 16882
rect 15710 16830 15762 16882
rect 17614 16830 17666 16882
rect 20190 16830 20242 16882
rect 20750 16830 20802 16882
rect 31614 16830 31666 16882
rect 32510 16830 32562 16882
rect 33070 16830 33122 16882
rect 8878 16718 8930 16770
rect 31950 16718 32002 16770
rect 37102 16718 37154 16770
rect 17502 16606 17554 16658
rect 30942 16606 30994 16658
rect 31614 16606 31666 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 23438 16270 23490 16322
rect 31054 16270 31106 16322
rect 34862 16270 34914 16322
rect 36430 16270 36482 16322
rect 10222 16158 10274 16210
rect 11006 16158 11058 16210
rect 31278 16158 31330 16210
rect 35870 16158 35922 16210
rect 37438 16158 37490 16210
rect 39566 16158 39618 16210
rect 9662 16046 9714 16098
rect 10558 16046 10610 16098
rect 10782 16046 10834 16098
rect 11230 16046 11282 16098
rect 11566 16046 11618 16098
rect 12910 16046 12962 16098
rect 13806 16046 13858 16098
rect 15710 16046 15762 16098
rect 23326 16046 23378 16098
rect 31390 16046 31442 16098
rect 34414 16046 34466 16098
rect 36094 16046 36146 16098
rect 40350 16046 40402 16098
rect 11006 15934 11058 15986
rect 11454 15934 11506 15986
rect 12574 15934 12626 15986
rect 13470 15934 13522 15986
rect 18398 15934 18450 15986
rect 33854 15934 33906 15986
rect 34302 15934 34354 15986
rect 34526 15934 34578 15986
rect 34974 15934 35026 15986
rect 35086 15934 35138 15986
rect 19966 15822 20018 15874
rect 22990 15822 23042 15874
rect 23438 15822 23490 15874
rect 37102 15822 37154 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 19854 15486 19906 15538
rect 25342 15486 25394 15538
rect 33182 15486 33234 15538
rect 35982 15486 36034 15538
rect 23214 15374 23266 15426
rect 23326 15374 23378 15426
rect 23550 15374 23602 15426
rect 23998 15374 24050 15426
rect 25790 15374 25842 15426
rect 27806 15374 27858 15426
rect 31726 15374 31778 15426
rect 35422 15374 35474 15426
rect 36878 15374 36930 15426
rect 19630 15262 19682 15314
rect 20750 15262 20802 15314
rect 23662 15262 23714 15314
rect 24222 15262 24274 15314
rect 24670 15262 24722 15314
rect 25230 15262 25282 15314
rect 29038 15262 29090 15314
rect 32510 15262 32562 15314
rect 34190 15262 34242 15314
rect 37998 15262 38050 15314
rect 20414 15150 20466 15202
rect 24446 15150 24498 15202
rect 24558 15150 24610 15202
rect 29598 15150 29650 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 23326 14702 23378 14754
rect 25454 14702 25506 14754
rect 5742 14590 5794 14642
rect 15150 14590 15202 14642
rect 20078 14590 20130 14642
rect 25006 14590 25058 14642
rect 25566 14590 25618 14642
rect 28702 14590 28754 14642
rect 31950 14590 32002 14642
rect 1934 14478 1986 14530
rect 22990 14478 23042 14530
rect 23662 14478 23714 14530
rect 24446 14478 24498 14530
rect 29150 14478 29202 14530
rect 2606 14366 2658 14418
rect 14254 14366 14306 14418
rect 14366 14366 14418 14418
rect 15486 14366 15538 14418
rect 24222 14366 24274 14418
rect 4846 14254 4898 14306
rect 6190 14254 6242 14306
rect 14590 14254 14642 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 9998 13918 10050 13970
rect 11678 13918 11730 13970
rect 12014 13918 12066 13970
rect 12462 13918 12514 13970
rect 14254 13918 14306 13970
rect 16046 13918 16098 13970
rect 30046 13918 30098 13970
rect 35422 13918 35474 13970
rect 35646 13918 35698 13970
rect 14926 13806 14978 13858
rect 15598 13806 15650 13858
rect 27246 13806 27298 13858
rect 9550 13694 9602 13746
rect 9774 13694 9826 13746
rect 10222 13694 10274 13746
rect 13694 13694 13746 13746
rect 14142 13694 14194 13746
rect 14366 13694 14418 13746
rect 14590 13694 14642 13746
rect 15374 13694 15426 13746
rect 26574 13694 26626 13746
rect 34974 13694 35026 13746
rect 36318 13694 36370 13746
rect 36542 13694 36594 13746
rect 5182 13582 5234 13634
rect 9886 13582 9938 13634
rect 15486 13582 15538 13634
rect 29374 13582 29426 13634
rect 34750 13582 34802 13634
rect 35534 13582 35586 13634
rect 15150 13470 15202 13522
rect 35982 13470 36034 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 24110 13134 24162 13186
rect 35870 13134 35922 13186
rect 5742 13022 5794 13074
rect 10222 13022 10274 13074
rect 12910 13022 12962 13074
rect 15038 13022 15090 13074
rect 15710 13022 15762 13074
rect 17838 13022 17890 13074
rect 21870 13022 21922 13074
rect 36094 13022 36146 13074
rect 36990 13022 37042 13074
rect 39118 13022 39170 13074
rect 6078 12910 6130 12962
rect 6414 12910 6466 12962
rect 6974 12910 7026 12962
rect 8430 12910 8482 12962
rect 9886 12910 9938 12962
rect 12238 12910 12290 12962
rect 14926 12910 14978 12962
rect 18622 12910 18674 12962
rect 23438 12910 23490 12962
rect 25678 12910 25730 12962
rect 39790 12910 39842 12962
rect 4958 12798 5010 12850
rect 5070 12798 5122 12850
rect 5630 12798 5682 12850
rect 5854 12798 5906 12850
rect 7422 12798 7474 12850
rect 8766 12798 8818 12850
rect 9774 12798 9826 12850
rect 12462 12798 12514 12850
rect 14590 12798 14642 12850
rect 23998 12798 24050 12850
rect 36094 12798 36146 12850
rect 7198 12686 7250 12738
rect 7534 12686 7586 12738
rect 19070 12686 19122 12738
rect 23774 12686 23826 12738
rect 24446 12686 24498 12738
rect 25454 12686 25506 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 5294 12350 5346 12402
rect 6638 12350 6690 12402
rect 8542 12350 8594 12402
rect 8654 12350 8706 12402
rect 8766 12350 8818 12402
rect 9774 12350 9826 12402
rect 11454 12350 11506 12402
rect 20750 12350 20802 12402
rect 22206 12350 22258 12402
rect 23438 12350 23490 12402
rect 24558 12350 24610 12402
rect 5518 12238 5570 12290
rect 8318 12238 8370 12290
rect 9550 12238 9602 12290
rect 11006 12238 11058 12290
rect 21086 12238 21138 12290
rect 22654 12238 22706 12290
rect 23662 12238 23714 12290
rect 24110 12238 24162 12290
rect 24670 12238 24722 12290
rect 5630 12126 5682 12178
rect 8990 12126 9042 12178
rect 9774 12126 9826 12178
rect 9998 12126 10050 12178
rect 10110 12126 10162 12178
rect 10670 12126 10722 12178
rect 20526 12126 20578 12178
rect 22094 12126 22146 12178
rect 22430 12126 22482 12178
rect 23102 12126 23154 12178
rect 23214 12126 23266 12178
rect 23998 12126 24050 12178
rect 24334 12126 24386 12178
rect 21646 12014 21698 12066
rect 22318 12014 22370 12066
rect 23774 12014 23826 12066
rect 36654 12014 36706 12066
rect 21310 11902 21362 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 13918 11454 13970 11506
rect 14926 11454 14978 11506
rect 22206 11454 22258 11506
rect 25230 11454 25282 11506
rect 34526 11454 34578 11506
rect 4398 11342 4450 11394
rect 4846 11342 4898 11394
rect 5742 11342 5794 11394
rect 6078 11342 6130 11394
rect 6638 11342 6690 11394
rect 6750 11342 6802 11394
rect 6862 11342 6914 11394
rect 14030 11342 14082 11394
rect 14254 11342 14306 11394
rect 14366 11342 14418 11394
rect 21758 11342 21810 11394
rect 21982 11342 22034 11394
rect 22430 11342 22482 11394
rect 22654 11342 22706 11394
rect 23662 11342 23714 11394
rect 23998 11342 24050 11394
rect 24334 11342 24386 11394
rect 24670 11342 24722 11394
rect 28142 11342 28194 11394
rect 34750 11342 34802 11394
rect 35422 11342 35474 11394
rect 4174 11230 4226 11282
rect 5070 11230 5122 11282
rect 5966 11230 6018 11282
rect 13918 11230 13970 11282
rect 23438 11230 23490 11282
rect 24222 11230 24274 11282
rect 27358 11230 27410 11282
rect 4286 11118 4338 11170
rect 5854 11118 5906 11170
rect 6190 11118 6242 11170
rect 7086 11118 7138 11170
rect 7646 11118 7698 11170
rect 28590 11118 28642 11170
rect 35198 11118 35250 11170
rect 35310 11118 35362 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 11678 10782 11730 10834
rect 12014 10782 12066 10834
rect 14366 10782 14418 10834
rect 15262 10782 15314 10834
rect 25342 10782 25394 10834
rect 31726 10782 31778 10834
rect 2606 10670 2658 10722
rect 13806 10670 13858 10722
rect 35422 10670 35474 10722
rect 35646 10670 35698 10722
rect 1934 10558 1986 10610
rect 11790 10558 11842 10610
rect 12126 10558 12178 10610
rect 13246 10558 13298 10610
rect 13582 10558 13634 10610
rect 14030 10558 14082 10610
rect 14590 10558 14642 10610
rect 14926 10558 14978 10610
rect 28478 10558 28530 10610
rect 34862 10558 34914 10610
rect 35086 10558 35138 10610
rect 4734 10446 4786 10498
rect 5182 10446 5234 10498
rect 11902 10446 11954 10498
rect 13918 10446 13970 10498
rect 14478 10446 14530 10498
rect 18286 10446 18338 10498
rect 19742 10446 19794 10498
rect 29150 10446 29202 10498
rect 31278 10446 31330 10498
rect 35534 10446 35586 10498
rect 34526 10334 34578 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 17278 9998 17330 10050
rect 20414 9998 20466 10050
rect 29598 9998 29650 10050
rect 29710 9998 29762 10050
rect 31390 9998 31442 10050
rect 11230 9886 11282 9938
rect 12910 9886 12962 9938
rect 15038 9886 15090 9938
rect 18734 9886 18786 9938
rect 12238 9774 12290 9826
rect 13806 9774 13858 9826
rect 14142 9774 14194 9826
rect 14926 9774 14978 9826
rect 17502 9774 17554 9826
rect 18286 9774 18338 9826
rect 19182 9774 19234 9826
rect 19630 9774 19682 9826
rect 29374 9774 29426 9826
rect 29934 9774 29986 9826
rect 30158 9774 30210 9826
rect 30606 9774 30658 9826
rect 31054 9774 31106 9826
rect 31838 9774 31890 9826
rect 32062 9774 32114 9826
rect 33966 9774 34018 9826
rect 11342 9662 11394 9714
rect 11566 9662 11618 9714
rect 12014 9662 12066 9714
rect 12350 9662 12402 9714
rect 14590 9662 14642 9714
rect 17838 9662 17890 9714
rect 18174 9662 18226 9714
rect 18846 9662 18898 9714
rect 30494 9662 30546 9714
rect 30830 9662 30882 9714
rect 31950 9662 32002 9714
rect 33742 9662 33794 9714
rect 12462 9550 12514 9602
rect 20190 9550 20242 9602
rect 20302 9550 20354 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 12462 9214 12514 9266
rect 12686 9214 12738 9266
rect 18622 9214 18674 9266
rect 18846 9214 18898 9266
rect 19854 9214 19906 9266
rect 31390 9214 31442 9266
rect 12798 9102 12850 9154
rect 20078 9102 20130 9154
rect 32062 9102 32114 9154
rect 33294 9102 33346 9154
rect 35534 9102 35586 9154
rect 17614 8990 17666 9042
rect 17838 8990 17890 9042
rect 18062 8990 18114 9042
rect 18398 8990 18450 9042
rect 18510 8990 18562 9042
rect 19630 8990 19682 9042
rect 31614 8990 31666 9042
rect 32286 8990 32338 9042
rect 33070 8990 33122 9042
rect 33742 8990 33794 9042
rect 34862 8990 34914 9042
rect 17950 8878 18002 8930
rect 19742 8878 19794 8930
rect 32174 8878 32226 8930
rect 33518 8878 33570 8930
rect 37662 8878 37714 8930
rect 38110 8878 38162 8930
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 7758 8318 7810 8370
rect 9886 8318 9938 8370
rect 15262 8318 15314 8370
rect 15822 8318 15874 8370
rect 18958 8318 19010 8370
rect 21422 8318 21474 8370
rect 23102 8318 23154 8370
rect 7086 8206 7138 8258
rect 15486 8206 15538 8258
rect 18062 8206 18114 8258
rect 18398 8206 18450 8258
rect 19294 8206 19346 8258
rect 19854 8206 19906 8258
rect 20078 8206 20130 8258
rect 20414 8206 20466 8258
rect 23438 8206 23490 8258
rect 13470 8094 13522 8146
rect 18286 8094 18338 8146
rect 10558 7982 10610 8034
rect 13806 7982 13858 8034
rect 17838 7982 17890 8034
rect 18734 7982 18786 8034
rect 18958 7982 19010 8034
rect 20078 7982 20130 8034
rect 23214 7982 23266 8034
rect 23886 7982 23938 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 25342 7646 25394 7698
rect 32062 7646 32114 7698
rect 22542 7534 22594 7586
rect 21870 7422 21922 7474
rect 32398 7422 32450 7474
rect 24670 7310 24722 7362
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 29822 6638 29874 6690
rect 33518 6638 33570 6690
rect 14814 6526 14866 6578
rect 15150 6526 15202 6578
rect 18286 6526 18338 6578
rect 30382 6526 30434 6578
rect 32398 6526 32450 6578
rect 18622 6414 18674 6466
rect 30830 6414 30882 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 20750 6078 20802 6130
rect 25454 6078 25506 6130
rect 26238 6078 26290 6130
rect 30046 6078 30098 6130
rect 30270 6078 30322 6130
rect 31166 6078 31218 6130
rect 36430 6078 36482 6130
rect 10894 5966 10946 6018
rect 18174 5966 18226 6018
rect 28702 5966 28754 6018
rect 28814 5966 28866 6018
rect 29150 5966 29202 6018
rect 35198 5966 35250 6018
rect 10222 5854 10274 5906
rect 13470 5854 13522 5906
rect 17390 5854 17442 5906
rect 27470 5854 27522 5906
rect 28478 5854 28530 5906
rect 29374 5854 29426 5906
rect 29598 5854 29650 5906
rect 30158 5854 30210 5906
rect 30606 5854 30658 5906
rect 35982 5854 36034 5906
rect 13022 5742 13074 5794
rect 20302 5742 20354 5794
rect 25678 5742 25730 5794
rect 26798 5742 26850 5794
rect 27694 5742 27746 5794
rect 29262 5742 29314 5794
rect 33070 5742 33122 5794
rect 25342 5630 25394 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 25230 5182 25282 5234
rect 27358 5182 27410 5234
rect 27806 5182 27858 5234
rect 29150 5182 29202 5234
rect 31278 5182 31330 5234
rect 32622 5182 32674 5234
rect 15934 5070 15986 5122
rect 19742 5070 19794 5122
rect 24558 5070 24610 5122
rect 31950 5070 32002 5122
rect 16046 4958 16098 5010
rect 19630 4958 19682 5010
rect 16942 4846 16994 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 22990 4510 23042 4562
rect 13134 4398 13186 4450
rect 21758 4398 21810 4450
rect 12462 4286 12514 4338
rect 15710 4286 15762 4338
rect 22542 4286 22594 4338
rect 15262 4174 15314 4226
rect 19630 4174 19682 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 1792 45200 1904 46000
rect 5600 45200 5712 46000
rect 9408 45200 9520 46000
rect 13216 45200 13328 46000
rect 17024 45200 17136 46000
rect 17388 45276 17892 45332
rect 1820 22148 1876 45200
rect 5628 43708 5684 45200
rect 9436 43708 9492 45200
rect 5628 43652 5908 43708
rect 9436 43652 9716 43708
rect 5068 41972 5124 41982
rect 5852 41972 5908 43652
rect 5068 41970 5908 41972
rect 5068 41918 5070 41970
rect 5122 41918 5854 41970
rect 5906 41918 5908 41970
rect 5068 41916 5908 41918
rect 5068 41906 5124 41916
rect 5852 41906 5908 41916
rect 6188 42082 6244 42094
rect 6188 42030 6190 42082
rect 6242 42030 6244 42082
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 6188 40628 6244 42030
rect 8876 41972 8932 41982
rect 9660 41972 9716 43652
rect 8876 41970 9716 41972
rect 8876 41918 8878 41970
rect 8930 41918 9662 41970
rect 9714 41918 9716 41970
rect 8876 41916 9716 41918
rect 8876 41906 8932 41916
rect 9660 41906 9716 41916
rect 9996 42082 10052 42094
rect 9996 42030 9998 42082
rect 10050 42030 10052 42082
rect 6188 40572 6580 40628
rect 2268 40402 2324 40414
rect 2268 40350 2270 40402
rect 2322 40350 2324 40402
rect 2044 38052 2100 38062
rect 2268 38052 2324 40350
rect 2940 40404 2996 40414
rect 2940 40310 2996 40348
rect 5628 40404 5684 40414
rect 6188 40404 6244 40414
rect 5628 40402 6244 40404
rect 5628 40350 5630 40402
rect 5682 40350 6190 40402
rect 6242 40350 6244 40402
rect 5628 40348 6244 40350
rect 5628 40338 5684 40348
rect 5068 40292 5124 40302
rect 5068 40198 5124 40236
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 2716 38948 2772 38958
rect 2716 38162 2772 38892
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 2716 38110 2718 38162
rect 2770 38110 2772 38162
rect 2716 38098 2772 38110
rect 4844 38162 4900 38174
rect 4844 38110 4846 38162
rect 4898 38110 4900 38162
rect 2044 38050 2324 38052
rect 2044 37998 2046 38050
rect 2098 37998 2324 38050
rect 2044 37996 2324 37998
rect 2044 37986 2100 37996
rect 2268 37828 2324 37996
rect 2268 37762 2324 37772
rect 3052 37828 3108 37838
rect 3052 37266 3108 37772
rect 3724 37380 3780 37390
rect 3724 37286 3780 37324
rect 3052 37214 3054 37266
rect 3106 37214 3108 37266
rect 3052 37202 3108 37214
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4844 35812 4900 38110
rect 6188 38052 6244 40348
rect 6412 38052 6468 38062
rect 6188 38050 6468 38052
rect 6188 37998 6414 38050
rect 6466 37998 6468 38050
rect 6188 37996 6468 37998
rect 5740 37828 5796 37838
rect 5740 37734 5796 37772
rect 6300 37828 6356 37996
rect 6412 37986 6468 37996
rect 5852 37154 5908 37166
rect 5852 37102 5854 37154
rect 5906 37102 5908 37154
rect 5852 36596 5908 37102
rect 5852 36530 5908 36540
rect 6300 37154 6356 37772
rect 6300 37102 6302 37154
rect 6354 37102 6356 37154
rect 4844 35746 4900 35756
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 2716 32562 2772 32574
rect 2716 32510 2718 32562
rect 2770 32510 2772 32562
rect 2268 31780 2324 31790
rect 2268 31686 2324 31724
rect 2716 31780 2772 32510
rect 2716 31714 2772 31724
rect 3388 32450 3444 32462
rect 3388 32398 3390 32450
rect 3442 32398 3444 32450
rect 2940 31668 2996 31678
rect 2828 31666 2996 31668
rect 2828 31614 2942 31666
rect 2994 31614 2996 31666
rect 2828 31612 2996 31614
rect 2828 28420 2884 31612
rect 2940 31602 2996 31612
rect 3388 30884 3444 32398
rect 5516 32452 5572 32462
rect 5964 32452 6020 32462
rect 6300 32452 6356 37102
rect 6524 36820 6580 40572
rect 9772 40402 9828 40414
rect 9772 40350 9774 40402
rect 9826 40350 9828 40402
rect 6860 40292 6916 40302
rect 6860 40290 8036 40292
rect 6860 40238 6862 40290
rect 6914 40238 8036 40290
rect 6860 40236 8036 40238
rect 6860 40226 6916 40236
rect 7980 39506 8036 40236
rect 8988 40290 9044 40302
rect 8988 40238 8990 40290
rect 9042 40238 9044 40290
rect 8988 40068 9044 40238
rect 8988 40002 9044 40012
rect 7980 39454 7982 39506
rect 8034 39454 8036 39506
rect 7980 39442 8036 39454
rect 8316 39508 8372 39518
rect 8316 39414 8372 39452
rect 7196 39284 7252 39294
rect 7196 38162 7252 39228
rect 7196 38110 7198 38162
rect 7250 38110 7252 38162
rect 7196 38098 7252 38110
rect 9324 38164 9380 38174
rect 9324 38162 9716 38164
rect 9324 38110 9326 38162
rect 9378 38110 9716 38162
rect 9324 38108 9716 38110
rect 9324 38098 9380 38108
rect 9660 37604 9716 38108
rect 9772 37828 9828 40350
rect 9996 40404 10052 42030
rect 13244 41860 13300 45200
rect 17052 45108 17108 45200
rect 17388 45108 17444 45276
rect 17052 45052 17444 45108
rect 17836 43708 17892 45276
rect 20832 45200 20944 46000
rect 21196 45276 21700 45332
rect 20860 45108 20916 45200
rect 21196 45108 21252 45276
rect 20860 45052 21252 45108
rect 17836 43652 18340 43708
rect 18284 42194 18340 43652
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 18284 42142 18286 42194
rect 18338 42142 18340 42194
rect 18284 42130 18340 42142
rect 13244 41794 13300 41804
rect 13468 41970 13524 41982
rect 13468 41918 13470 41970
rect 13522 41918 13524 41970
rect 11564 40516 11620 40526
rect 11452 40460 11564 40516
rect 11340 40404 11396 40414
rect 9996 40348 10612 40404
rect 9772 37734 9828 37772
rect 10332 38836 10388 38846
rect 9660 37548 9940 37604
rect 9884 37378 9940 37548
rect 9884 37326 9886 37378
rect 9938 37326 9940 37378
rect 9884 37314 9940 37326
rect 10332 37380 10388 38780
rect 10332 37286 10388 37324
rect 6524 36754 6580 36764
rect 9996 37042 10052 37054
rect 9996 36990 9998 37042
rect 10050 36990 10052 37042
rect 6972 36596 7028 36606
rect 6972 36502 7028 36540
rect 9996 36596 10052 36990
rect 9996 36530 10052 36540
rect 7084 36260 7140 36270
rect 7084 36166 7140 36204
rect 10220 36260 10276 36270
rect 10220 35810 10276 36204
rect 10220 35758 10222 35810
rect 10274 35758 10276 35810
rect 10220 35746 10276 35758
rect 10444 35476 10500 35486
rect 10332 35474 10500 35476
rect 10332 35422 10446 35474
rect 10498 35422 10500 35474
rect 10332 35420 10500 35422
rect 10332 35364 10388 35420
rect 10444 35410 10500 35420
rect 6636 33460 6692 33470
rect 6636 33366 6692 33404
rect 8988 33460 9044 33470
rect 8764 33236 8820 33246
rect 8316 33234 8820 33236
rect 8316 33182 8766 33234
rect 8818 33182 8820 33234
rect 8316 33180 8820 33182
rect 8316 32786 8372 33180
rect 8764 33170 8820 33180
rect 8316 32734 8318 32786
rect 8370 32734 8372 32786
rect 8316 32722 8372 32734
rect 8988 32788 9044 33404
rect 9548 33346 9604 33358
rect 9548 33294 9550 33346
rect 9602 33294 9604 33346
rect 9548 33124 9604 33294
rect 10332 33346 10388 35308
rect 10332 33294 10334 33346
rect 10386 33294 10388 33346
rect 10332 33282 10388 33294
rect 10556 33348 10612 40348
rect 11340 40310 11396 40348
rect 11452 39956 11508 40460
rect 11564 40422 11620 40460
rect 12012 40516 12068 40526
rect 11676 40404 11732 40414
rect 11676 40310 11732 40348
rect 11228 39900 11508 39956
rect 11228 39730 11284 39900
rect 11228 39678 11230 39730
rect 11282 39678 11284 39730
rect 11228 39666 11284 39678
rect 12012 39730 12068 40460
rect 12124 40514 12180 40526
rect 12124 40462 12126 40514
rect 12178 40462 12180 40514
rect 12124 40404 12180 40462
rect 12348 40516 12404 40526
rect 12348 40422 12404 40460
rect 12124 40338 12180 40348
rect 12572 40402 12628 40414
rect 12572 40350 12574 40402
rect 12626 40350 12628 40402
rect 12460 40292 12516 40302
rect 12460 40198 12516 40236
rect 12012 39678 12014 39730
rect 12066 39678 12068 39730
rect 12012 39666 12068 39678
rect 11004 39620 11060 39630
rect 11004 39526 11060 39564
rect 12572 39620 12628 40350
rect 13468 40180 13524 41918
rect 17276 41970 17332 41982
rect 21084 41972 21140 41982
rect 17276 41918 17278 41970
rect 17330 41918 17332 41970
rect 14476 41860 14532 41870
rect 14476 41766 14532 41804
rect 15708 40628 15764 40638
rect 16716 40628 16772 40638
rect 15708 40626 16772 40628
rect 15708 40574 15710 40626
rect 15762 40574 16718 40626
rect 16770 40574 16772 40626
rect 15708 40572 16772 40574
rect 15708 40562 15764 40572
rect 16716 40562 16772 40572
rect 14700 40514 14756 40526
rect 14700 40462 14702 40514
rect 14754 40462 14756 40514
rect 13468 40114 13524 40124
rect 13916 40404 13972 40414
rect 12572 39554 12628 39564
rect 12684 39508 12740 39518
rect 10668 39396 10724 39406
rect 10668 39302 10724 39340
rect 11676 39394 11732 39406
rect 11676 39342 11678 39394
rect 11730 39342 11732 39394
rect 11676 38948 11732 39342
rect 11900 39394 11956 39406
rect 12124 39396 12180 39406
rect 11900 39342 11902 39394
rect 11954 39342 11956 39394
rect 11900 39284 11956 39342
rect 11900 39218 11956 39228
rect 12012 39394 12180 39396
rect 12012 39342 12126 39394
rect 12178 39342 12180 39394
rect 12012 39340 12180 39342
rect 11676 38882 11732 38892
rect 12012 39060 12068 39340
rect 12124 39330 12180 39340
rect 12012 38050 12068 39004
rect 12572 38948 12628 38958
rect 12572 38854 12628 38892
rect 12684 38946 12740 39452
rect 13916 39058 13972 40348
rect 14364 40402 14420 40414
rect 14364 40350 14366 40402
rect 14418 40350 14420 40402
rect 14252 39620 14308 39630
rect 14028 39508 14084 39518
rect 14028 39414 14084 39452
rect 13916 39006 13918 39058
rect 13970 39006 13972 39058
rect 13916 38994 13972 39006
rect 12684 38894 12686 38946
rect 12738 38894 12740 38946
rect 12684 38882 12740 38894
rect 13804 38836 13860 38846
rect 13804 38742 13860 38780
rect 14028 38836 14084 38846
rect 14028 38668 14084 38780
rect 14028 38612 14196 38668
rect 12012 37998 12014 38050
rect 12066 37998 12068 38050
rect 12012 37986 12068 37998
rect 11676 37938 11732 37950
rect 11676 37886 11678 37938
rect 11730 37886 11732 37938
rect 10668 37492 10724 37502
rect 11116 37492 11172 37502
rect 10668 37490 11172 37492
rect 10668 37438 10670 37490
rect 10722 37438 11118 37490
rect 11170 37438 11172 37490
rect 10668 37436 11172 37438
rect 10668 37426 10724 37436
rect 11116 37426 11172 37436
rect 11004 37266 11060 37278
rect 11004 37214 11006 37266
rect 11058 37214 11060 37266
rect 11004 37044 11060 37214
rect 11004 36978 11060 36988
rect 11228 37268 11284 37278
rect 10780 35924 10836 35934
rect 11228 35924 11284 37212
rect 11564 37266 11620 37278
rect 11564 37214 11566 37266
rect 11618 37214 11620 37266
rect 11564 37156 11620 37214
rect 11564 37090 11620 37100
rect 11676 37044 11732 37886
rect 11788 37826 11844 37838
rect 11788 37774 11790 37826
rect 11842 37774 11844 37826
rect 11788 37268 11844 37774
rect 12460 37826 12516 37838
rect 12460 37774 12462 37826
rect 12514 37774 12516 37826
rect 11788 37202 11844 37212
rect 12236 37378 12292 37390
rect 12236 37326 12238 37378
rect 12290 37326 12292 37378
rect 12236 37268 12292 37326
rect 12236 37202 12292 37212
rect 12348 37266 12404 37278
rect 12348 37214 12350 37266
rect 12402 37214 12404 37266
rect 11676 36978 11732 36988
rect 12348 37044 12404 37214
rect 12460 37156 12516 37774
rect 12460 37090 12516 37100
rect 12348 36978 12404 36988
rect 12012 36820 12068 36830
rect 12012 36594 12068 36764
rect 13468 36820 13524 36830
rect 12012 36542 12014 36594
rect 12066 36542 12068 36594
rect 12012 36530 12068 36542
rect 12348 36596 12404 36606
rect 12348 36502 12404 36540
rect 12908 36596 12964 36606
rect 12908 36502 12964 36540
rect 12572 36484 12628 36494
rect 12572 36390 12628 36428
rect 13244 36484 13300 36494
rect 10780 35922 11284 35924
rect 10780 35870 10782 35922
rect 10834 35870 11284 35922
rect 10780 35868 11284 35870
rect 10780 35858 10836 35868
rect 13020 35812 13076 35822
rect 13020 35718 13076 35756
rect 13244 35700 13300 36428
rect 13468 36484 13524 36764
rect 14140 36708 14196 38612
rect 14252 37378 14308 39564
rect 14364 39508 14420 40350
rect 14700 40180 14756 40462
rect 15484 40514 15540 40526
rect 15484 40462 15486 40514
rect 15538 40462 15540 40514
rect 14364 39442 14420 39452
rect 14476 40124 14700 40180
rect 14476 38834 14532 40124
rect 14700 40114 14756 40124
rect 15372 40402 15428 40414
rect 15372 40350 15374 40402
rect 15426 40350 15428 40402
rect 15372 39956 15428 40350
rect 15148 39900 15428 39956
rect 15484 40180 15540 40462
rect 16940 40516 16996 40526
rect 16940 40422 16996 40460
rect 14924 39620 14980 39630
rect 15148 39620 15204 39900
rect 14924 39618 15204 39620
rect 14924 39566 14926 39618
rect 14978 39566 15204 39618
rect 14924 39564 15204 39566
rect 15260 39620 15316 39630
rect 15484 39620 15540 40124
rect 16604 40402 16660 40414
rect 16604 40350 16606 40402
rect 16658 40350 16660 40402
rect 16044 39732 16100 39742
rect 16044 39638 16100 39676
rect 15260 39618 15540 39620
rect 15260 39566 15262 39618
rect 15314 39566 15540 39618
rect 15260 39564 15540 39566
rect 15596 39620 15652 39630
rect 14812 39508 14868 39518
rect 14588 39396 14644 39406
rect 14588 39302 14644 39340
rect 14476 38782 14478 38834
rect 14530 38782 14532 38834
rect 14476 38770 14532 38782
rect 14252 37326 14254 37378
rect 14306 37326 14308 37378
rect 14252 37314 14308 37326
rect 14476 37266 14532 37278
rect 14476 37214 14478 37266
rect 14530 37214 14532 37266
rect 14476 37156 14532 37214
rect 14476 37090 14532 37100
rect 14588 37044 14644 37054
rect 14252 36708 14308 36718
rect 14140 36706 14308 36708
rect 14140 36654 14254 36706
rect 14306 36654 14308 36706
rect 14140 36652 14308 36654
rect 14252 36642 14308 36652
rect 13468 36390 13524 36428
rect 13804 36596 13860 36606
rect 13804 36482 13860 36540
rect 14476 36484 14532 36494
rect 13804 36430 13806 36482
rect 13858 36430 13860 36482
rect 13804 36418 13860 36430
rect 13916 36482 14532 36484
rect 13916 36430 14478 36482
rect 14530 36430 14532 36482
rect 13916 36428 14532 36430
rect 13692 36372 13748 36382
rect 13692 36278 13748 36316
rect 13916 36036 13972 36428
rect 14476 36418 14532 36428
rect 13580 35980 13972 36036
rect 13580 35922 13636 35980
rect 13580 35870 13582 35922
rect 13634 35870 13636 35922
rect 13580 35858 13636 35870
rect 14588 35922 14644 36988
rect 14812 36594 14868 39452
rect 14924 38948 14980 39564
rect 15260 39554 15316 39564
rect 15148 39284 15204 39294
rect 15148 39058 15204 39228
rect 15148 39006 15150 39058
rect 15202 39006 15204 39058
rect 15148 38994 15204 39006
rect 15372 38948 15428 39564
rect 15596 39526 15652 39564
rect 15820 39508 15876 39518
rect 15484 39396 15540 39406
rect 15484 39394 15652 39396
rect 15484 39342 15486 39394
rect 15538 39342 15652 39394
rect 15484 39340 15652 39342
rect 15484 39330 15540 39340
rect 15484 38948 15540 38958
rect 15372 38946 15540 38948
rect 15372 38894 15486 38946
rect 15538 38894 15540 38946
rect 15372 38892 15540 38894
rect 14924 38882 14980 38892
rect 15484 38882 15540 38892
rect 15036 38836 15092 38846
rect 15036 38742 15092 38780
rect 15596 38836 15652 39340
rect 15708 39060 15764 39070
rect 15708 38966 15764 39004
rect 15596 38770 15652 38780
rect 15820 38722 15876 39452
rect 15932 39394 15988 39406
rect 15932 39342 15934 39394
rect 15986 39342 15988 39394
rect 15932 39060 15988 39342
rect 16156 39394 16212 39406
rect 16156 39342 16158 39394
rect 16210 39342 16212 39394
rect 16156 39284 16212 39342
rect 16380 39396 16436 39406
rect 16604 39396 16660 40350
rect 17276 40068 17332 41918
rect 20748 41970 21140 41972
rect 20748 41918 21086 41970
rect 21138 41918 21140 41970
rect 20748 41916 21140 41918
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 17276 40002 17332 40012
rect 17836 40404 17892 40414
rect 17836 39618 17892 40348
rect 20076 40404 20132 40414
rect 20300 40404 20356 40414
rect 20132 40402 20356 40404
rect 20132 40350 20302 40402
rect 20354 40350 20356 40402
rect 20132 40348 20356 40350
rect 20076 40310 20132 40348
rect 20300 40338 20356 40348
rect 20748 39730 20804 41916
rect 21084 41906 21140 41916
rect 21644 41860 21700 45276
rect 24640 45200 24752 46000
rect 28448 45200 28560 46000
rect 32256 45200 32368 46000
rect 32620 45276 33124 45332
rect 23212 41972 23268 41982
rect 22092 41860 22148 41870
rect 21644 41858 22148 41860
rect 21644 41806 22094 41858
rect 22146 41806 22148 41858
rect 21644 41804 22148 41806
rect 22092 41794 22148 41804
rect 21420 40404 21476 40414
rect 21084 40292 21140 40302
rect 21084 40198 21140 40236
rect 20748 39678 20750 39730
rect 20802 39678 20804 39730
rect 20748 39666 20804 39678
rect 21420 39730 21476 40348
rect 23212 40290 23268 41916
rect 24668 41860 24724 45200
rect 28476 42196 28532 45200
rect 32284 45108 32340 45200
rect 32620 45108 32676 45276
rect 32284 45052 32676 45108
rect 33068 43708 33124 45276
rect 36064 45200 36176 46000
rect 39872 45200 39984 46000
rect 43680 45200 43792 46000
rect 33068 43652 33572 43708
rect 28476 42130 28532 42140
rect 33516 42194 33572 43652
rect 33516 42142 33518 42194
rect 33570 42142 33572 42194
rect 33516 42130 33572 42142
rect 24892 41972 24948 41982
rect 28700 41972 28756 41982
rect 24892 41878 24948 41916
rect 28140 41970 28756 41972
rect 28140 41918 28702 41970
rect 28754 41918 28756 41970
rect 28140 41916 28756 41918
rect 24668 41794 24724 41804
rect 25900 41860 25956 41870
rect 25900 41766 25956 41804
rect 25340 40404 25396 40414
rect 25340 40310 25396 40348
rect 23212 40238 23214 40290
rect 23266 40238 23268 40290
rect 23212 40226 23268 40238
rect 26012 40290 26068 40302
rect 26012 40238 26014 40290
rect 26066 40238 26068 40290
rect 21420 39678 21422 39730
rect 21474 39678 21476 39730
rect 21420 39666 21476 39678
rect 17836 39566 17838 39618
rect 17890 39566 17892 39618
rect 16828 39508 16884 39518
rect 16828 39414 16884 39452
rect 16436 39340 16660 39396
rect 16940 39396 16996 39406
rect 16380 39302 16436 39340
rect 16940 39302 16996 39340
rect 17052 39394 17108 39406
rect 17052 39342 17054 39394
rect 17106 39342 17108 39394
rect 16156 39218 16212 39228
rect 17052 39284 17108 39342
rect 17052 39218 17108 39228
rect 15932 38994 15988 39004
rect 15820 38670 15822 38722
rect 15874 38670 15876 38722
rect 15820 38658 15876 38670
rect 17836 38500 17892 39566
rect 18620 39620 18676 39630
rect 18620 39526 18676 39564
rect 26012 39396 26068 40238
rect 28140 40290 28196 41916
rect 28700 41906 28756 41916
rect 30380 41972 30436 41982
rect 30380 41878 30436 41916
rect 31388 41972 31444 41982
rect 28140 40238 28142 40290
rect 28194 40238 28196 40290
rect 28140 40226 28196 40238
rect 28588 40404 28644 40414
rect 26012 39330 26068 39340
rect 28364 39620 28420 39630
rect 28588 39620 28644 40348
rect 29260 40290 29316 40302
rect 29260 40238 29262 40290
rect 29314 40238 29316 40290
rect 29260 39732 29316 40238
rect 31388 40290 31444 41916
rect 32508 41972 32564 41982
rect 32508 41878 32564 41916
rect 33740 41972 33796 41982
rect 31388 40238 31390 40290
rect 31442 40238 31444 40290
rect 31388 40226 31444 40238
rect 31612 40516 31668 40526
rect 29260 39666 29316 39676
rect 31612 39730 31668 40460
rect 31612 39678 31614 39730
rect 31666 39678 31668 39730
rect 31612 39666 31668 39678
rect 31948 40402 32004 40414
rect 31948 40350 31950 40402
rect 32002 40350 32004 40402
rect 28420 39564 28644 39620
rect 30268 39620 30324 39630
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 16828 38444 17892 38500
rect 16268 37378 16324 37390
rect 16268 37326 16270 37378
rect 16322 37326 16324 37378
rect 14812 36542 14814 36594
rect 14866 36542 14868 36594
rect 14812 36530 14868 36542
rect 15596 37266 15652 37278
rect 15596 37214 15598 37266
rect 15650 37214 15652 37266
rect 15596 36596 15652 37214
rect 15596 36530 15652 36540
rect 15036 36484 15092 36494
rect 15036 36370 15092 36428
rect 15484 36484 15540 36494
rect 15484 36390 15540 36428
rect 15036 36318 15038 36370
rect 15090 36318 15092 36370
rect 15036 36306 15092 36318
rect 16268 36372 16324 37326
rect 16716 37156 16772 37166
rect 16716 37062 16772 37100
rect 16268 36306 16324 36316
rect 14588 35870 14590 35922
rect 14642 35870 14644 35922
rect 14588 35858 14644 35870
rect 14812 36258 14868 36270
rect 14812 36206 14814 36258
rect 14866 36206 14868 36258
rect 14700 35810 14756 35822
rect 14700 35758 14702 35810
rect 14754 35758 14756 35810
rect 13244 35606 13300 35644
rect 13916 35700 13972 35710
rect 13916 34354 13972 35644
rect 14588 35698 14644 35710
rect 14588 35646 14590 35698
rect 14642 35646 14644 35698
rect 13916 34302 13918 34354
rect 13970 34302 13972 34354
rect 13916 34290 13972 34302
rect 14252 35364 14308 35374
rect 14252 34692 14308 35308
rect 14588 35028 14644 35646
rect 14700 35364 14756 35758
rect 14700 35298 14756 35308
rect 14588 34972 14756 35028
rect 14700 34804 14756 34972
rect 14812 35026 14868 36206
rect 15484 35812 15540 35822
rect 15484 35810 16660 35812
rect 15484 35758 15486 35810
rect 15538 35758 16660 35810
rect 15484 35756 16660 35758
rect 15484 35746 15540 35756
rect 14812 34974 14814 35026
rect 14866 34974 14868 35026
rect 14812 34962 14868 34974
rect 15036 35588 15092 35598
rect 15036 34914 15092 35532
rect 16604 35138 16660 35756
rect 16604 35086 16606 35138
rect 16658 35086 16660 35138
rect 16604 35074 16660 35086
rect 16716 35476 16772 35486
rect 16716 35026 16772 35420
rect 16716 34974 16718 35026
rect 16770 34974 16772 35026
rect 16716 34962 16772 34974
rect 15036 34862 15038 34914
rect 15090 34862 15092 34914
rect 15036 34850 15092 34862
rect 14812 34804 14868 34814
rect 14700 34748 14812 34804
rect 14812 34710 14868 34748
rect 14588 34692 14644 34702
rect 14252 34690 14644 34692
rect 14252 34638 14590 34690
rect 14642 34638 14644 34690
rect 14252 34636 14644 34638
rect 14252 34354 14308 34636
rect 14588 34626 14644 34636
rect 14252 34302 14254 34354
rect 14306 34302 14308 34354
rect 14252 34290 14308 34302
rect 10556 33292 10724 33348
rect 9996 33124 10052 33134
rect 9548 33122 10052 33124
rect 9548 33070 9998 33122
rect 10050 33070 10052 33122
rect 9548 33068 10052 33070
rect 8428 32676 8484 32686
rect 8428 32582 8484 32620
rect 8988 32674 9044 32732
rect 9772 32788 9828 32798
rect 9772 32694 9828 32732
rect 8988 32622 8990 32674
rect 9042 32622 9044 32674
rect 8988 32610 9044 32622
rect 5516 32450 5908 32452
rect 5516 32398 5518 32450
rect 5570 32398 5908 32450
rect 5516 32396 5908 32398
rect 5516 32386 5572 32396
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 5068 31892 5124 31902
rect 5068 31890 5684 31892
rect 5068 31838 5070 31890
rect 5122 31838 5684 31890
rect 5068 31836 5684 31838
rect 5068 31826 5124 31836
rect 3388 30818 3444 30828
rect 4956 30884 5012 30894
rect 5012 30828 5124 30884
rect 4956 30818 5012 30828
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 5068 29650 5124 30828
rect 5068 29598 5070 29650
rect 5122 29598 5124 29650
rect 5068 29586 5124 29598
rect 5628 29538 5684 31836
rect 5628 29486 5630 29538
rect 5682 29486 5684 29538
rect 3388 29428 3444 29438
rect 3276 28980 3332 28990
rect 3276 28866 3332 28924
rect 3276 28814 3278 28866
rect 3330 28814 3332 28866
rect 3276 28802 3332 28814
rect 3164 28644 3220 28654
rect 3164 28550 3220 28588
rect 2940 28420 2996 28430
rect 2828 28418 2996 28420
rect 2828 28366 2942 28418
rect 2994 28366 2996 28418
rect 2828 28364 2996 28366
rect 2940 28354 2996 28364
rect 3388 26908 3444 29372
rect 3724 29426 3780 29438
rect 3724 29374 3726 29426
rect 3778 29374 3780 29426
rect 3612 28644 3668 28654
rect 3500 28532 3556 28542
rect 3500 28438 3556 28476
rect 3612 28082 3668 28588
rect 3612 28030 3614 28082
rect 3666 28030 3668 28082
rect 3388 26852 3556 26908
rect 2940 25284 2996 25294
rect 2940 24050 2996 25228
rect 2940 23998 2942 24050
rect 2994 23998 2996 24050
rect 2940 23986 2996 23998
rect 3164 24500 3220 24510
rect 2268 23940 2324 23950
rect 2268 23846 2324 23884
rect 3164 23266 3220 24444
rect 3164 23214 3166 23266
rect 3218 23214 3220 23266
rect 3164 23202 3220 23214
rect 2492 23156 2548 23166
rect 2492 23062 2548 23100
rect 1820 22082 1876 22092
rect 1820 19234 1876 19246
rect 1820 19182 1822 19234
rect 1874 19182 1876 19234
rect 1820 18564 1876 19182
rect 1820 18498 1876 18508
rect 2604 19122 2660 19134
rect 2604 19070 2606 19122
rect 2658 19070 2660 19122
rect 2604 18452 2660 19070
rect 3500 18564 3556 26852
rect 3612 21924 3668 28030
rect 3724 28530 3780 29374
rect 3948 29428 4004 29438
rect 3948 29426 4340 29428
rect 3948 29374 3950 29426
rect 4002 29374 4340 29426
rect 3948 29372 4340 29374
rect 3948 29362 4004 29372
rect 3836 29314 3892 29326
rect 3836 29262 3838 29314
rect 3890 29262 3892 29314
rect 3836 28980 3892 29262
rect 3836 28914 3892 28924
rect 4284 28866 4340 29372
rect 4396 29426 4452 29438
rect 4396 29374 4398 29426
rect 4450 29374 4452 29426
rect 4396 29204 4452 29374
rect 4620 29428 4676 29438
rect 4620 29334 4676 29372
rect 4844 29426 4900 29438
rect 4844 29374 4846 29426
rect 4898 29374 4900 29426
rect 4396 29138 4452 29148
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4284 28814 4286 28866
rect 4338 28814 4340 28866
rect 3724 28478 3726 28530
rect 3778 28478 3780 28530
rect 3724 27860 3780 28478
rect 4060 28756 4116 28766
rect 4060 28530 4116 28700
rect 4060 28478 4062 28530
rect 4114 28478 4116 28530
rect 4060 28308 4116 28478
rect 4284 28532 4340 28814
rect 4284 28466 4340 28476
rect 4396 28868 4452 28878
rect 4396 28308 4452 28812
rect 4508 28644 4564 28654
rect 4508 28550 4564 28588
rect 4732 28644 4788 28654
rect 4732 28550 4788 28588
rect 4060 28252 4228 28308
rect 4172 27970 4228 28252
rect 4172 27918 4174 27970
rect 4226 27918 4228 27970
rect 4172 27906 4228 27918
rect 4284 28252 4452 28308
rect 4508 28420 4564 28430
rect 3724 27794 3780 27804
rect 4284 27858 4340 28252
rect 4508 28082 4564 28364
rect 4508 28030 4510 28082
rect 4562 28030 4564 28082
rect 4508 28018 4564 28030
rect 4620 28084 4676 28094
rect 4844 28084 4900 29374
rect 5180 29426 5236 29438
rect 5180 29374 5182 29426
rect 5234 29374 5236 29426
rect 5068 28980 5124 28990
rect 5068 28532 5124 28924
rect 5180 28866 5236 29374
rect 5628 29428 5684 29486
rect 5628 29362 5684 29372
rect 5740 31554 5796 31566
rect 5740 31502 5742 31554
rect 5794 31502 5796 31554
rect 5740 31108 5796 31502
rect 5180 28814 5182 28866
rect 5234 28814 5236 28866
rect 5180 28802 5236 28814
rect 5516 29202 5572 29214
rect 5516 29150 5518 29202
rect 5570 29150 5572 29202
rect 5068 28466 5124 28476
rect 4620 28082 4900 28084
rect 4620 28030 4622 28082
rect 4674 28030 4900 28082
rect 4620 28028 4900 28030
rect 4956 28420 5012 28430
rect 4956 28084 5012 28364
rect 5068 28084 5124 28094
rect 4956 28082 5124 28084
rect 4956 28030 5070 28082
rect 5122 28030 5124 28082
rect 4956 28028 5124 28030
rect 4620 28018 4676 28028
rect 5068 28018 5124 28028
rect 5404 27972 5460 27982
rect 5516 27972 5572 29150
rect 5628 28420 5684 28430
rect 5628 28326 5684 28364
rect 5180 27970 5572 27972
rect 5180 27918 5406 27970
rect 5458 27918 5572 27970
rect 5180 27916 5572 27918
rect 4284 27806 4286 27858
rect 4338 27806 4340 27858
rect 4284 27748 4340 27806
rect 4732 27860 4788 27870
rect 4732 27766 4788 27804
rect 4284 27682 4340 27692
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 5180 26964 5236 27916
rect 5404 27906 5460 27916
rect 5292 27748 5348 27758
rect 5348 27692 5572 27748
rect 5292 27682 5348 27692
rect 5180 26908 5348 26964
rect 5292 26852 5460 26908
rect 3836 26740 3892 26750
rect 3836 26402 3892 26684
rect 3836 26350 3838 26402
rect 3890 26350 3892 26402
rect 3836 26338 3892 26350
rect 3724 26066 3780 26078
rect 3724 26014 3726 26066
rect 3778 26014 3780 26066
rect 3724 24500 3780 26014
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 3724 24434 3780 24444
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 5068 24052 5124 24062
rect 5068 23958 5124 23996
rect 5292 23156 5348 23166
rect 5292 23042 5348 23100
rect 5292 22990 5294 23042
rect 5346 22990 5348 23042
rect 5292 22978 5348 22990
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 5404 22372 5460 26852
rect 5516 25506 5572 27692
rect 5740 27076 5796 31052
rect 5852 30212 5908 32396
rect 5964 32450 6356 32452
rect 5964 32398 5966 32450
rect 6018 32398 6356 32450
rect 5964 32396 6356 32398
rect 8092 32562 8148 32574
rect 8092 32510 8094 32562
rect 8146 32510 8148 32562
rect 5964 31780 6020 32396
rect 5964 31108 6020 31724
rect 5964 31042 6020 31052
rect 5852 30146 5908 30156
rect 6636 30436 6692 30446
rect 6076 29316 6132 29326
rect 6076 29222 6132 29260
rect 6300 28980 6356 28990
rect 5964 28644 6020 28654
rect 5964 28550 6020 28588
rect 6300 28532 6356 28924
rect 6412 28868 6468 28878
rect 6412 28774 6468 28812
rect 6412 28532 6468 28542
rect 6300 28530 6468 28532
rect 6300 28478 6414 28530
rect 6466 28478 6468 28530
rect 6300 28476 6468 28478
rect 6412 28466 6468 28476
rect 6524 28532 6580 28542
rect 6524 28438 6580 28476
rect 5964 28420 6020 28430
rect 5964 27860 6020 28364
rect 5740 27020 5908 27076
rect 5516 25454 5518 25506
rect 5570 25454 5572 25506
rect 5516 25442 5572 25454
rect 5740 25284 5796 25294
rect 5740 25190 5796 25228
rect 5852 23940 5908 27020
rect 5964 26290 6020 27804
rect 6636 26514 6692 30380
rect 8092 30436 8148 32510
rect 8876 32338 8932 32350
rect 8876 32286 8878 32338
rect 8930 32286 8932 32338
rect 8092 30370 8148 30380
rect 8764 30436 8820 30446
rect 8764 30342 8820 30380
rect 8764 30212 8820 30222
rect 8876 30212 8932 32286
rect 9996 31892 10052 33068
rect 10444 33122 10500 33134
rect 10444 33070 10446 33122
rect 10498 33070 10500 33122
rect 10444 32676 10500 33070
rect 10444 32610 10500 32620
rect 10556 33122 10612 33134
rect 10556 33070 10558 33122
rect 10610 33070 10612 33122
rect 9996 31826 10052 31836
rect 10332 32452 10388 32462
rect 10556 32452 10612 33070
rect 10332 32450 10612 32452
rect 10332 32398 10334 32450
rect 10386 32398 10612 32450
rect 10332 32396 10612 32398
rect 9100 30324 9156 30334
rect 9100 30230 9156 30268
rect 9660 30212 9716 30222
rect 8540 30210 8932 30212
rect 8540 30158 8766 30210
rect 8818 30158 8932 30210
rect 8540 30156 8932 30158
rect 9436 30210 9716 30212
rect 9436 30158 9662 30210
rect 9714 30158 9716 30210
rect 9436 30156 9716 30158
rect 6972 29652 7028 29662
rect 6972 28754 7028 29596
rect 6972 28702 6974 28754
rect 7026 28702 7028 28754
rect 6972 28532 7028 28702
rect 7980 28644 8036 28654
rect 7980 28550 8036 28588
rect 6972 28466 7028 28476
rect 8316 28532 8372 28542
rect 7868 28420 7924 28430
rect 8204 28420 8260 28430
rect 7868 28418 8260 28420
rect 7868 28366 7870 28418
rect 7922 28366 8206 28418
rect 8258 28366 8260 28418
rect 7868 28364 8260 28366
rect 7868 28354 7924 28364
rect 8204 28084 8260 28364
rect 8204 28018 8260 28028
rect 6636 26462 6638 26514
rect 6690 26462 6692 26514
rect 6636 26450 6692 26462
rect 5964 26238 5966 26290
rect 6018 26238 6020 26290
rect 5964 26226 6020 26238
rect 6412 26404 6468 26414
rect 6300 25732 6356 25742
rect 5964 25730 6356 25732
rect 5964 25678 6302 25730
rect 6354 25678 6356 25730
rect 5964 25676 6356 25678
rect 5964 25506 6020 25676
rect 6300 25666 6356 25676
rect 5964 25454 5966 25506
rect 6018 25454 6020 25506
rect 5964 25442 6020 25454
rect 6188 25394 6244 25406
rect 6188 25342 6190 25394
rect 6242 25342 6244 25394
rect 6188 25284 6244 25342
rect 6188 25218 6244 25228
rect 6412 24050 6468 26348
rect 6524 26178 6580 26190
rect 6524 26126 6526 26178
rect 6578 26126 6580 26178
rect 6524 25730 6580 26126
rect 6524 25678 6526 25730
rect 6578 25678 6580 25730
rect 6524 25666 6580 25678
rect 8316 25620 8372 28476
rect 8540 25732 8596 30156
rect 8764 30146 8820 30156
rect 8652 29540 8708 29550
rect 8652 29538 8932 29540
rect 8652 29486 8654 29538
rect 8706 29486 8932 29538
rect 8652 29484 8932 29486
rect 8652 29474 8708 29484
rect 8876 28756 8932 29484
rect 8764 28644 8820 28654
rect 8764 28550 8820 28588
rect 8876 28642 8932 28700
rect 8876 28590 8878 28642
rect 8930 28590 8932 28642
rect 8876 28578 8932 28590
rect 8988 29428 9044 29438
rect 9436 29428 9492 30156
rect 9660 30146 9716 30156
rect 10108 30212 10164 30222
rect 10108 30118 10164 30156
rect 8988 29426 9492 29428
rect 8988 29374 8990 29426
rect 9042 29374 9492 29426
rect 8988 29372 9492 29374
rect 9996 29428 10052 29466
rect 8988 26628 9044 29372
rect 9996 29362 10052 29372
rect 9660 29316 9716 29326
rect 9100 29314 9828 29316
rect 9100 29262 9662 29314
rect 9714 29262 9828 29314
rect 9100 29260 9828 29262
rect 9100 28530 9156 29260
rect 9660 29250 9716 29260
rect 9660 28868 9716 28878
rect 9660 28774 9716 28812
rect 9548 28756 9604 28766
rect 9100 28478 9102 28530
rect 9154 28478 9156 28530
rect 9100 28466 9156 28478
rect 9212 28642 9268 28654
rect 9212 28590 9214 28642
rect 9266 28590 9268 28642
rect 9212 28532 9268 28590
rect 9212 28466 9268 28476
rect 9548 27858 9604 28700
rect 9548 27806 9550 27858
rect 9602 27806 9604 27858
rect 9548 27794 9604 27806
rect 9772 27858 9828 29260
rect 9884 29204 9940 29214
rect 9884 28644 9940 29148
rect 9884 28550 9940 28588
rect 10108 28532 10164 28542
rect 9996 28084 10052 28094
rect 9996 27970 10052 28028
rect 9996 27918 9998 27970
rect 10050 27918 10052 27970
rect 9996 27906 10052 27918
rect 9772 27806 9774 27858
rect 9826 27806 9828 27858
rect 8988 26562 9044 26572
rect 9772 26292 9828 27806
rect 10108 27858 10164 28476
rect 10108 27806 10110 27858
rect 10162 27806 10164 27858
rect 10108 27794 10164 27806
rect 10332 26516 10388 32396
rect 10444 31108 10500 31118
rect 10444 31014 10500 31052
rect 10668 30212 10724 33292
rect 11004 33346 11060 33358
rect 11004 33294 11006 33346
rect 11058 33294 11060 33346
rect 11004 33124 11060 33294
rect 11452 33124 11508 33134
rect 11004 33122 11508 33124
rect 11004 33070 11454 33122
rect 11506 33070 11508 33122
rect 11004 33068 11508 33070
rect 10556 30210 10724 30212
rect 10556 30158 10670 30210
rect 10722 30158 10724 30210
rect 10556 30156 10724 30158
rect 10556 29428 10612 30156
rect 10668 30146 10724 30156
rect 10780 29538 10836 29550
rect 10780 29486 10782 29538
rect 10834 29486 10836 29538
rect 10556 29426 10724 29428
rect 10556 29374 10558 29426
rect 10610 29374 10724 29426
rect 10556 29372 10724 29374
rect 10556 29362 10612 29372
rect 10444 28644 10500 28654
rect 10444 28642 10612 28644
rect 10444 28590 10446 28642
rect 10498 28590 10612 28642
rect 10444 28588 10612 28590
rect 10444 28578 10500 28588
rect 10556 28082 10612 28588
rect 10556 28030 10558 28082
rect 10610 28030 10612 28082
rect 10556 28018 10612 28030
rect 10668 27188 10724 29372
rect 10780 28980 10836 29486
rect 10780 28914 10836 28924
rect 10892 28756 10948 28766
rect 10668 27122 10724 27132
rect 10780 28530 10836 28542
rect 10780 28478 10782 28530
rect 10834 28478 10836 28530
rect 10780 26740 10836 28478
rect 10892 28084 10948 28700
rect 11228 28644 11284 28654
rect 11340 28644 11396 33068
rect 11452 33058 11508 33068
rect 13468 31890 13524 31902
rect 13468 31838 13470 31890
rect 13522 31838 13524 31890
rect 12012 30324 12068 30334
rect 11900 30212 11956 30222
rect 11452 29428 11508 29438
rect 11452 29334 11508 29372
rect 11900 29426 11956 30156
rect 11900 29374 11902 29426
rect 11954 29374 11956 29426
rect 11900 29362 11956 29374
rect 11284 28588 11396 28644
rect 11564 29316 11620 29326
rect 11564 28642 11620 29260
rect 11676 29204 11732 29214
rect 11676 29110 11732 29148
rect 11564 28590 11566 28642
rect 11618 28590 11620 28642
rect 11228 28550 11284 28588
rect 11564 28578 11620 28590
rect 12012 28532 12068 30268
rect 13468 30212 13524 31838
rect 16380 31892 16436 31902
rect 16380 31778 16436 31836
rect 16380 31726 16382 31778
rect 16434 31726 16436 31778
rect 16380 31714 16436 31726
rect 16828 31892 16884 38444
rect 22764 38164 22820 38174
rect 25564 38164 25620 38174
rect 22764 38050 22820 38108
rect 22764 37998 22766 38050
rect 22818 37998 22820 38050
rect 22764 37986 22820 37998
rect 25452 38162 25620 38164
rect 25452 38110 25566 38162
rect 25618 38110 25620 38162
rect 25452 38108 25620 38110
rect 23436 37938 23492 37950
rect 23436 37886 23438 37938
rect 23490 37886 23492 37938
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19628 37154 19684 37166
rect 19628 37102 19630 37154
rect 19682 37102 19684 37154
rect 18396 36484 18452 36494
rect 18396 36390 18452 36428
rect 19068 36484 19124 36494
rect 19068 36390 19124 36428
rect 19292 36482 19348 36494
rect 19292 36430 19294 36482
rect 19346 36430 19348 36482
rect 17724 36372 17780 36382
rect 17724 35810 17780 36316
rect 17724 35758 17726 35810
rect 17778 35758 17780 35810
rect 17724 35746 17780 35758
rect 18060 36258 18116 36270
rect 18060 36206 18062 36258
rect 18114 36206 18116 36258
rect 17276 35700 17332 35710
rect 17276 31948 17332 35644
rect 18060 35588 18116 36206
rect 18284 36260 18340 36270
rect 18732 36260 18788 36270
rect 18284 36258 18452 36260
rect 18284 36206 18286 36258
rect 18338 36206 18452 36258
rect 18284 36204 18452 36206
rect 18284 36194 18340 36204
rect 18060 35522 18116 35532
rect 18172 35698 18228 35710
rect 18172 35646 18174 35698
rect 18226 35646 18228 35698
rect 18172 35140 18228 35646
rect 18396 35700 18452 36204
rect 18732 36258 18900 36260
rect 18732 36206 18734 36258
rect 18786 36206 18900 36258
rect 18732 36204 18900 36206
rect 18732 36194 18788 36204
rect 18284 35140 18340 35150
rect 18172 35138 18340 35140
rect 18172 35086 18286 35138
rect 18338 35086 18340 35138
rect 18172 35084 18340 35086
rect 18284 35074 18340 35084
rect 18396 34804 18452 35644
rect 18844 35476 18900 36204
rect 19292 35924 19348 36430
rect 19628 36372 19684 37102
rect 20300 37156 20356 37166
rect 19628 36306 19684 36316
rect 19964 36372 20020 36382
rect 19964 36278 20020 36316
rect 20300 36372 20356 37100
rect 20972 36484 21028 36494
rect 20748 36372 20804 36382
rect 20300 36370 20468 36372
rect 20300 36318 20302 36370
rect 20354 36318 20468 36370
rect 20300 36316 20468 36318
rect 20300 36306 20356 36316
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 18844 35382 18900 35420
rect 19068 35868 19348 35924
rect 18620 35140 18676 35150
rect 18620 35046 18676 35084
rect 18396 34710 18452 34748
rect 18956 34692 19012 34702
rect 18956 34598 19012 34636
rect 19068 34354 19124 35868
rect 20300 35812 20356 35822
rect 19180 35700 19236 35710
rect 19516 35700 19572 35710
rect 19964 35700 20020 35710
rect 19180 35698 19572 35700
rect 19180 35646 19182 35698
rect 19234 35646 19518 35698
rect 19570 35646 19572 35698
rect 19180 35644 19572 35646
rect 19180 35634 19236 35644
rect 19516 35634 19572 35644
rect 19852 35698 20020 35700
rect 19852 35646 19966 35698
rect 20018 35646 20020 35698
rect 19852 35644 20020 35646
rect 19068 34302 19070 34354
rect 19122 34302 19124 34354
rect 19068 34290 19124 34302
rect 19180 35140 19236 35150
rect 19180 34356 19236 35084
rect 19852 35140 19908 35644
rect 19964 35634 20020 35644
rect 20076 35700 20132 35710
rect 20076 35606 20132 35644
rect 20300 35698 20356 35756
rect 20300 35646 20302 35698
rect 20354 35646 20356 35698
rect 20300 35308 20356 35646
rect 19852 35074 19908 35084
rect 19964 35252 20356 35308
rect 19292 35028 19348 35038
rect 19292 35026 19684 35028
rect 19292 34974 19294 35026
rect 19346 34974 19684 35026
rect 19292 34972 19684 34974
rect 19292 34962 19348 34972
rect 19628 34916 19684 34972
rect 19740 34916 19796 34926
rect 19628 34914 19796 34916
rect 19628 34862 19742 34914
rect 19794 34862 19796 34914
rect 19628 34860 19796 34862
rect 19740 34850 19796 34860
rect 19516 34804 19572 34814
rect 19516 34710 19572 34748
rect 19964 34802 20020 35252
rect 19964 34750 19966 34802
rect 20018 34750 20020 34802
rect 19964 34738 20020 34750
rect 20076 34802 20132 34814
rect 20076 34750 20078 34802
rect 20130 34750 20132 34802
rect 20076 34692 20132 34750
rect 20076 34636 20244 34692
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19180 34242 19236 34300
rect 20076 34356 20132 34366
rect 20188 34356 20244 34636
rect 20132 34300 20244 34356
rect 20076 34290 20132 34300
rect 19180 34190 19182 34242
rect 19234 34190 19236 34242
rect 19180 34178 19236 34190
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 15596 31668 15652 31678
rect 15596 31666 15876 31668
rect 15596 31614 15598 31666
rect 15650 31614 15876 31666
rect 15596 31612 15876 31614
rect 15596 31602 15652 31612
rect 15820 31218 15876 31612
rect 15820 31166 15822 31218
rect 15874 31166 15876 31218
rect 15820 31154 15876 31166
rect 15484 30996 15540 31006
rect 15484 30902 15540 30940
rect 16492 30996 16548 31006
rect 15932 30882 15988 30894
rect 15932 30830 15934 30882
rect 15986 30830 15988 30882
rect 13580 30212 13636 30222
rect 13468 30210 13636 30212
rect 13468 30158 13582 30210
rect 13634 30158 13636 30210
rect 13468 30156 13636 30158
rect 12124 29540 12180 29550
rect 12124 29426 12180 29484
rect 12124 29374 12126 29426
rect 12178 29374 12180 29426
rect 12124 29362 12180 29374
rect 12684 29314 12740 29326
rect 12684 29262 12686 29314
rect 12738 29262 12740 29314
rect 12012 28438 12068 28476
rect 12572 28644 12628 28654
rect 10892 27990 10948 28028
rect 10780 26674 10836 26684
rect 12124 27860 12180 27870
rect 10332 26460 10836 26516
rect 10108 26404 10164 26414
rect 10164 26348 10276 26404
rect 10108 26338 10164 26348
rect 9772 26226 9828 26236
rect 8540 25676 8820 25732
rect 8316 25554 8372 25564
rect 8652 25508 8708 25518
rect 8428 25506 8708 25508
rect 8428 25454 8654 25506
rect 8706 25454 8708 25506
rect 8428 25452 8708 25454
rect 6412 23998 6414 24050
rect 6466 23998 6468 24050
rect 6412 23986 6468 23998
rect 6748 25284 6804 25294
rect 5852 23846 5908 23884
rect 5404 22306 5460 22316
rect 5852 23044 5908 23054
rect 3612 21858 3668 21868
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4956 19908 5012 19918
rect 5068 19908 5124 19918
rect 4956 19906 5068 19908
rect 4956 19854 4958 19906
rect 5010 19854 5068 19906
rect 4956 19852 5068 19854
rect 4956 19842 5012 19852
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4732 19348 4788 19358
rect 4732 19254 4788 19292
rect 4060 18564 4116 18574
rect 3500 18562 4116 18564
rect 3500 18510 4062 18562
rect 4114 18510 4116 18562
rect 3500 18508 4116 18510
rect 2604 18386 2660 18396
rect 3948 18340 4004 18350
rect 3948 18246 4004 18284
rect 4060 17892 4116 18508
rect 5068 18564 5124 19852
rect 5852 19908 5908 22988
rect 5852 19842 5908 19852
rect 6412 22932 6468 22942
rect 6412 21924 6468 22876
rect 5740 19346 5796 19358
rect 5740 19294 5742 19346
rect 5794 19294 5796 19346
rect 5292 18564 5348 18574
rect 4844 18340 4900 18350
rect 4844 18246 4900 18284
rect 4284 18228 4340 18238
rect 4284 18134 4340 18172
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4508 17892 4564 17902
rect 4060 17836 4508 17892
rect 4508 17778 4564 17836
rect 4508 17726 4510 17778
rect 4562 17726 4564 17778
rect 4508 17714 4564 17726
rect 5068 16996 5124 18508
rect 5180 18508 5292 18564
rect 5180 18450 5236 18508
rect 5292 18498 5348 18508
rect 5740 18564 5796 19294
rect 6076 19348 6132 19358
rect 6076 19234 6132 19292
rect 6076 19182 6078 19234
rect 6130 19182 6132 19234
rect 6076 19170 6132 19182
rect 5740 18498 5796 18508
rect 6076 18564 6132 18574
rect 5180 18398 5182 18450
rect 5234 18398 5236 18450
rect 5180 18386 5236 18398
rect 5628 18338 5684 18350
rect 5628 18286 5630 18338
rect 5682 18286 5684 18338
rect 5628 17666 5684 18286
rect 5964 18228 6020 18238
rect 5964 17778 6020 18172
rect 5964 17726 5966 17778
rect 6018 17726 6020 17778
rect 5964 17714 6020 17726
rect 5628 17614 5630 17666
rect 5682 17614 5684 17666
rect 5628 17602 5684 17614
rect 6076 17666 6132 18508
rect 6076 17614 6078 17666
rect 6130 17614 6132 17666
rect 6076 17602 6132 17614
rect 5068 16930 5124 16940
rect 5852 17442 5908 17454
rect 5852 17390 5854 17442
rect 5906 17390 5908 17442
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 5852 15988 5908 17390
rect 6188 17442 6244 17454
rect 6188 17390 6190 17442
rect 6242 17390 6244 17442
rect 5852 15922 5908 15932
rect 6076 16996 6132 17006
rect 6076 16882 6132 16940
rect 6076 16830 6078 16882
rect 6130 16830 6132 16882
rect 6076 15148 6132 16830
rect 6188 16884 6244 17390
rect 6188 16818 6244 16828
rect 5964 15092 6132 15148
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 5740 14642 5796 14654
rect 5740 14590 5742 14642
rect 5794 14590 5796 14642
rect 1932 14530 1988 14542
rect 1932 14478 1934 14530
rect 1986 14478 1988 14530
rect 1932 13524 1988 14478
rect 1932 10610 1988 13468
rect 2604 14418 2660 14430
rect 2604 14366 2606 14418
rect 2658 14366 2660 14418
rect 2604 13076 2660 14366
rect 4844 14308 4900 14318
rect 4844 14214 4900 14252
rect 5180 13634 5236 13646
rect 5180 13582 5182 13634
rect 5234 13582 5236 13634
rect 5180 13524 5236 13582
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 2604 13010 2660 13020
rect 4956 12850 5012 12862
rect 4956 12798 4958 12850
rect 5010 12798 5012 12850
rect 4956 12740 5012 12798
rect 5068 12852 5124 12862
rect 5068 12758 5124 12796
rect 4956 12674 5012 12684
rect 5068 11844 5124 11854
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4844 11732 4900 11742
rect 4396 11396 4452 11406
rect 4396 11302 4452 11340
rect 4844 11394 4900 11676
rect 4844 11342 4846 11394
rect 4898 11342 4900 11394
rect 4172 11284 4228 11294
rect 4172 11190 4228 11228
rect 2604 11172 2660 11182
rect 2604 10722 2660 11116
rect 4284 11172 4340 11182
rect 4284 11078 4340 11116
rect 2604 10670 2606 10722
rect 2658 10670 2660 10722
rect 2604 10658 2660 10670
rect 1932 10558 1934 10610
rect 1986 10558 1988 10610
rect 1932 10546 1988 10558
rect 4732 10500 4788 10510
rect 4844 10500 4900 11342
rect 5068 11282 5124 11788
rect 5068 11230 5070 11282
rect 5122 11230 5124 11282
rect 5068 11218 5124 11230
rect 4732 10498 4900 10500
rect 4732 10446 4734 10498
rect 4786 10446 4900 10498
rect 4732 10444 4900 10446
rect 5180 10498 5236 13468
rect 5740 13300 5796 14590
rect 5964 13524 6020 15092
rect 6188 14308 6244 14318
rect 6188 14214 6244 14252
rect 5964 13458 6020 13468
rect 5740 13244 6020 13300
rect 5740 13076 5796 13086
rect 5740 12982 5796 13020
rect 5628 12852 5684 12862
rect 5292 12850 5684 12852
rect 5292 12798 5630 12850
rect 5682 12798 5684 12850
rect 5292 12796 5684 12798
rect 5292 12402 5348 12796
rect 5292 12350 5294 12402
rect 5346 12350 5348 12402
rect 5292 12338 5348 12350
rect 5628 12404 5684 12796
rect 5852 12852 5908 12862
rect 5852 12758 5908 12796
rect 5964 12740 6020 13244
rect 6076 12964 6132 12974
rect 6076 12870 6132 12908
rect 6412 12964 6468 21868
rect 6748 21364 6804 25228
rect 8204 24836 8260 24846
rect 7644 24722 7700 24734
rect 7644 24670 7646 24722
rect 7698 24670 7700 24722
rect 6860 24052 6916 24062
rect 6860 23938 6916 23996
rect 7308 24052 7364 24062
rect 7308 23958 7364 23996
rect 6860 23886 6862 23938
rect 6914 23886 6916 23938
rect 6860 23874 6916 23886
rect 7420 23716 7476 23726
rect 7420 23622 7476 23660
rect 6860 23156 6916 23166
rect 6860 21586 6916 23100
rect 7644 23156 7700 24670
rect 8204 24722 8260 24780
rect 8204 24670 8206 24722
rect 8258 24670 8260 24722
rect 8204 24658 8260 24670
rect 7644 23090 7700 23100
rect 8428 23716 8484 25452
rect 8652 25442 8708 25452
rect 8764 25396 8820 25676
rect 8876 25620 8932 25630
rect 8876 25526 8932 25564
rect 8988 25396 9044 25406
rect 8764 25394 9044 25396
rect 8764 25342 8990 25394
rect 9042 25342 9044 25394
rect 8764 25340 9044 25342
rect 8988 24388 9044 25340
rect 8988 24322 9044 24332
rect 6860 21534 6862 21586
rect 6914 21534 6916 21586
rect 6860 21522 6916 21534
rect 7308 21586 7364 21598
rect 7308 21534 7310 21586
rect 7362 21534 7364 21586
rect 6748 21298 6804 21308
rect 6748 17444 6804 17454
rect 6748 16994 6804 17388
rect 6748 16942 6750 16994
rect 6802 16942 6804 16994
rect 6748 16930 6804 16942
rect 7308 13412 7364 21534
rect 7420 21588 7476 21598
rect 7420 21494 7476 21532
rect 8428 20802 8484 23660
rect 9996 21588 10052 21598
rect 10220 21588 10276 26348
rect 10780 26402 10836 26460
rect 10780 26350 10782 26402
rect 10834 26350 10836 26402
rect 10780 25732 10836 26350
rect 11116 26292 11172 26302
rect 11172 26236 11284 26292
rect 11116 26226 11172 26236
rect 10556 24388 10612 24398
rect 10444 23714 10500 23726
rect 10444 23662 10446 23714
rect 10498 23662 10500 23714
rect 9996 21586 10276 21588
rect 9996 21534 9998 21586
rect 10050 21534 10276 21586
rect 9996 21532 10276 21534
rect 10332 21698 10388 21710
rect 10332 21646 10334 21698
rect 10386 21646 10388 21698
rect 9996 21522 10052 21532
rect 8428 20750 8430 20802
rect 8482 20750 8484 20802
rect 8428 20738 8484 20750
rect 9436 20802 9492 20814
rect 9436 20750 9438 20802
rect 9490 20750 9492 20802
rect 9212 20690 9268 20702
rect 9212 20638 9214 20690
rect 9266 20638 9268 20690
rect 8428 20578 8484 20590
rect 8428 20526 8430 20578
rect 8482 20526 8484 20578
rect 8428 20018 8484 20526
rect 9212 20356 9268 20638
rect 9324 20580 9380 20590
rect 9324 20486 9380 20524
rect 8988 20300 9268 20356
rect 8988 20242 9044 20300
rect 8988 20190 8990 20242
rect 9042 20190 9044 20242
rect 8988 20178 9044 20190
rect 8540 20132 8596 20142
rect 8540 20038 8596 20076
rect 8428 19966 8430 20018
rect 8482 19966 8484 20018
rect 8428 19348 8484 19966
rect 8876 20020 8932 20030
rect 8876 19926 8932 19964
rect 8428 19282 8484 19292
rect 9436 18452 9492 20750
rect 9996 20804 10052 20814
rect 9996 20132 10052 20748
rect 9884 20130 10052 20132
rect 9884 20078 9998 20130
rect 10050 20078 10052 20130
rect 9884 20076 10052 20078
rect 9884 19458 9940 20076
rect 9996 20066 10052 20076
rect 10108 20578 10164 20590
rect 10108 20526 10110 20578
rect 10162 20526 10164 20578
rect 10108 19908 10164 20526
rect 10220 20244 10276 20254
rect 10332 20244 10388 21646
rect 10220 20242 10388 20244
rect 10220 20190 10222 20242
rect 10274 20190 10388 20242
rect 10220 20188 10388 20190
rect 10220 20132 10276 20188
rect 10220 20066 10276 20076
rect 10444 20130 10500 23662
rect 10556 20802 10612 24332
rect 10780 23938 10836 25676
rect 10780 23886 10782 23938
rect 10834 23886 10836 23938
rect 10780 23874 10836 23886
rect 11116 23938 11172 23950
rect 11116 23886 11118 23938
rect 11170 23886 11172 23938
rect 10556 20750 10558 20802
rect 10610 20750 10612 20802
rect 10556 20738 10612 20750
rect 10780 23156 10836 23166
rect 11116 23156 11172 23886
rect 10780 23154 11172 23156
rect 10780 23102 10782 23154
rect 10834 23102 11172 23154
rect 10780 23100 11172 23102
rect 10780 20468 10836 23100
rect 10892 20804 10948 20814
rect 10892 20710 10948 20748
rect 11228 20690 11284 26236
rect 11788 25508 11844 25518
rect 11788 25414 11844 25452
rect 12124 24724 12180 27804
rect 12572 27412 12628 28588
rect 12572 27346 12628 27356
rect 12684 26852 12740 29262
rect 13468 28642 13524 28654
rect 13468 28590 13470 28642
rect 13522 28590 13524 28642
rect 12684 26786 12740 26796
rect 12796 28532 12852 28542
rect 12236 26404 12292 26414
rect 12236 26292 12292 26348
rect 12684 26292 12740 26302
rect 12236 26290 12516 26292
rect 12236 26238 12238 26290
rect 12290 26238 12516 26290
rect 12236 26236 12516 26238
rect 12236 26226 12292 26236
rect 12236 25732 12292 25742
rect 12236 25638 12292 25676
rect 12460 25730 12516 26236
rect 12684 26198 12740 26236
rect 12460 25678 12462 25730
rect 12514 25678 12516 25730
rect 12460 25666 12516 25678
rect 12684 25508 12740 25518
rect 12796 25508 12852 28476
rect 13468 27860 13524 28590
rect 13580 28532 13636 30156
rect 14028 30098 14084 30110
rect 14028 30046 14030 30098
rect 14082 30046 14084 30098
rect 13916 29428 13972 29438
rect 13916 28642 13972 29372
rect 13916 28590 13918 28642
rect 13970 28590 13972 28642
rect 13916 28578 13972 28590
rect 14028 28644 14084 30046
rect 15932 30100 15988 30830
rect 16492 30882 16548 30940
rect 16492 30830 16494 30882
rect 16546 30830 16548 30882
rect 15932 30034 15988 30044
rect 16044 30210 16100 30222
rect 16044 30158 16046 30210
rect 16098 30158 16100 30210
rect 16044 29988 16100 30158
rect 16044 29922 16100 29932
rect 16492 29988 16548 30830
rect 16828 30884 16884 31836
rect 16828 30322 16884 30828
rect 16828 30270 16830 30322
rect 16882 30270 16884 30322
rect 16828 30258 16884 30270
rect 16940 31892 17332 31948
rect 20412 31948 20468 36316
rect 20748 35028 20804 36316
rect 20972 35810 21028 36428
rect 20972 35758 20974 35810
rect 21026 35758 21028 35810
rect 20972 35746 21028 35758
rect 21756 36372 21812 36382
rect 21756 35812 21812 36316
rect 21644 35698 21700 35710
rect 21644 35646 21646 35698
rect 21698 35646 21700 35698
rect 20748 35026 21364 35028
rect 20748 34974 20750 35026
rect 20802 34974 21364 35026
rect 20748 34972 21364 34974
rect 20748 34962 20804 34972
rect 21308 34914 21364 34972
rect 21308 34862 21310 34914
rect 21362 34862 21364 34914
rect 21308 34850 21364 34862
rect 21644 34916 21700 35646
rect 21756 35586 21812 35756
rect 21756 35534 21758 35586
rect 21810 35534 21812 35586
rect 21756 35522 21812 35534
rect 23436 35476 23492 37886
rect 25228 37268 25284 37278
rect 25452 37268 25508 38108
rect 25564 38098 25620 38108
rect 26012 38164 26068 38174
rect 26012 38070 26068 38108
rect 28364 38164 28420 39564
rect 28364 38098 28420 38108
rect 25564 37380 25620 37390
rect 25564 37378 25732 37380
rect 25564 37326 25566 37378
rect 25618 37326 25732 37378
rect 25564 37324 25732 37326
rect 25564 37314 25620 37324
rect 25116 37266 25508 37268
rect 25116 37214 25230 37266
rect 25282 37214 25508 37266
rect 25116 37212 25508 37214
rect 24556 36708 24612 36718
rect 24556 36594 24612 36652
rect 24556 36542 24558 36594
rect 24610 36542 24612 36594
rect 24556 36530 24612 36542
rect 24780 36484 24836 36494
rect 25116 36484 25172 37212
rect 25228 37202 25284 37212
rect 25564 36708 25620 36718
rect 25564 36614 25620 36652
rect 25676 36484 25732 37324
rect 28700 37154 28756 37166
rect 28700 37102 28702 37154
rect 28754 37102 28756 37154
rect 26460 36708 26516 36718
rect 24780 36482 25172 36484
rect 24780 36430 24782 36482
rect 24834 36430 25172 36482
rect 24780 36428 25172 36430
rect 25564 36428 26404 36484
rect 24780 36418 24836 36428
rect 24108 36372 24164 36382
rect 24108 36278 24164 36316
rect 25228 35700 25284 35710
rect 25228 35606 25284 35644
rect 23436 35410 23492 35420
rect 24220 35476 24276 35486
rect 24276 35420 24388 35476
rect 24220 35410 24276 35420
rect 21644 34850 21700 34860
rect 21644 34692 21700 34702
rect 21644 34690 21924 34692
rect 21644 34638 21646 34690
rect 21698 34638 21924 34690
rect 21644 34636 21924 34638
rect 21644 34626 21700 34636
rect 20412 31892 21140 31948
rect 16492 29922 16548 29932
rect 16940 29652 16996 31892
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 18284 30884 18340 30894
rect 16716 29596 16996 29652
rect 17500 30100 17556 30110
rect 17500 29650 17556 30044
rect 17500 29598 17502 29650
rect 17554 29598 17556 29650
rect 14476 29540 14532 29550
rect 14476 29446 14532 29484
rect 15484 29538 15540 29550
rect 15484 29486 15486 29538
rect 15538 29486 15540 29538
rect 14364 29428 14420 29438
rect 14364 29334 14420 29372
rect 15484 29428 15540 29486
rect 15484 29204 15540 29372
rect 16156 29540 16212 29550
rect 15596 29316 15652 29326
rect 15596 29222 15652 29260
rect 15484 29138 15540 29148
rect 15708 29202 15764 29214
rect 15708 29150 15710 29202
rect 15762 29150 15764 29202
rect 15708 28980 15764 29150
rect 15708 28914 15764 28924
rect 15932 29092 15988 29102
rect 15932 28756 15988 29036
rect 16156 28868 16212 29484
rect 16268 29426 16324 29438
rect 16268 29374 16270 29426
rect 16322 29374 16324 29426
rect 16268 29092 16324 29374
rect 16268 29026 16324 29036
rect 16380 29426 16436 29438
rect 16380 29374 16382 29426
rect 16434 29374 16436 29426
rect 16380 28980 16436 29374
rect 16156 28812 16324 28868
rect 15932 28690 15988 28700
rect 14028 28578 14084 28588
rect 15148 28644 15204 28654
rect 13580 28466 13636 28476
rect 13468 27794 13524 27804
rect 14140 27188 14196 27198
rect 14140 27094 14196 27132
rect 15036 27186 15092 27198
rect 15036 27134 15038 27186
rect 15090 27134 15092 27186
rect 14924 27074 14980 27086
rect 14924 27022 14926 27074
rect 14978 27022 14980 27074
rect 14476 26962 14532 26974
rect 14476 26910 14478 26962
rect 14530 26910 14532 26962
rect 14476 26908 14532 26910
rect 14364 26852 14532 26908
rect 14364 26516 14420 26852
rect 14364 26422 14420 26460
rect 14476 26628 14532 26638
rect 14476 26404 14532 26572
rect 14476 26402 14644 26404
rect 14476 26350 14478 26402
rect 14530 26350 14644 26402
rect 14476 26348 14644 26350
rect 14476 26338 14532 26348
rect 12684 25506 12852 25508
rect 12684 25454 12686 25506
rect 12738 25454 12852 25506
rect 12684 25452 12852 25454
rect 12684 25442 12740 25452
rect 12460 24836 12516 24846
rect 12460 24742 12516 24780
rect 12348 24724 12404 24734
rect 11676 24722 12404 24724
rect 11676 24670 12350 24722
rect 12402 24670 12404 24722
rect 11676 24668 12404 24670
rect 11676 23826 11732 24668
rect 12348 24658 12404 24668
rect 11676 23774 11678 23826
rect 11730 23774 11732 23826
rect 11340 23714 11396 23726
rect 11340 23662 11342 23714
rect 11394 23662 11396 23714
rect 11340 23156 11396 23662
rect 11340 23090 11396 23100
rect 11676 23154 11732 23774
rect 11676 23102 11678 23154
rect 11730 23102 11732 23154
rect 11676 23090 11732 23102
rect 12684 23156 12740 23166
rect 12684 23062 12740 23100
rect 12796 21700 12852 25452
rect 14364 25508 14420 25518
rect 14364 25414 14420 25452
rect 12908 25396 12964 25406
rect 12908 25394 13076 25396
rect 12908 25342 12910 25394
rect 12962 25342 13076 25394
rect 12908 25340 13076 25342
rect 12908 25330 12964 25340
rect 13020 22260 13076 25340
rect 14476 24724 14532 24734
rect 13804 23154 13860 23166
rect 13804 23102 13806 23154
rect 13858 23102 13860 23154
rect 13804 22596 13860 23102
rect 14476 23042 14532 24668
rect 14476 22990 14478 23042
rect 14530 22990 14532 23042
rect 14476 22978 14532 22990
rect 13020 22194 13076 22204
rect 13356 22540 13860 22596
rect 12908 21700 12964 21710
rect 12796 21698 12964 21700
rect 12796 21646 12910 21698
rect 12962 21646 12964 21698
rect 12796 21644 12964 21646
rect 12908 21634 12964 21644
rect 11340 21588 11396 21598
rect 11340 21494 11396 21532
rect 13356 21586 13412 22540
rect 13468 22372 13524 22382
rect 14364 22372 14420 22382
rect 13468 22278 13524 22316
rect 14140 22370 14420 22372
rect 14140 22318 14366 22370
rect 14418 22318 14420 22370
rect 14140 22316 14420 22318
rect 13692 22146 13748 22158
rect 13692 22094 13694 22146
rect 13746 22094 13748 22146
rect 13580 21812 13636 21822
rect 13580 21718 13636 21756
rect 13356 21534 13358 21586
rect 13410 21534 13412 21586
rect 11228 20638 11230 20690
rect 11282 20638 11284 20690
rect 11228 20626 11284 20638
rect 11340 20914 11396 20926
rect 11340 20862 11342 20914
rect 11394 20862 11396 20914
rect 11340 20692 11396 20862
rect 11340 20626 11396 20636
rect 10780 20412 11060 20468
rect 10444 20078 10446 20130
rect 10498 20078 10500 20130
rect 10444 20020 10500 20078
rect 10780 20020 10836 20030
rect 10444 20018 10836 20020
rect 10444 19966 10782 20018
rect 10834 19966 10836 20018
rect 10444 19964 10836 19966
rect 10780 19954 10836 19964
rect 10220 19908 10276 19918
rect 9884 19406 9886 19458
rect 9938 19406 9940 19458
rect 9884 19394 9940 19406
rect 9996 19852 10220 19908
rect 9772 19124 9828 19134
rect 9436 18386 9492 18396
rect 9548 19122 9828 19124
rect 9548 19070 9774 19122
rect 9826 19070 9828 19122
rect 9548 19068 9828 19070
rect 9548 17668 9604 19068
rect 9772 19058 9828 19068
rect 8876 17612 9604 17668
rect 8876 16770 8932 17612
rect 8876 16718 8878 16770
rect 8930 16718 8932 16770
rect 8876 16706 8932 16718
rect 9436 17442 9492 17454
rect 9436 17390 9438 17442
rect 9490 17390 9492 17442
rect 9436 15148 9492 17390
rect 9548 16100 9604 17612
rect 9884 17668 9940 17678
rect 9996 17668 10052 19852
rect 10220 19842 10276 19852
rect 10332 19908 10388 19918
rect 10892 19908 10948 19918
rect 10332 19906 10500 19908
rect 10332 19854 10334 19906
rect 10386 19854 10500 19906
rect 10332 19852 10500 19854
rect 10332 19842 10388 19852
rect 10444 18900 10500 19852
rect 10892 19814 10948 19852
rect 11004 19684 11060 20412
rect 10892 19628 11060 19684
rect 11228 20244 11284 20254
rect 10444 18844 10836 18900
rect 10220 18676 10276 18686
rect 9884 17666 10052 17668
rect 9884 17614 9886 17666
rect 9938 17614 10052 17666
rect 9884 17612 10052 17614
rect 10108 18564 10164 18574
rect 10108 17666 10164 18508
rect 10108 17614 10110 17666
rect 10162 17614 10164 17666
rect 9884 17602 9940 17612
rect 10108 17602 10164 17614
rect 10220 17668 10276 18620
rect 10556 18674 10612 18686
rect 10556 18622 10558 18674
rect 10610 18622 10612 18674
rect 10556 18564 10612 18622
rect 10444 18452 10500 18462
rect 10444 17892 10500 18396
rect 10220 17666 10388 17668
rect 10220 17614 10222 17666
rect 10274 17614 10388 17666
rect 10220 17612 10388 17614
rect 10220 17602 10276 17612
rect 9660 16996 9716 17006
rect 10220 16996 10276 17006
rect 9716 16994 10276 16996
rect 9716 16942 10222 16994
rect 10274 16942 10276 16994
rect 9716 16940 10276 16942
rect 9660 16902 9716 16940
rect 10220 16930 10276 16940
rect 10220 16212 10276 16222
rect 10332 16212 10388 17612
rect 10444 17666 10500 17836
rect 10444 17614 10446 17666
rect 10498 17614 10500 17666
rect 10444 17602 10500 17614
rect 10220 16210 10388 16212
rect 10220 16158 10222 16210
rect 10274 16158 10388 16210
rect 10220 16156 10388 16158
rect 10220 16146 10276 16156
rect 9660 16100 9716 16110
rect 9548 16098 9716 16100
rect 9548 16046 9662 16098
rect 9714 16046 9716 16098
rect 9548 16044 9716 16046
rect 9660 16034 9716 16044
rect 10556 16098 10612 18508
rect 10668 18676 10724 18686
rect 10668 18562 10724 18620
rect 10668 18510 10670 18562
rect 10722 18510 10724 18562
rect 10668 18498 10724 18510
rect 10556 16046 10558 16098
rect 10610 16046 10612 16098
rect 10556 16034 10612 16046
rect 10780 16098 10836 18844
rect 10780 16046 10782 16098
rect 10834 16046 10836 16098
rect 10780 16034 10836 16046
rect 10892 15148 10948 19628
rect 11228 18676 11284 20188
rect 11452 19908 11508 19918
rect 11452 19348 11508 19852
rect 11452 19282 11508 19292
rect 11284 18620 11396 18676
rect 11228 18610 11284 18620
rect 11004 18450 11060 18462
rect 11004 18398 11006 18450
rect 11058 18398 11060 18450
rect 11004 18340 11060 18398
rect 11004 18274 11060 18284
rect 11228 17666 11284 17678
rect 11228 17614 11230 17666
rect 11282 17614 11284 17666
rect 11004 17554 11060 17566
rect 11004 17502 11006 17554
rect 11058 17502 11060 17554
rect 11004 16210 11060 17502
rect 11116 17444 11172 17454
rect 11116 17350 11172 17388
rect 11004 16158 11006 16210
rect 11058 16158 11060 16210
rect 11004 16146 11060 16158
rect 11228 16098 11284 17614
rect 11228 16046 11230 16098
rect 11282 16046 11284 16098
rect 11228 16034 11284 16046
rect 11004 15988 11060 15998
rect 11340 15988 11396 18620
rect 11452 17780 11508 17790
rect 11452 17666 11508 17724
rect 12012 17780 12068 17790
rect 12012 17686 12068 17724
rect 11452 17614 11454 17666
rect 11506 17614 11508 17666
rect 11452 17602 11508 17614
rect 11564 16884 11620 16894
rect 11564 16098 11620 16828
rect 11564 16046 11566 16098
rect 11618 16046 11620 16098
rect 11452 15988 11508 15998
rect 11340 15986 11508 15988
rect 11340 15934 11454 15986
rect 11506 15934 11508 15986
rect 11340 15932 11508 15934
rect 11004 15894 11060 15932
rect 11452 15922 11508 15932
rect 8764 15092 9492 15148
rect 10668 15092 10948 15148
rect 11564 15148 11620 16046
rect 12908 16100 12964 16110
rect 12908 16006 12964 16044
rect 11900 15988 11956 15998
rect 11564 15092 11732 15148
rect 8540 13972 8596 13982
rect 6972 13076 7028 13086
rect 6972 12964 7028 13020
rect 6412 12962 6692 12964
rect 6412 12910 6414 12962
rect 6466 12910 6692 12962
rect 6412 12908 6692 12910
rect 6412 12898 6468 12908
rect 5964 12674 6020 12684
rect 6636 12516 6692 12908
rect 5628 12348 5796 12404
rect 5516 12290 5572 12302
rect 5516 12238 5518 12290
rect 5570 12238 5572 12290
rect 5516 11844 5572 12238
rect 5628 12180 5684 12190
rect 5628 12086 5684 12124
rect 5516 11778 5572 11788
rect 5740 11394 5796 12348
rect 6636 12402 6692 12460
rect 6636 12350 6638 12402
rect 6690 12350 6692 12402
rect 6636 12338 6692 12350
rect 6748 12962 7028 12964
rect 6748 12910 6974 12962
rect 7026 12910 7028 12962
rect 6748 12908 7028 12910
rect 6748 12180 6804 12908
rect 6972 12898 7028 12908
rect 7196 12740 7252 12750
rect 5740 11342 5742 11394
rect 5794 11342 5796 11394
rect 5740 11330 5796 11342
rect 6076 11844 6132 11854
rect 6748 11844 6804 12124
rect 6076 11394 6132 11788
rect 6076 11342 6078 11394
rect 6130 11342 6132 11394
rect 6076 11330 6132 11342
rect 6636 11788 6804 11844
rect 6860 12738 7252 12740
rect 6860 12686 7198 12738
rect 7250 12686 7252 12738
rect 6860 12684 7252 12686
rect 6860 11844 6916 12684
rect 7196 12674 7252 12684
rect 6636 11394 6692 11788
rect 6636 11342 6638 11394
rect 6690 11342 6692 11394
rect 6636 11330 6692 11342
rect 6748 11396 6804 11406
rect 6748 11302 6804 11340
rect 6860 11394 6916 11788
rect 7308 11732 7364 13356
rect 8428 13412 8484 13422
rect 8428 12962 8484 13356
rect 8428 12910 8430 12962
rect 8482 12910 8484 12962
rect 8428 12898 8484 12910
rect 7420 12852 7476 12862
rect 7420 12758 7476 12796
rect 7532 12738 7588 12750
rect 7532 12686 7534 12738
rect 7586 12686 7588 12738
rect 7532 12292 7588 12686
rect 8540 12402 8596 13916
rect 8764 13076 8820 15092
rect 10668 14308 10724 15092
rect 10668 14242 10724 14252
rect 9996 13972 10052 13982
rect 9996 13878 10052 13916
rect 11676 13970 11732 15092
rect 11676 13918 11678 13970
rect 11730 13918 11732 13970
rect 8540 12350 8542 12402
rect 8594 12350 8596 12402
rect 8540 12338 8596 12350
rect 8652 12964 8708 12974
rect 8652 12402 8708 12908
rect 8764 12850 8820 13020
rect 9548 13746 9604 13758
rect 9548 13694 9550 13746
rect 9602 13694 9604 13746
rect 8988 12964 9044 12974
rect 8764 12798 8766 12850
rect 8818 12798 8820 12850
rect 8764 12786 8820 12798
rect 8876 12852 8932 12862
rect 8652 12350 8654 12402
rect 8706 12350 8708 12402
rect 8652 12338 8708 12350
rect 8764 12404 8820 12414
rect 8876 12404 8932 12796
rect 8764 12402 8932 12404
rect 8764 12350 8766 12402
rect 8818 12350 8932 12402
rect 8764 12348 8932 12350
rect 8764 12338 8820 12348
rect 7532 12226 7588 12236
rect 8316 12292 8372 12302
rect 8316 12198 8372 12236
rect 8988 12178 9044 12908
rect 9548 12964 9604 13694
rect 9548 12898 9604 12908
rect 9772 13746 9828 13758
rect 9772 13694 9774 13746
rect 9826 13694 9828 13746
rect 9772 12852 9828 13694
rect 10220 13748 10276 13758
rect 9884 13634 9940 13646
rect 9884 13582 9886 13634
rect 9938 13582 9940 13634
rect 9884 13188 9940 13582
rect 9884 13132 10052 13188
rect 9660 12850 9828 12852
rect 9660 12798 9774 12850
rect 9826 12798 9828 12850
rect 9660 12796 9828 12798
rect 8988 12126 8990 12178
rect 9042 12126 9044 12178
rect 8988 12114 9044 12126
rect 9436 12404 9492 12414
rect 7308 11666 7364 11676
rect 6860 11342 6862 11394
rect 6914 11342 6916 11394
rect 6860 11330 6916 11342
rect 5964 11284 6020 11294
rect 5964 11190 6020 11228
rect 5852 11172 5908 11182
rect 5852 11078 5908 11116
rect 6188 11170 6244 11182
rect 6188 11118 6190 11170
rect 6242 11118 6244 11170
rect 6188 10836 6244 11118
rect 7084 11170 7140 11182
rect 7084 11118 7086 11170
rect 7138 11118 7140 11170
rect 7084 11060 7140 11118
rect 7084 10994 7140 11004
rect 7644 11170 7700 11182
rect 7644 11118 7646 11170
rect 7698 11118 7700 11170
rect 7644 11060 7700 11118
rect 7644 10994 7700 11004
rect 6188 10770 6244 10780
rect 5180 10446 5182 10498
rect 5234 10446 5236 10498
rect 4732 10434 4788 10444
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 5180 8036 5236 10446
rect 7756 9940 7812 9950
rect 7756 8370 7812 9884
rect 9436 9940 9492 12348
rect 9548 12292 9604 12302
rect 9548 12198 9604 12236
rect 9436 9874 9492 9884
rect 9660 12180 9716 12796
rect 9772 12786 9828 12796
rect 9884 12962 9940 12974
rect 9884 12910 9886 12962
rect 9938 12910 9940 12962
rect 9884 12852 9940 12910
rect 9884 12786 9940 12796
rect 9996 12628 10052 13132
rect 10220 13074 10276 13692
rect 10220 13022 10222 13074
rect 10274 13022 10276 13074
rect 10220 13010 10276 13022
rect 9884 12572 10052 12628
rect 9772 12404 9828 12442
rect 9772 12338 9828 12348
rect 9660 8428 9716 12124
rect 9772 12178 9828 12190
rect 9772 12126 9774 12178
rect 9826 12126 9828 12178
rect 9772 12068 9828 12126
rect 9884 12180 9940 12572
rect 10108 12516 10164 12526
rect 9996 12180 10052 12190
rect 9884 12178 10052 12180
rect 9884 12126 9998 12178
rect 10050 12126 10052 12178
rect 9884 12124 10052 12126
rect 9996 12114 10052 12124
rect 10108 12178 10164 12460
rect 11452 12516 11508 12526
rect 11004 12404 11060 12414
rect 11004 12290 11060 12348
rect 11452 12402 11508 12460
rect 11452 12350 11454 12402
rect 11506 12350 11508 12402
rect 11452 12338 11508 12350
rect 11004 12238 11006 12290
rect 11058 12238 11060 12290
rect 10108 12126 10110 12178
rect 10162 12126 10164 12178
rect 10108 12114 10164 12126
rect 10668 12180 10724 12190
rect 10668 12086 10724 12124
rect 9772 12002 9828 12012
rect 11004 12068 11060 12238
rect 11004 12002 11060 12012
rect 11676 10836 11732 13918
rect 11900 11172 11956 15932
rect 12572 15988 12628 15998
rect 12572 15894 12628 15932
rect 12460 15092 12516 15102
rect 12012 13972 12068 13982
rect 12460 13972 12516 15036
rect 12012 13970 12516 13972
rect 12012 13918 12014 13970
rect 12066 13918 12462 13970
rect 12514 13918 12516 13970
rect 12012 13916 12516 13918
rect 12012 13906 12068 13916
rect 12236 13076 12292 13916
rect 12460 13906 12516 13916
rect 12908 13076 12964 13086
rect 12236 13074 12964 13076
rect 12236 13022 12910 13074
rect 12962 13022 12964 13074
rect 12236 13020 12964 13022
rect 12236 12962 12292 13020
rect 12908 13010 12964 13020
rect 12236 12910 12238 12962
rect 12290 12910 12292 12962
rect 12236 12898 12292 12910
rect 12460 12852 12516 12862
rect 12460 12758 12516 12796
rect 13244 12516 13300 12526
rect 12012 11172 12068 11182
rect 11900 11116 12012 11172
rect 11676 10742 11732 10780
rect 12012 10834 12068 11116
rect 12012 10782 12014 10834
rect 12066 10782 12068 10834
rect 12012 10770 12068 10782
rect 12908 11172 12964 11182
rect 11788 10612 11844 10622
rect 11788 10518 11844 10556
rect 12124 10610 12180 10622
rect 12124 10558 12126 10610
rect 12178 10558 12180 10610
rect 11900 10498 11956 10510
rect 11900 10446 11902 10498
rect 11954 10446 11956 10498
rect 11900 10276 11956 10446
rect 11340 10220 11956 10276
rect 11228 9940 11284 9950
rect 10892 9938 11284 9940
rect 10892 9886 11230 9938
rect 11282 9886 11284 9938
rect 10892 9884 11284 9886
rect 9660 8372 9940 8428
rect 7756 8318 7758 8370
rect 7810 8318 7812 8370
rect 7756 8306 7812 8318
rect 9884 8370 9940 8372
rect 9884 8318 9886 8370
rect 9938 8318 9940 8370
rect 9884 8306 9940 8318
rect 5180 7970 5236 7980
rect 7084 8258 7140 8270
rect 7084 8206 7086 8258
rect 7138 8206 7140 8258
rect 7084 8036 7140 8206
rect 7084 7970 7140 7980
rect 10556 8036 10612 8046
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 10220 5908 10276 5918
rect 10220 5814 10276 5852
rect 10556 5908 10612 7980
rect 10892 6018 10948 9884
rect 11228 9874 11284 9884
rect 11340 9714 11396 10220
rect 12012 10164 12068 10174
rect 11340 9662 11342 9714
rect 11394 9662 11396 9714
rect 11340 9650 11396 9662
rect 11564 9716 11620 9726
rect 11564 9622 11620 9660
rect 12012 9714 12068 10108
rect 12012 9662 12014 9714
rect 12066 9662 12068 9714
rect 12012 9650 12068 9662
rect 12124 9940 12180 10558
rect 12124 9380 12180 9884
rect 12236 10612 12292 10622
rect 12236 9940 12292 10556
rect 12908 10164 12964 11116
rect 13244 10836 13300 12460
rect 13356 12404 13412 21534
rect 13692 20244 13748 22094
rect 13804 22146 13860 22158
rect 13804 22094 13806 22146
rect 13858 22094 13860 22146
rect 13804 20802 13860 22094
rect 13804 20750 13806 20802
rect 13858 20750 13860 20802
rect 13804 20738 13860 20750
rect 14028 20690 14084 20702
rect 14028 20638 14030 20690
rect 14082 20638 14084 20690
rect 14028 20580 14084 20638
rect 14028 20514 14084 20524
rect 13692 20178 13748 20188
rect 13804 18452 13860 18462
rect 13468 18450 13860 18452
rect 13468 18398 13806 18450
rect 13858 18398 13860 18450
rect 13468 18396 13860 18398
rect 13468 15986 13524 18396
rect 13804 18386 13860 18396
rect 14028 17668 14084 17678
rect 14028 17574 14084 17612
rect 13804 16100 13860 16110
rect 13804 16006 13860 16044
rect 13468 15934 13470 15986
rect 13522 15934 13524 15986
rect 13468 15148 13524 15934
rect 14140 15148 14196 22316
rect 14364 22306 14420 22316
rect 14476 22260 14532 22270
rect 14476 22166 14532 22204
rect 14588 20020 14644 26348
rect 14924 26292 14980 27022
rect 14924 26226 14980 26236
rect 15036 23380 15092 27134
rect 15148 24724 15204 28588
rect 16044 28644 16100 28654
rect 16044 28550 16100 28588
rect 16268 28642 16324 28812
rect 16268 28590 16270 28642
rect 16322 28590 16324 28642
rect 16268 28578 16324 28590
rect 16380 28642 16436 28924
rect 16380 28590 16382 28642
rect 16434 28590 16436 28642
rect 16380 28578 16436 28590
rect 16716 28196 16772 29596
rect 17500 29586 17556 29598
rect 17612 29538 17668 29550
rect 17612 29486 17614 29538
rect 17666 29486 17668 29538
rect 17388 29428 17444 29438
rect 17164 29426 17444 29428
rect 17164 29374 17390 29426
rect 17442 29374 17444 29426
rect 17164 29372 17444 29374
rect 16828 29316 16884 29326
rect 17164 29316 17220 29372
rect 17388 29362 17444 29372
rect 17500 29428 17556 29438
rect 16828 29314 17220 29316
rect 16828 29262 16830 29314
rect 16882 29262 17220 29314
rect 16828 29260 17220 29262
rect 16828 29250 16884 29260
rect 17388 28980 17444 28990
rect 17276 28756 17332 28766
rect 17276 28662 17332 28700
rect 16828 28418 16884 28430
rect 16828 28366 16830 28418
rect 16882 28366 16884 28418
rect 16828 28308 16884 28366
rect 16828 28252 17220 28308
rect 16716 28140 16884 28196
rect 15484 27746 15540 27758
rect 15484 27694 15486 27746
rect 15538 27694 15540 27746
rect 15260 27188 15316 27198
rect 15484 27188 15540 27694
rect 15820 27188 15876 27198
rect 16156 27188 16212 27198
rect 15316 27186 15876 27188
rect 15316 27134 15822 27186
rect 15874 27134 15876 27186
rect 15316 27132 15876 27134
rect 15260 27074 15316 27132
rect 15820 27122 15876 27132
rect 15932 27132 16156 27188
rect 15260 27022 15262 27074
rect 15314 27022 15316 27074
rect 15260 27010 15316 27022
rect 15596 26852 15652 26862
rect 15260 26516 15316 26526
rect 15260 26402 15316 26460
rect 15260 26350 15262 26402
rect 15314 26350 15316 26402
rect 15260 26338 15316 26350
rect 15596 25506 15652 26796
rect 15820 26404 15876 26414
rect 15932 26404 15988 27132
rect 16156 27094 16212 27132
rect 15820 26402 15988 26404
rect 15820 26350 15822 26402
rect 15874 26350 15988 26402
rect 15820 26348 15988 26350
rect 15820 26338 15876 26348
rect 15596 25454 15598 25506
rect 15650 25454 15652 25506
rect 15596 25442 15652 25454
rect 16044 26292 16100 26302
rect 16044 24946 16100 26236
rect 16268 26292 16324 26302
rect 16156 26180 16212 26190
rect 16156 26086 16212 26124
rect 16044 24894 16046 24946
rect 16098 24894 16100 24946
rect 16044 24882 16100 24894
rect 15148 24658 15204 24668
rect 16156 24836 16212 24846
rect 16268 24836 16324 26236
rect 16156 24834 16324 24836
rect 16156 24782 16158 24834
rect 16210 24782 16324 24834
rect 16156 24780 16324 24782
rect 16380 25284 16436 25294
rect 16156 24388 16212 24780
rect 15932 24332 16212 24388
rect 15036 23314 15092 23324
rect 15148 23938 15204 23950
rect 15148 23886 15150 23938
rect 15202 23886 15204 23938
rect 14700 22932 14756 22942
rect 15148 22932 15204 23886
rect 14700 22930 15204 22932
rect 14700 22878 14702 22930
rect 14754 22878 15204 22930
rect 14700 22876 15204 22878
rect 14700 22866 14756 22876
rect 15148 22484 15204 22876
rect 15148 22418 15204 22428
rect 15372 23380 15428 23390
rect 15372 22372 15428 23324
rect 15932 23378 15988 24332
rect 16380 24276 16436 25228
rect 15932 23326 15934 23378
rect 15986 23326 15988 23378
rect 15932 22708 15988 23326
rect 15932 22642 15988 22652
rect 16044 24220 16436 24276
rect 16044 23042 16100 24220
rect 16828 24052 16884 28140
rect 17164 27074 17220 28252
rect 17388 27970 17444 28924
rect 17388 27918 17390 27970
rect 17442 27918 17444 27970
rect 17388 27906 17444 27918
rect 17500 27748 17556 29372
rect 17612 28644 17668 29486
rect 17836 29428 17892 29438
rect 17836 29426 18004 29428
rect 17836 29374 17838 29426
rect 17890 29374 18004 29426
rect 17836 29372 18004 29374
rect 17836 29362 17892 29372
rect 17612 28578 17668 28588
rect 17612 27860 17668 27870
rect 17612 27858 17780 27860
rect 17612 27806 17614 27858
rect 17666 27806 17780 27858
rect 17612 27804 17780 27806
rect 17612 27794 17668 27804
rect 17164 27022 17166 27074
rect 17218 27022 17220 27074
rect 17164 26516 17220 27022
rect 17388 27692 17556 27748
rect 17276 26852 17332 26862
rect 17276 26758 17332 26796
rect 17388 26850 17444 27692
rect 17724 27074 17780 27804
rect 17724 27022 17726 27074
rect 17778 27022 17780 27074
rect 17724 26964 17780 27022
rect 17724 26898 17780 26908
rect 17836 27858 17892 27870
rect 17836 27806 17838 27858
rect 17890 27806 17892 27858
rect 17836 27188 17892 27806
rect 17388 26798 17390 26850
rect 17442 26798 17444 26850
rect 17388 26786 17444 26798
rect 17164 26460 17780 26516
rect 17724 26402 17780 26460
rect 17724 26350 17726 26402
rect 17778 26350 17780 26402
rect 17724 26338 17780 26350
rect 17388 26292 17444 26302
rect 17388 26198 17444 26236
rect 17612 26290 17668 26302
rect 17612 26238 17614 26290
rect 17666 26238 17668 26290
rect 17612 26180 17668 26238
rect 17836 26180 17892 27132
rect 17948 26852 18004 29372
rect 18060 29426 18116 29438
rect 18060 29374 18062 29426
rect 18114 29374 18116 29426
rect 18060 28756 18116 29374
rect 18060 28690 18116 28700
rect 18172 29428 18228 29438
rect 18172 28082 18228 29372
rect 18172 28030 18174 28082
rect 18226 28030 18228 28082
rect 18172 28018 18228 28030
rect 18060 27972 18116 27982
rect 18060 27878 18116 27916
rect 17948 26786 18004 26796
rect 18060 26964 18116 26974
rect 18060 26404 18116 26908
rect 18284 26516 18340 30828
rect 18620 30882 18676 30894
rect 20748 30884 20804 30894
rect 18620 30830 18622 30882
rect 18674 30830 18676 30882
rect 18620 29650 18676 30830
rect 20188 30882 20804 30884
rect 20188 30830 20750 30882
rect 20802 30830 20804 30882
rect 20188 30828 20804 30830
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 18620 29598 18622 29650
rect 18674 29598 18676 29650
rect 18620 29540 18676 29598
rect 18956 29652 19012 29662
rect 19628 29652 19684 29662
rect 20188 29652 20244 30828
rect 20748 30818 20804 30828
rect 20300 29988 20356 29998
rect 20300 29894 20356 29932
rect 18956 29650 19684 29652
rect 18956 29598 18958 29650
rect 19010 29598 19630 29650
rect 19682 29598 19684 29650
rect 18956 29596 19684 29598
rect 18956 29586 19012 29596
rect 19628 29586 19684 29596
rect 19964 29596 20244 29652
rect 18620 29474 18676 29484
rect 19852 29538 19908 29550
rect 19852 29486 19854 29538
rect 19906 29486 19908 29538
rect 18844 29426 18900 29438
rect 18844 29374 18846 29426
rect 18898 29374 18900 29426
rect 18396 28756 18452 28766
rect 18396 28662 18452 28700
rect 18508 28644 18564 28654
rect 18564 28588 18676 28644
rect 18508 28578 18564 28588
rect 18284 26450 18340 26460
rect 18508 26852 18564 26862
rect 18060 26338 18116 26348
rect 18172 26292 18228 26302
rect 18172 26198 18228 26236
rect 18508 26290 18564 26796
rect 18508 26238 18510 26290
rect 18562 26238 18564 26290
rect 18508 26226 18564 26238
rect 17612 26124 17892 26180
rect 17612 26068 17668 26124
rect 17500 26012 17668 26068
rect 17500 25506 17556 26012
rect 17500 25454 17502 25506
rect 17554 25454 17556 25506
rect 17500 25442 17556 25454
rect 17612 25730 17668 25742
rect 17612 25678 17614 25730
rect 17666 25678 17668 25730
rect 17164 25396 17220 25406
rect 17164 25302 17220 25340
rect 16940 24052 16996 24062
rect 16828 24050 16996 24052
rect 16828 23998 16942 24050
rect 16994 23998 16996 24050
rect 16828 23996 16996 23998
rect 16940 23986 16996 23996
rect 17164 23938 17220 23950
rect 17164 23886 17166 23938
rect 17218 23886 17220 23938
rect 16044 22990 16046 23042
rect 16098 22990 16100 23042
rect 15372 21810 15428 22316
rect 15708 22596 15764 22606
rect 15708 22258 15764 22540
rect 15932 22484 15988 22494
rect 15932 22390 15988 22428
rect 15708 22206 15710 22258
rect 15762 22206 15764 22258
rect 15708 22194 15764 22206
rect 15372 21758 15374 21810
rect 15426 21758 15428 21810
rect 15372 21746 15428 21758
rect 15148 20804 15204 20814
rect 15148 20802 15540 20804
rect 15148 20750 15150 20802
rect 15202 20750 15540 20802
rect 15148 20748 15540 20750
rect 15148 20738 15204 20748
rect 15036 20692 15092 20702
rect 15036 20598 15092 20636
rect 15484 20242 15540 20748
rect 15484 20190 15486 20242
rect 15538 20190 15540 20242
rect 15484 20178 15540 20190
rect 14588 19926 14644 19964
rect 14812 20132 14868 20142
rect 14812 20130 15204 20132
rect 14812 20078 14814 20130
rect 14866 20078 15204 20130
rect 14812 20076 15204 20078
rect 14252 18676 14308 18686
rect 14252 18582 14308 18620
rect 14700 18674 14756 18686
rect 14700 18622 14702 18674
rect 14754 18622 14756 18674
rect 14476 18564 14532 18574
rect 14476 18470 14532 18508
rect 14364 18452 14420 18462
rect 14364 18358 14420 18396
rect 14476 18004 14532 18014
rect 14476 17780 14532 17948
rect 14476 17714 14532 17724
rect 14700 17778 14756 18622
rect 14812 18676 14868 20076
rect 15148 19458 15204 20076
rect 16044 20130 16100 22990
rect 16268 23826 16324 23838
rect 16268 23774 16270 23826
rect 16322 23774 16324 23826
rect 16156 22596 16212 22606
rect 16268 22596 16324 23774
rect 17164 22596 17220 23886
rect 17612 23828 17668 25678
rect 18172 25396 18228 25406
rect 18172 25302 18228 25340
rect 18620 25060 18676 28588
rect 18844 28532 18900 29374
rect 19068 29426 19124 29438
rect 19068 29374 19070 29426
rect 19122 29374 19124 29426
rect 19068 29316 19124 29374
rect 19292 29428 19348 29438
rect 19292 29334 19348 29372
rect 19068 29250 19124 29260
rect 19852 29092 19908 29486
rect 19964 29314 20020 29596
rect 20300 29316 20356 29326
rect 19964 29262 19966 29314
rect 20018 29262 20020 29314
rect 19964 29250 20020 29262
rect 20076 29314 20356 29316
rect 20076 29262 20302 29314
rect 20354 29262 20356 29314
rect 20076 29260 20356 29262
rect 20076 29092 20132 29260
rect 19852 29036 20132 29092
rect 18844 27748 18900 28476
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 18844 27692 19124 27748
rect 18844 26964 18900 26974
rect 18844 26514 18900 26908
rect 18844 26462 18846 26514
rect 18898 26462 18900 26514
rect 18844 26450 18900 26462
rect 18732 26290 18788 26302
rect 18732 26238 18734 26290
rect 18786 26238 18788 26290
rect 18732 26068 18788 26238
rect 18956 26292 19012 26302
rect 18956 26198 19012 26236
rect 18732 25284 18788 26012
rect 18732 25218 18788 25228
rect 18620 25004 19012 25060
rect 18956 24946 19012 25004
rect 18956 24894 18958 24946
rect 19010 24894 19012 24946
rect 18956 23940 19012 24894
rect 17724 23828 17780 23838
rect 17612 23826 17780 23828
rect 17612 23774 17726 23826
rect 17778 23774 17780 23826
rect 17612 23772 17780 23774
rect 17500 23156 17556 23166
rect 17612 23156 17668 23772
rect 17724 23762 17780 23772
rect 17500 23154 17668 23156
rect 17500 23102 17502 23154
rect 17554 23102 17668 23154
rect 17500 23100 17668 23102
rect 17500 23090 17556 23100
rect 16156 22594 16324 22596
rect 16156 22542 16158 22594
rect 16210 22542 16324 22594
rect 16156 22540 16324 22542
rect 16940 22540 17164 22596
rect 16156 20914 16212 22540
rect 16156 20862 16158 20914
rect 16210 20862 16212 20914
rect 16156 20850 16212 20862
rect 16940 20914 16996 22540
rect 17164 22530 17220 22540
rect 17276 23044 17332 23054
rect 17164 22372 17220 22382
rect 17276 22372 17332 22988
rect 17220 22316 17332 22372
rect 17948 23042 18004 23054
rect 17948 22990 17950 23042
rect 18002 22990 18004 23042
rect 17164 22278 17220 22316
rect 17052 22260 17108 22270
rect 17052 22166 17108 22204
rect 16940 20862 16942 20914
rect 16994 20862 16996 20914
rect 16940 20850 16996 20862
rect 17052 21812 17108 21822
rect 17052 20802 17108 21756
rect 17052 20750 17054 20802
rect 17106 20750 17108 20802
rect 17052 20738 17108 20750
rect 17276 20690 17332 20702
rect 17276 20638 17278 20690
rect 17330 20638 17332 20690
rect 17276 20188 17332 20638
rect 16044 20078 16046 20130
rect 16098 20078 16100 20130
rect 16044 20066 16100 20078
rect 16940 20132 17332 20188
rect 15148 19406 15150 19458
rect 15202 19406 15204 19458
rect 15148 19394 15204 19406
rect 15820 20018 15876 20030
rect 15820 19966 15822 20018
rect 15874 19966 15876 20018
rect 15036 19124 15092 19134
rect 14812 18562 14868 18620
rect 14812 18510 14814 18562
rect 14866 18510 14868 18562
rect 14812 18498 14868 18510
rect 14924 19122 15092 19124
rect 14924 19070 15038 19122
rect 15090 19070 15092 19122
rect 14924 19068 15092 19070
rect 14924 17892 14980 19068
rect 15036 19058 15092 19068
rect 15036 18564 15092 18574
rect 15036 18450 15092 18508
rect 15036 18398 15038 18450
rect 15090 18398 15092 18450
rect 15036 18386 15092 18398
rect 15484 18450 15540 18462
rect 15484 18398 15486 18450
rect 15538 18398 15540 18450
rect 15260 18228 15316 18238
rect 15260 18134 15316 18172
rect 15036 17892 15092 17902
rect 14924 17836 15036 17892
rect 15036 17826 15092 17836
rect 14700 17726 14702 17778
rect 14754 17726 14756 17778
rect 14700 17714 14756 17726
rect 15484 17668 15540 18398
rect 15708 18452 15764 18462
rect 15708 18358 15764 18396
rect 15484 17602 15540 17612
rect 15260 16884 15316 16894
rect 15708 16884 15764 16894
rect 15260 16882 15764 16884
rect 15260 16830 15262 16882
rect 15314 16830 15710 16882
rect 15762 16830 15764 16882
rect 15260 16828 15764 16830
rect 15260 16818 15316 16828
rect 15708 16098 15764 16828
rect 15708 16046 15710 16098
rect 15762 16046 15764 16098
rect 15708 15876 15764 16046
rect 15708 15810 15764 15820
rect 13468 15092 13748 15148
rect 14140 15092 15092 15148
rect 13692 13972 13748 15092
rect 14252 14420 14308 14430
rect 13692 13746 13748 13916
rect 13692 13694 13694 13746
rect 13746 13694 13748 13746
rect 13692 13682 13748 13694
rect 14028 14418 14308 14420
rect 14028 14366 14254 14418
rect 14306 14366 14308 14418
rect 14028 14364 14308 14366
rect 14028 12852 14084 14364
rect 14252 14354 14308 14364
rect 14364 14418 14420 15092
rect 15036 14644 15092 15092
rect 15148 14644 15204 14654
rect 15036 14642 15764 14644
rect 15036 14590 15150 14642
rect 15202 14590 15764 14642
rect 15036 14588 15764 14590
rect 15148 14578 15204 14588
rect 14364 14366 14366 14418
rect 14418 14366 14420 14418
rect 14364 14354 14420 14366
rect 15484 14420 15540 14430
rect 15540 14364 15652 14420
rect 15484 14326 15540 14364
rect 14588 14308 14644 14318
rect 14588 14306 14980 14308
rect 14588 14254 14590 14306
rect 14642 14254 14980 14306
rect 14588 14252 14980 14254
rect 14588 14242 14644 14252
rect 14252 13972 14308 13982
rect 14252 13970 14644 13972
rect 14252 13918 14254 13970
rect 14306 13918 14644 13970
rect 14252 13916 14644 13918
rect 14252 13906 14308 13916
rect 14140 13746 14196 13758
rect 14140 13694 14142 13746
rect 14194 13694 14196 13746
rect 14140 13636 14196 13694
rect 14364 13748 14420 13758
rect 14364 13654 14420 13692
rect 14588 13746 14644 13916
rect 14924 13858 14980 14252
rect 14924 13806 14926 13858
rect 14978 13806 14980 13858
rect 14924 13794 14980 13806
rect 15596 13858 15652 14364
rect 15596 13806 15598 13858
rect 15650 13806 15652 13858
rect 14588 13694 14590 13746
rect 14642 13694 14644 13746
rect 14588 13682 14644 13694
rect 15036 13748 15092 13758
rect 15372 13748 15428 13758
rect 15092 13746 15428 13748
rect 15092 13694 15374 13746
rect 15426 13694 15428 13746
rect 15092 13692 15428 13694
rect 14140 13570 14196 13580
rect 14924 13636 14980 13646
rect 14924 12962 14980 13580
rect 15036 13074 15092 13692
rect 15372 13682 15428 13692
rect 15484 13634 15540 13646
rect 15484 13582 15486 13634
rect 15538 13582 15540 13634
rect 15148 13524 15204 13534
rect 15372 13524 15428 13534
rect 15148 13522 15372 13524
rect 15148 13470 15150 13522
rect 15202 13470 15372 13522
rect 15148 13468 15372 13470
rect 15148 13458 15204 13468
rect 15372 13458 15428 13468
rect 15036 13022 15038 13074
rect 15090 13022 15092 13074
rect 15036 13010 15092 13022
rect 15484 13076 15540 13582
rect 15596 13636 15652 13806
rect 15596 13570 15652 13580
rect 15484 13010 15540 13020
rect 15708 13074 15764 14588
rect 15820 14420 15876 19966
rect 16156 18338 16212 18350
rect 16156 18286 16158 18338
rect 16210 18286 16212 18338
rect 16156 18228 16212 18286
rect 15820 14354 15876 14364
rect 16044 18172 16156 18228
rect 16044 13970 16100 18172
rect 16156 18162 16212 18172
rect 16828 17892 16884 17902
rect 16828 17778 16884 17836
rect 16828 17726 16830 17778
rect 16882 17726 16884 17778
rect 16828 17714 16884 17726
rect 16044 13918 16046 13970
rect 16098 13918 16100 13970
rect 16044 13524 16100 13918
rect 16044 13458 16100 13468
rect 15708 13022 15710 13074
rect 15762 13022 15764 13074
rect 15708 13010 15764 13022
rect 14924 12910 14926 12962
rect 14978 12910 14980 12962
rect 14924 12898 14980 12910
rect 14084 12796 14196 12852
rect 14028 12786 14084 12796
rect 13356 12338 13412 12348
rect 13916 11508 13972 11518
rect 13244 10610 13300 10780
rect 13580 11506 13972 11508
rect 13580 11454 13918 11506
rect 13970 11454 13972 11506
rect 13580 11452 13972 11454
rect 13244 10558 13246 10610
rect 13298 10558 13300 10610
rect 13244 10546 13300 10558
rect 13468 10612 13524 10622
rect 12236 9884 12740 9940
rect 12236 9826 12292 9884
rect 12236 9774 12238 9826
rect 12290 9774 12292 9826
rect 12236 9762 12292 9774
rect 12348 9716 12404 9726
rect 12572 9716 12628 9726
rect 12348 9622 12404 9660
rect 12460 9660 12572 9716
rect 12460 9602 12516 9660
rect 12572 9650 12628 9660
rect 12460 9550 12462 9602
rect 12514 9550 12516 9602
rect 12460 9538 12516 9550
rect 12124 9324 12516 9380
rect 12460 9266 12516 9324
rect 12460 9214 12462 9266
rect 12514 9214 12516 9266
rect 12460 9202 12516 9214
rect 12684 9266 12740 9884
rect 12908 9938 12964 10108
rect 12908 9886 12910 9938
rect 12962 9886 12964 9938
rect 12908 9874 12964 9886
rect 12684 9214 12686 9266
rect 12738 9214 12740 9266
rect 12684 9202 12740 9214
rect 12796 9716 12852 9726
rect 12796 9154 12852 9660
rect 12796 9102 12798 9154
rect 12850 9102 12852 9154
rect 12796 9090 12852 9102
rect 13468 8146 13524 10556
rect 13580 10610 13636 11452
rect 13916 11442 13972 11452
rect 14028 11394 14084 11406
rect 14028 11342 14030 11394
rect 14082 11342 14084 11394
rect 13916 11284 13972 11294
rect 13916 11190 13972 11228
rect 14028 10948 14084 11342
rect 14140 11284 14196 12796
rect 14588 12850 14644 12862
rect 14588 12798 14590 12850
rect 14642 12798 14644 12850
rect 14252 11676 14532 11732
rect 14252 11394 14308 11676
rect 14252 11342 14254 11394
rect 14306 11342 14308 11394
rect 14252 11330 14308 11342
rect 14364 11508 14420 11518
rect 14364 11394 14420 11452
rect 14364 11342 14366 11394
rect 14418 11342 14420 11394
rect 14364 11330 14420 11342
rect 14140 11218 14196 11228
rect 14028 10892 14420 10948
rect 13916 10780 14196 10836
rect 13804 10724 13860 10734
rect 13916 10724 13972 10780
rect 13804 10722 13972 10724
rect 13804 10670 13806 10722
rect 13858 10670 13972 10722
rect 13804 10668 13972 10670
rect 13804 10658 13860 10668
rect 13580 10558 13582 10610
rect 13634 10558 13636 10610
rect 13580 10546 13636 10558
rect 14028 10610 14084 10622
rect 14028 10558 14030 10610
rect 14082 10558 14084 10610
rect 13916 10498 13972 10510
rect 13916 10446 13918 10498
rect 13970 10446 13972 10498
rect 13804 9940 13860 9950
rect 13804 9826 13860 9884
rect 13804 9774 13806 9826
rect 13858 9774 13860 9826
rect 13804 9762 13860 9774
rect 13916 8428 13972 10446
rect 14028 9940 14084 10558
rect 14028 9874 14084 9884
rect 14140 9940 14196 10780
rect 14364 10834 14420 10892
rect 14364 10782 14366 10834
rect 14418 10782 14420 10834
rect 14364 10052 14420 10782
rect 14476 10498 14532 11676
rect 14588 10948 14644 12798
rect 14924 11508 14980 11518
rect 14924 11414 14980 11452
rect 14588 10892 14980 10948
rect 14588 10612 14644 10622
rect 14588 10518 14644 10556
rect 14924 10610 14980 10892
rect 15260 10836 15316 10846
rect 15260 10742 15316 10780
rect 14924 10558 14926 10610
rect 14978 10558 14980 10610
rect 14476 10446 14478 10498
rect 14530 10446 14532 10498
rect 14476 10434 14532 10446
rect 14924 10388 14980 10558
rect 14924 10322 14980 10332
rect 14364 9996 15092 10052
rect 14140 9884 14980 9940
rect 14140 9826 14196 9884
rect 14140 9774 14142 9826
rect 14194 9774 14196 9826
rect 14140 9762 14196 9774
rect 14924 9826 14980 9884
rect 14924 9774 14926 9826
rect 14978 9774 14980 9826
rect 14924 9762 14980 9774
rect 15036 9938 15092 9996
rect 15036 9886 15038 9938
rect 15090 9886 15092 9938
rect 13468 8094 13470 8146
rect 13522 8094 13524 8146
rect 13468 8082 13524 8094
rect 13580 8372 13972 8428
rect 14588 9714 14644 9726
rect 14588 9662 14590 9714
rect 14642 9662 14644 9714
rect 10892 5966 10894 6018
rect 10946 5966 10948 6018
rect 10892 5954 10948 5966
rect 13020 6804 13076 6814
rect 10556 5842 10612 5852
rect 13020 5794 13076 6748
rect 13468 5908 13524 5918
rect 13468 5814 13524 5852
rect 13020 5742 13022 5794
rect 13074 5742 13076 5794
rect 13020 5730 13076 5742
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 13580 5012 13636 8372
rect 14588 8148 14644 9662
rect 15036 8428 15092 9886
rect 15820 9828 15876 9838
rect 14588 8082 14644 8092
rect 14812 8372 15316 8428
rect 13804 8034 13860 8046
rect 13804 7982 13806 8034
rect 13858 7982 13860 8034
rect 13804 6804 13860 7982
rect 13804 6738 13860 6748
rect 14812 6578 14868 8372
rect 15260 8370 15316 8372
rect 15260 8318 15262 8370
rect 15314 8318 15316 8370
rect 15260 8306 15316 8318
rect 15820 8370 15876 9772
rect 15820 8318 15822 8370
rect 15874 8318 15876 8370
rect 15820 8306 15876 8318
rect 15484 8258 15540 8270
rect 15484 8206 15486 8258
rect 15538 8206 15540 8258
rect 15484 6804 15540 8206
rect 15484 6738 15540 6748
rect 16044 6804 16100 6814
rect 14812 6526 14814 6578
rect 14866 6526 14868 6578
rect 14812 6514 14868 6526
rect 15148 6580 15204 6590
rect 15148 6578 15316 6580
rect 15148 6526 15150 6578
rect 15202 6526 15316 6578
rect 15148 6524 15316 6526
rect 15148 6514 15204 6524
rect 13132 4956 13636 5012
rect 15260 5124 15316 6524
rect 13132 4450 13188 4956
rect 13132 4398 13134 4450
rect 13186 4398 13188 4450
rect 13132 4386 13188 4398
rect 12460 4340 12516 4350
rect 12460 4246 12516 4284
rect 15260 4226 15316 5068
rect 15932 5124 15988 5134
rect 15932 5030 15988 5068
rect 16044 5010 16100 6748
rect 16044 4958 16046 5010
rect 16098 4958 16100 5010
rect 16044 4946 16100 4958
rect 16940 4898 16996 20132
rect 17836 19348 17892 19358
rect 17836 19254 17892 19292
rect 17948 18004 18004 22990
rect 18844 22596 18900 22606
rect 18844 22260 18900 22540
rect 18956 22372 19012 23884
rect 19068 23378 19124 27692
rect 20188 27076 20244 29260
rect 20300 29250 20356 29260
rect 20636 27300 20692 27310
rect 20300 27188 20356 27198
rect 20636 27188 20692 27244
rect 20300 27186 20692 27188
rect 20300 27134 20302 27186
rect 20354 27134 20692 27186
rect 20300 27132 20692 27134
rect 20300 27122 20356 27132
rect 20188 27010 20244 27020
rect 20524 26964 20580 26974
rect 20524 26870 20580 26908
rect 20636 26962 20692 27132
rect 20636 26910 20638 26962
rect 20690 26910 20692 26962
rect 20636 26898 20692 26910
rect 20860 26852 20916 26862
rect 20860 26850 21028 26852
rect 20860 26798 20862 26850
rect 20914 26798 21028 26850
rect 20860 26796 21028 26798
rect 20860 26786 20916 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19852 26516 19908 26526
rect 19852 26422 19908 26460
rect 19180 26404 19236 26414
rect 19180 26290 19236 26348
rect 20972 26402 21028 26796
rect 20972 26350 20974 26402
rect 21026 26350 21028 26402
rect 20972 26338 21028 26350
rect 19180 26238 19182 26290
rect 19234 26238 19236 26290
rect 19180 23716 19236 26238
rect 20188 26292 20244 26302
rect 20188 26198 20244 26236
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 21084 24052 21140 31892
rect 21420 30996 21476 31006
rect 21420 30902 21476 30940
rect 21868 27748 21924 34636
rect 24332 32786 24388 35420
rect 25564 34804 25620 36428
rect 25788 36370 25844 36428
rect 25788 36318 25790 36370
rect 25842 36318 25844 36370
rect 25788 36306 25844 36318
rect 26348 36370 26404 36428
rect 26460 36482 26516 36652
rect 28700 36708 28756 37102
rect 28700 36642 28756 36652
rect 26460 36430 26462 36482
rect 26514 36430 26516 36482
rect 26460 36418 26516 36430
rect 26348 36318 26350 36370
rect 26402 36318 26404 36370
rect 26348 36306 26404 36318
rect 25676 36258 25732 36270
rect 25676 36206 25678 36258
rect 25730 36206 25732 36258
rect 25676 34916 25732 36206
rect 26124 36260 26180 36270
rect 26124 36258 26292 36260
rect 26124 36206 26126 36258
rect 26178 36206 26292 36258
rect 26124 36204 26292 36206
rect 26124 36194 26180 36204
rect 25900 35698 25956 35710
rect 25900 35646 25902 35698
rect 25954 35646 25956 35698
rect 25900 35026 25956 35646
rect 25900 34974 25902 35026
rect 25954 34974 25956 35026
rect 25900 34962 25956 34974
rect 25788 34916 25844 34926
rect 25676 34914 25844 34916
rect 25676 34862 25790 34914
rect 25842 34862 25844 34914
rect 25676 34860 25844 34862
rect 25788 34850 25844 34860
rect 26012 34916 26068 34926
rect 26012 34822 26068 34860
rect 25564 34748 25732 34804
rect 24332 32734 24334 32786
rect 24386 32734 24388 32786
rect 24332 32722 24388 32734
rect 24220 32674 24276 32686
rect 24668 32676 24724 32686
rect 24220 32622 24222 32674
rect 24274 32622 24276 32674
rect 24220 32564 24276 32622
rect 24220 32498 24276 32508
rect 24556 32620 24668 32676
rect 24444 32340 24500 32350
rect 24220 32338 24500 32340
rect 24220 32286 24446 32338
rect 24498 32286 24500 32338
rect 24220 32284 24500 32286
rect 24108 31668 24164 31678
rect 24108 31574 24164 31612
rect 24220 31218 24276 32284
rect 24444 32274 24500 32284
rect 24556 32116 24612 32620
rect 24668 32610 24724 32620
rect 25228 32676 25284 32686
rect 25228 32582 25284 32620
rect 25340 32564 25396 32574
rect 25340 32470 25396 32508
rect 25452 32562 25508 32574
rect 25452 32510 25454 32562
rect 25506 32510 25508 32562
rect 25452 32340 25508 32510
rect 24444 32060 24612 32116
rect 25116 32284 25452 32340
rect 24444 31666 24500 32060
rect 25116 31948 25172 32284
rect 25452 32246 25508 32284
rect 25676 32562 25732 34748
rect 26236 34802 26292 36204
rect 26236 34750 26238 34802
rect 26290 34750 26292 34802
rect 26236 34738 26292 34750
rect 26908 35810 26964 35822
rect 26908 35758 26910 35810
rect 26962 35758 26964 35810
rect 25676 32510 25678 32562
rect 25730 32510 25732 32562
rect 25676 31948 25732 32510
rect 24892 31892 24948 31902
rect 24444 31614 24446 31666
rect 24498 31614 24500 31666
rect 24444 31602 24500 31614
rect 24556 31890 24948 31892
rect 24556 31838 24894 31890
rect 24946 31838 24948 31890
rect 24556 31836 24948 31838
rect 24220 31166 24222 31218
rect 24274 31166 24276 31218
rect 24220 31154 24276 31166
rect 24444 31106 24500 31118
rect 24444 31054 24446 31106
rect 24498 31054 24500 31106
rect 23996 30884 24052 30894
rect 24444 30884 24500 31054
rect 23996 30882 24500 30884
rect 23996 30830 23998 30882
rect 24050 30830 24500 30882
rect 23996 30828 24500 30830
rect 24556 31106 24612 31836
rect 24892 31826 24948 31836
rect 25004 31892 25172 31948
rect 25228 31892 25732 31948
rect 25004 31778 25060 31892
rect 25004 31726 25006 31778
rect 25058 31726 25060 31778
rect 25004 31714 25060 31726
rect 24780 31668 24836 31678
rect 24556 31054 24558 31106
rect 24610 31054 24612 31106
rect 23548 29316 23604 29326
rect 23548 28754 23604 29260
rect 23548 28702 23550 28754
rect 23602 28702 23604 28754
rect 23548 28690 23604 28702
rect 23996 28980 24052 30828
rect 24556 30322 24612 31054
rect 24556 30270 24558 30322
rect 24610 30270 24612 30322
rect 24556 30258 24612 30270
rect 24668 31612 24780 31668
rect 22876 28644 22932 28654
rect 22876 28550 22932 28588
rect 21868 27746 22036 27748
rect 21868 27694 21870 27746
rect 21922 27694 22036 27746
rect 21868 27692 22036 27694
rect 21868 27682 21924 27692
rect 21756 27186 21812 27198
rect 21756 27134 21758 27186
rect 21810 27134 21812 27186
rect 21756 27076 21812 27134
rect 21980 27188 22036 27692
rect 21980 27122 22036 27132
rect 22540 27188 22596 27198
rect 21756 27010 21812 27020
rect 22540 27074 22596 27132
rect 22540 27022 22542 27074
rect 22594 27022 22596 27074
rect 22540 27010 22596 27022
rect 21084 23986 21140 23996
rect 21308 26964 21364 26974
rect 19292 23940 19348 23950
rect 19292 23846 19348 23884
rect 19628 23716 19684 23726
rect 19180 23714 19684 23716
rect 19180 23662 19630 23714
rect 19682 23662 19684 23714
rect 19180 23660 19684 23662
rect 19068 23326 19070 23378
rect 19122 23326 19124 23378
rect 19068 23314 19124 23326
rect 19180 23266 19236 23278
rect 19180 23214 19182 23266
rect 19234 23214 19236 23266
rect 19180 22820 19236 23214
rect 19180 22754 19236 22764
rect 19404 23154 19460 23166
rect 19404 23102 19406 23154
rect 19458 23102 19460 23154
rect 19404 22596 19460 23102
rect 19404 22502 19460 22540
rect 19068 22372 19124 22382
rect 18956 22370 19124 22372
rect 18956 22318 19070 22370
rect 19122 22318 19124 22370
rect 18956 22316 19124 22318
rect 19068 22306 19124 22316
rect 18844 21698 18900 22204
rect 18844 21646 18846 21698
rect 18898 21646 18900 21698
rect 18844 21634 18900 21646
rect 19068 21700 19124 21710
rect 19068 21606 19124 21644
rect 18956 21474 19012 21486
rect 18956 21422 18958 21474
rect 19010 21422 19012 21474
rect 17948 17938 18004 17948
rect 18060 20690 18116 20702
rect 18060 20638 18062 20690
rect 18114 20638 18116 20690
rect 17500 17892 17556 17902
rect 17276 17668 17332 17678
rect 17332 17612 17444 17668
rect 17276 17602 17332 17612
rect 17276 17444 17332 17454
rect 17276 16884 17332 17388
rect 17276 16818 17332 16828
rect 17388 16660 17444 17612
rect 17500 17106 17556 17836
rect 17500 17054 17502 17106
rect 17554 17054 17556 17106
rect 17500 17042 17556 17054
rect 17612 16882 17668 16894
rect 17612 16830 17614 16882
rect 17666 16830 17668 16882
rect 17500 16660 17556 16670
rect 17388 16658 17556 16660
rect 17388 16606 17502 16658
rect 17554 16606 17556 16658
rect 17388 16604 17556 16606
rect 17500 16594 17556 16604
rect 17612 15540 17668 16830
rect 17612 15474 17668 15484
rect 18060 15204 18116 20638
rect 18060 15138 18116 15148
rect 18396 16884 18452 16894
rect 18396 15986 18452 16828
rect 18956 16100 19012 21422
rect 19516 20188 19572 23660
rect 19628 23650 19684 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20188 23492 20244 23502
rect 19852 23156 19908 23166
rect 19628 23100 19852 23156
rect 19628 22482 19684 23100
rect 19852 23062 19908 23100
rect 20188 23154 20244 23436
rect 20188 23102 20190 23154
rect 20242 23102 20244 23154
rect 20188 23090 20244 23102
rect 20412 23380 20468 23390
rect 20412 23154 20468 23324
rect 21084 23266 21140 23278
rect 21084 23214 21086 23266
rect 21138 23214 21140 23266
rect 20412 23102 20414 23154
rect 20466 23102 20468 23154
rect 20412 23090 20468 23102
rect 20748 23156 20804 23166
rect 20748 23062 20804 23100
rect 19628 22430 19630 22482
rect 19682 22430 19684 22482
rect 19628 22418 19684 22430
rect 19740 22820 19796 22830
rect 19740 22148 19796 22764
rect 21084 22820 21140 23214
rect 21084 22754 21140 22764
rect 19180 20132 19572 20188
rect 19628 22092 19796 22148
rect 19628 20188 19684 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 21308 20188 21364 26908
rect 22204 26964 22260 26974
rect 22204 26870 22260 26908
rect 22876 26180 22932 26190
rect 21532 25508 21588 25518
rect 21532 23380 21588 25452
rect 22764 25396 22820 25406
rect 22764 23826 22820 25340
rect 22764 23774 22766 23826
rect 22818 23774 22820 23826
rect 21532 23286 21588 23324
rect 22540 23714 22596 23726
rect 22540 23662 22542 23714
rect 22594 23662 22596 23714
rect 21532 22372 21588 22382
rect 21756 22372 21812 22382
rect 21532 22370 21812 22372
rect 21532 22318 21534 22370
rect 21586 22318 21758 22370
rect 21810 22318 21812 22370
rect 21532 22316 21812 22318
rect 21532 22148 21588 22316
rect 21756 22306 21812 22316
rect 21532 22082 21588 22092
rect 19628 20132 19796 20188
rect 19068 20020 19124 20030
rect 19068 18564 19124 19964
rect 19068 18470 19124 18508
rect 19180 18228 19236 20132
rect 19740 20020 19796 20132
rect 20412 20132 21364 20188
rect 19740 19926 19796 19964
rect 19964 20018 20020 20030
rect 19964 19966 19966 20018
rect 20018 19966 20020 20018
rect 19852 19906 19908 19918
rect 19852 19854 19854 19906
rect 19906 19854 19908 19906
rect 19852 19236 19908 19854
rect 19964 19572 20020 19966
rect 20412 20018 20468 20132
rect 20412 19966 20414 20018
rect 20466 19966 20468 20018
rect 19964 19516 20356 19572
rect 19404 19180 19908 19236
rect 20188 19348 20244 19358
rect 19292 18452 19348 18462
rect 19404 18452 19460 19180
rect 19964 19122 20020 19134
rect 19964 19070 19966 19122
rect 20018 19070 20020 19122
rect 19964 19012 20020 19070
rect 19628 18956 20020 19012
rect 19516 18676 19572 18686
rect 19628 18676 19684 18956
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19516 18674 19684 18676
rect 19516 18622 19518 18674
rect 19570 18622 19684 18674
rect 19516 18620 19684 18622
rect 20188 18674 20244 19292
rect 20188 18622 20190 18674
rect 20242 18622 20244 18674
rect 19516 18610 19572 18620
rect 20188 18610 20244 18622
rect 19628 18452 19684 18462
rect 19404 18450 19684 18452
rect 19404 18398 19630 18450
rect 19682 18398 19684 18450
rect 19404 18396 19684 18398
rect 19292 18358 19348 18396
rect 19628 18386 19684 18396
rect 20188 18452 20244 18462
rect 20300 18452 20356 19516
rect 20244 18396 20356 18452
rect 20188 18386 20244 18396
rect 19516 18228 19572 18238
rect 20300 18228 20356 18238
rect 19180 18226 19572 18228
rect 19180 18174 19518 18226
rect 19570 18174 19572 18226
rect 19180 18172 19572 18174
rect 19516 18162 19572 18172
rect 20188 18172 20300 18228
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20188 16882 20244 18172
rect 20300 18162 20356 18172
rect 20188 16830 20190 16882
rect 20242 16830 20244 16882
rect 20188 16818 20244 16830
rect 20412 16660 20468 19966
rect 20636 19234 20692 19246
rect 20636 19182 20638 19234
rect 20690 19182 20692 19234
rect 20636 19012 20692 19182
rect 21420 19012 21476 19022
rect 20636 19010 21476 19012
rect 20636 18958 21422 19010
rect 21474 18958 21476 19010
rect 20636 18956 21476 18958
rect 20636 16884 20692 18956
rect 21420 18946 21476 18956
rect 20748 18452 20804 18462
rect 20748 18358 20804 18396
rect 20636 16818 20692 16828
rect 20748 16882 20804 16894
rect 20748 16830 20750 16882
rect 20802 16830 20804 16882
rect 20748 16660 20804 16830
rect 20412 16604 20804 16660
rect 18956 16034 19012 16044
rect 18396 15934 18398 15986
rect 18450 15934 18452 15986
rect 18396 14644 18452 15934
rect 19964 15876 20020 15914
rect 19964 15810 20020 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19516 15540 19572 15550
rect 18396 14588 18564 14644
rect 17836 13076 17892 13086
rect 17836 12982 17892 13020
rect 18508 12964 18564 14588
rect 18620 12964 18676 12974
rect 18508 12962 18676 12964
rect 18508 12910 18622 12962
rect 18674 12910 18676 12962
rect 18508 12908 18676 12910
rect 18620 12740 18676 12908
rect 19068 12740 19124 12750
rect 18620 12738 19124 12740
rect 18620 12686 19070 12738
rect 19122 12686 19124 12738
rect 18620 12684 19124 12686
rect 17276 10724 17332 10734
rect 17276 10050 17332 10668
rect 18284 10500 18340 10510
rect 18284 10406 18340 10444
rect 17276 9998 17278 10050
rect 17330 9998 17332 10050
rect 17276 9986 17332 9998
rect 17836 10052 17892 10062
rect 17500 9828 17556 9838
rect 17500 9734 17556 9772
rect 17836 9714 17892 9996
rect 18732 9938 18788 9950
rect 18732 9886 18734 9938
rect 18786 9886 18788 9938
rect 18284 9826 18340 9838
rect 18284 9774 18286 9826
rect 18338 9774 18340 9826
rect 17836 9662 17838 9714
rect 17890 9662 17892 9714
rect 17836 9650 17892 9662
rect 18172 9714 18228 9726
rect 18172 9662 18174 9714
rect 18226 9662 18228 9714
rect 17612 9042 17668 9054
rect 17612 8990 17614 9042
rect 17666 8990 17668 9042
rect 17612 8428 17668 8990
rect 17836 9044 17892 9054
rect 17836 8950 17892 8988
rect 18060 9042 18116 9054
rect 18060 8990 18062 9042
rect 18114 8990 18116 9042
rect 17948 8930 18004 8942
rect 17948 8878 17950 8930
rect 18002 8878 18004 8930
rect 17612 8372 17892 8428
rect 17836 8036 17892 8372
rect 17836 7942 17892 7980
rect 16940 4846 16942 4898
rect 16994 4846 16996 4898
rect 16940 4834 16996 4846
rect 17388 6132 17444 6142
rect 17388 5906 17444 6076
rect 17948 6020 18004 8878
rect 18060 8258 18116 8990
rect 18060 8206 18062 8258
rect 18114 8206 18116 8258
rect 18060 8194 18116 8206
rect 18172 7812 18228 9662
rect 18284 9268 18340 9774
rect 18732 9604 18788 9886
rect 18284 9202 18340 9212
rect 18396 9548 18788 9604
rect 18844 9714 18900 9726
rect 18844 9662 18846 9714
rect 18898 9662 18900 9714
rect 18396 9042 18452 9548
rect 18732 9380 18788 9390
rect 18620 9324 18732 9380
rect 18620 9266 18676 9324
rect 18732 9314 18788 9324
rect 18620 9214 18622 9266
rect 18674 9214 18676 9266
rect 18620 9202 18676 9214
rect 18844 9266 18900 9662
rect 18844 9214 18846 9266
rect 18898 9214 18900 9266
rect 18396 8990 18398 9042
rect 18450 8990 18452 9042
rect 18396 8932 18452 8990
rect 18508 9044 18564 9054
rect 18508 8950 18564 8988
rect 18396 8258 18452 8876
rect 18844 8428 18900 9214
rect 18396 8206 18398 8258
rect 18450 8206 18452 8258
rect 18396 8194 18452 8206
rect 18732 8372 18900 8428
rect 18284 8148 18340 8158
rect 18284 8054 18340 8092
rect 18732 8034 18788 8372
rect 18956 8370 19012 8382
rect 18956 8318 18958 8370
rect 19010 8318 19012 8370
rect 18956 8260 19012 8318
rect 18956 8194 19012 8204
rect 18732 7982 18734 8034
rect 18786 7982 18788 8034
rect 18732 7812 18788 7982
rect 18844 8148 18900 8158
rect 18844 8036 18900 8092
rect 18956 8036 19012 8046
rect 18844 8034 19012 8036
rect 18844 7982 18958 8034
rect 19010 7982 19012 8034
rect 18844 7980 19012 7982
rect 18956 7970 19012 7980
rect 18172 7756 18788 7812
rect 18284 6578 18340 7756
rect 18284 6526 18286 6578
rect 18338 6526 18340 6578
rect 18284 6514 18340 6526
rect 18620 6466 18676 6478
rect 18620 6414 18622 6466
rect 18674 6414 18676 6466
rect 18172 6020 18228 6030
rect 17948 6018 18228 6020
rect 17948 5966 18174 6018
rect 18226 5966 18228 6018
rect 17948 5964 18228 5966
rect 18172 5954 18228 5964
rect 17388 5854 17390 5906
rect 17442 5854 17444 5906
rect 15708 4340 15764 4350
rect 15708 4246 15764 4284
rect 17388 4340 17444 5854
rect 18620 5796 18676 6414
rect 19068 6132 19124 12684
rect 19180 9826 19236 9838
rect 19180 9774 19182 9826
rect 19234 9774 19236 9826
rect 19180 8148 19236 9774
rect 19292 9604 19348 9614
rect 19292 8258 19348 9548
rect 19516 9492 19572 15484
rect 19852 15540 19908 15550
rect 19852 15446 19908 15484
rect 19628 15314 19684 15326
rect 19628 15262 19630 15314
rect 19682 15262 19684 15314
rect 19628 15092 19684 15262
rect 20748 15314 20804 16604
rect 20748 15262 20750 15314
rect 20802 15262 20804 15314
rect 20748 15250 20804 15262
rect 20412 15202 20468 15214
rect 20412 15150 20414 15202
rect 20466 15150 20468 15202
rect 19628 15026 19684 15036
rect 20076 15092 20132 15102
rect 20076 14642 20132 15036
rect 20076 14590 20078 14642
rect 20130 14590 20132 14642
rect 20076 14578 20132 14590
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20412 13636 20468 15150
rect 21868 15092 21924 15102
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19628 11396 19684 11406
rect 19628 10500 19684 11340
rect 20412 11172 20468 13580
rect 20412 11106 20468 11116
rect 20524 14532 20580 14542
rect 20524 12178 20580 14476
rect 21084 13076 21140 13086
rect 20748 12404 20804 12414
rect 20748 12310 20804 12348
rect 21084 12290 21140 13020
rect 21868 13076 21924 15036
rect 22540 15092 22596 23662
rect 22652 23380 22708 23390
rect 22652 23286 22708 23324
rect 22764 23268 22820 23774
rect 22876 25284 22932 26124
rect 23100 26178 23156 26190
rect 23100 26126 23102 26178
rect 23154 26126 23156 26178
rect 23100 26068 23156 26126
rect 23100 26002 23156 26012
rect 22876 23938 22932 25228
rect 23436 24052 23492 24062
rect 23436 23958 23492 23996
rect 23884 24052 23940 24062
rect 23884 23958 23940 23996
rect 22876 23886 22878 23938
rect 22930 23886 22932 23938
rect 22876 23492 22932 23886
rect 22876 23426 22932 23436
rect 23548 23380 23604 23390
rect 22764 23212 23380 23268
rect 23324 23154 23380 23212
rect 23324 23102 23326 23154
rect 23378 23102 23380 23154
rect 23324 23090 23380 23102
rect 23548 23154 23604 23324
rect 23548 23102 23550 23154
rect 23602 23102 23604 23154
rect 23548 23090 23604 23102
rect 23884 23044 23940 23054
rect 23884 22950 23940 22988
rect 22988 22930 23044 22942
rect 22988 22878 22990 22930
rect 23042 22878 23044 22930
rect 22988 20188 23044 22878
rect 23996 20188 24052 28924
rect 24220 25508 24276 25518
rect 24220 25414 24276 25452
rect 24444 25396 24500 25406
rect 24668 25396 24724 31612
rect 24780 31574 24836 31612
rect 25228 31666 25284 31892
rect 25228 31614 25230 31666
rect 25282 31614 25284 31666
rect 25228 31602 25284 31614
rect 24892 30212 24948 30222
rect 24892 30118 24948 30156
rect 25676 30212 25732 30222
rect 25340 30098 25396 30110
rect 25340 30046 25342 30098
rect 25394 30046 25396 30098
rect 25228 29540 25284 29550
rect 25340 29540 25396 30046
rect 25228 29538 25396 29540
rect 25228 29486 25230 29538
rect 25282 29486 25396 29538
rect 25228 29484 25396 29486
rect 25228 29474 25284 29484
rect 25564 29426 25620 29438
rect 25564 29374 25566 29426
rect 25618 29374 25620 29426
rect 25340 29316 25396 29326
rect 25340 29222 25396 29260
rect 25564 29316 25620 29374
rect 25564 29250 25620 29260
rect 25676 28754 25732 30156
rect 26908 30212 26964 35758
rect 27356 35588 27412 35598
rect 27356 35494 27412 35532
rect 29036 35028 29092 35038
rect 28140 34914 28196 34926
rect 28140 34862 28142 34914
rect 28194 34862 28196 34914
rect 27468 34802 27524 34814
rect 27468 34750 27470 34802
rect 27522 34750 27524 34802
rect 27468 34020 27524 34750
rect 27468 33954 27524 33964
rect 27356 33124 27412 33134
rect 27356 30882 27412 33068
rect 27356 30830 27358 30882
rect 27410 30830 27412 30882
rect 27356 30818 27412 30830
rect 28140 32340 28196 34862
rect 28364 34916 28420 34926
rect 28364 34822 28420 34860
rect 29036 34914 29092 34972
rect 29036 34862 29038 34914
rect 29090 34862 29092 34914
rect 29036 34850 29092 34862
rect 29372 34916 29428 34926
rect 29372 34822 29428 34860
rect 29260 34690 29316 34702
rect 29260 34638 29262 34690
rect 29314 34638 29316 34690
rect 29260 33348 29316 34638
rect 29372 33348 29428 33358
rect 29260 33346 29428 33348
rect 29260 33294 29374 33346
rect 29426 33294 29428 33346
rect 29260 33292 29428 33294
rect 26908 30146 26964 30156
rect 28140 30210 28196 32284
rect 29148 33122 29204 33134
rect 29148 33070 29150 33122
rect 29202 33070 29204 33122
rect 29148 32340 29204 33070
rect 29372 33124 29428 33292
rect 29372 33058 29428 33068
rect 29148 32274 29204 32284
rect 30268 30994 30324 39564
rect 30940 39620 30996 39630
rect 30940 39526 30996 39564
rect 31948 39620 32004 40350
rect 33740 39730 33796 41916
rect 36092 41860 36148 45200
rect 36316 41972 36372 41982
rect 36316 41878 36372 41916
rect 36092 41794 36148 41804
rect 37324 41860 37380 41870
rect 37324 41766 37380 41804
rect 39900 41860 39956 45200
rect 39900 41794 39956 41804
rect 40124 41970 40180 41982
rect 40124 41918 40126 41970
rect 40178 41918 40180 41970
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 39788 40964 39844 40974
rect 40124 40964 40180 41918
rect 41132 41860 41188 41870
rect 41132 41766 41188 41804
rect 43148 41412 43204 41422
rect 43708 41412 43764 45200
rect 43148 41410 43764 41412
rect 43148 41358 43150 41410
rect 43202 41358 43764 41410
rect 43148 41356 43764 41358
rect 43148 41346 43204 41356
rect 39788 40962 40180 40964
rect 39788 40910 39790 40962
rect 39842 40910 40180 40962
rect 39788 40908 40180 40910
rect 43932 41186 43988 41198
rect 43932 41134 43934 41186
rect 43986 41134 43988 41186
rect 37436 40402 37492 40414
rect 37436 40350 37438 40402
rect 37490 40350 37492 40402
rect 34636 40292 34692 40302
rect 36764 40292 36820 40302
rect 34636 40290 34804 40292
rect 34636 40238 34638 40290
rect 34690 40238 34804 40290
rect 34636 40236 34804 40238
rect 34636 40226 34692 40236
rect 33740 39678 33742 39730
rect 33794 39678 33796 39730
rect 33740 39666 33796 39678
rect 31948 39554 32004 39564
rect 34188 39620 34244 39630
rect 34188 39526 34244 39564
rect 31948 38162 32004 38174
rect 31948 38110 31950 38162
rect 32002 38110 32004 38162
rect 31612 37268 31668 37278
rect 31612 37174 31668 37212
rect 30828 37154 30884 37166
rect 30828 37102 30830 37154
rect 30882 37102 30884 37154
rect 30828 36596 30884 37102
rect 30828 36530 30884 36540
rect 31948 34916 32004 38110
rect 34076 37940 34132 37950
rect 34076 37938 34580 37940
rect 34076 37886 34078 37938
rect 34130 37886 34580 37938
rect 34076 37884 34580 37886
rect 34076 37874 34132 37884
rect 32060 37268 32116 37278
rect 32060 37174 32116 37212
rect 34412 37156 34468 37166
rect 34076 37154 34468 37156
rect 34076 37102 34414 37154
rect 34466 37102 34468 37154
rect 34076 37100 34468 37102
rect 34076 36820 34132 37100
rect 34412 37090 34468 37100
rect 33628 36764 34132 36820
rect 32284 36708 32340 36718
rect 32284 36594 32340 36652
rect 32284 36542 32286 36594
rect 32338 36542 32340 36594
rect 32284 36530 32340 36542
rect 33516 36708 33572 36718
rect 33516 36370 33572 36652
rect 33516 36318 33518 36370
rect 33570 36318 33572 36370
rect 33516 36306 33572 36318
rect 32396 36260 32452 36270
rect 32396 36166 32452 36204
rect 31948 34850 32004 34860
rect 33628 33460 33684 36764
rect 33852 36596 33908 36606
rect 33852 36502 33908 36540
rect 34076 36482 34132 36764
rect 34076 36430 34078 36482
rect 34130 36430 34132 36482
rect 34076 36418 34132 36430
rect 34412 36932 34468 36942
rect 34412 36482 34468 36876
rect 34524 36594 34580 37884
rect 34524 36542 34526 36594
rect 34578 36542 34580 36594
rect 34524 36530 34580 36542
rect 34412 36430 34414 36482
rect 34466 36430 34468 36482
rect 33740 36370 33796 36382
rect 33740 36318 33742 36370
rect 33794 36318 33796 36370
rect 33740 36036 33796 36318
rect 33852 36260 33908 36270
rect 33852 36166 33908 36204
rect 34412 36148 34468 36430
rect 34636 36482 34692 36494
rect 34636 36430 34638 36482
rect 34690 36430 34692 36482
rect 34636 36260 34692 36430
rect 34636 36194 34692 36204
rect 34412 36092 34580 36148
rect 33740 35980 34468 36036
rect 34412 35922 34468 35980
rect 34412 35870 34414 35922
rect 34466 35870 34468 35922
rect 34412 35858 34468 35870
rect 34524 35476 34580 36092
rect 34748 36036 34804 40236
rect 36764 40290 37156 40292
rect 36764 40238 36766 40290
rect 36818 40238 37156 40290
rect 36764 40236 37156 40238
rect 36764 40226 36820 40236
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 37100 38162 37156 40236
rect 37100 38110 37102 38162
rect 37154 38110 37156 38162
rect 37100 38098 37156 38110
rect 37436 39396 37492 40350
rect 38108 40404 38164 40414
rect 38108 40290 38164 40348
rect 38108 40238 38110 40290
rect 38162 40238 38164 40290
rect 37884 39620 37940 39630
rect 38108 39620 38164 40238
rect 37884 39618 38164 39620
rect 37884 39566 37886 39618
rect 37938 39566 38164 39618
rect 37884 39564 38164 39566
rect 37548 39396 37604 39406
rect 37884 39396 37940 39564
rect 37436 39394 37940 39396
rect 37436 39342 37550 39394
rect 37602 39342 37940 39394
rect 37436 39340 37940 39342
rect 38668 39506 38724 39518
rect 38668 39454 38670 39506
rect 38722 39454 38724 39506
rect 34860 38050 34916 38062
rect 34860 37998 34862 38050
rect 34914 37998 34916 38050
rect 34860 37828 34916 37998
rect 36988 37940 37044 37950
rect 35308 37828 35364 37838
rect 34860 37772 35308 37828
rect 35308 37268 35364 37772
rect 35308 37044 35364 37212
rect 36988 37044 37044 37884
rect 37324 37938 37380 37950
rect 37324 37886 37326 37938
rect 37378 37886 37380 37938
rect 37324 37492 37380 37886
rect 37436 37828 37492 39340
rect 37548 39330 37604 39340
rect 37436 37762 37492 37772
rect 37548 37938 37604 37950
rect 37548 37886 37550 37938
rect 37602 37886 37604 37938
rect 37324 37426 37380 37436
rect 35308 36988 35588 37044
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35420 36708 35476 36718
rect 35420 36594 35476 36652
rect 35420 36542 35422 36594
rect 35474 36542 35476 36594
rect 35420 36530 35476 36542
rect 34972 36372 35028 36382
rect 34972 36278 35028 36316
rect 34636 35980 34804 36036
rect 34636 35810 34692 35980
rect 34636 35758 34638 35810
rect 34690 35758 34692 35810
rect 34636 35588 34692 35758
rect 34636 35522 34692 35532
rect 34748 35698 34804 35710
rect 34748 35646 34750 35698
rect 34802 35646 34804 35698
rect 34412 35420 34580 35476
rect 33628 33458 34020 33460
rect 33628 33406 33630 33458
rect 33682 33406 34020 33458
rect 33628 33404 34020 33406
rect 33628 33394 33684 33404
rect 32284 33348 32340 33358
rect 32284 32676 32340 33292
rect 33180 33348 33236 33358
rect 33180 33254 33236 33292
rect 32284 32562 32340 32620
rect 32508 32676 32564 32686
rect 32508 32582 32564 32620
rect 32284 32510 32286 32562
rect 32338 32510 32340 32562
rect 32284 32498 32340 32510
rect 33180 32564 33236 32574
rect 33516 32564 33572 32574
rect 33180 32562 33516 32564
rect 33180 32510 33182 32562
rect 33234 32510 33516 32562
rect 33180 32508 33516 32510
rect 33180 32498 33236 32508
rect 33404 32228 33460 32238
rect 33292 31892 33348 31902
rect 32956 31668 33012 31678
rect 33292 31668 33348 31836
rect 33404 31890 33460 32172
rect 33516 31948 33572 32508
rect 33852 32450 33908 32462
rect 33852 32398 33854 32450
rect 33906 32398 33908 32450
rect 33852 32228 33908 32398
rect 33852 32162 33908 32172
rect 33964 31948 34020 33404
rect 34076 33348 34132 33358
rect 34076 33254 34132 33292
rect 34412 33234 34468 35420
rect 34748 33796 34804 35646
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35084 34916 35140 34926
rect 35084 34822 35140 34860
rect 34412 33182 34414 33234
rect 34466 33182 34468 33234
rect 34300 32676 34356 32686
rect 33516 31892 33684 31948
rect 33964 31892 34132 31948
rect 33404 31838 33406 31890
rect 33458 31838 33460 31890
rect 33404 31826 33460 31838
rect 30268 30942 30270 30994
rect 30322 30942 30324 30994
rect 29484 30882 29540 30894
rect 29484 30830 29486 30882
rect 29538 30830 29540 30882
rect 28140 30158 28142 30210
rect 28194 30158 28196 30210
rect 28140 30146 28196 30158
rect 28364 30210 28420 30222
rect 28364 30158 28366 30210
rect 28418 30158 28420 30210
rect 26236 29988 26292 29998
rect 26012 29316 26068 29326
rect 26012 29222 26068 29260
rect 25676 28702 25678 28754
rect 25730 28702 25732 28754
rect 25676 28690 25732 28702
rect 26124 28644 26180 28654
rect 26124 28550 26180 28588
rect 25452 27188 25508 27198
rect 25452 27094 25508 27132
rect 25900 27188 25956 27198
rect 25900 27074 25956 27132
rect 25900 27022 25902 27074
rect 25954 27022 25956 27074
rect 25900 27010 25956 27022
rect 24892 25508 24948 25518
rect 24892 25414 24948 25452
rect 24500 25340 24724 25396
rect 24444 25302 24500 25340
rect 24332 24052 24388 24062
rect 24332 23938 24388 23996
rect 24332 23886 24334 23938
rect 24386 23886 24388 23938
rect 24332 23874 24388 23886
rect 24892 24052 24948 24062
rect 24892 23938 24948 23996
rect 24892 23886 24894 23938
rect 24946 23886 24948 23938
rect 24892 23874 24948 23886
rect 24556 23716 24612 23726
rect 24444 23714 24612 23716
rect 24444 23662 24558 23714
rect 24610 23662 24612 23714
rect 24444 23660 24612 23662
rect 24444 23156 24500 23660
rect 24556 23650 24612 23660
rect 25228 23714 25284 23726
rect 25228 23662 25230 23714
rect 25282 23662 25284 23714
rect 24444 23062 24500 23100
rect 24668 21812 24724 21822
rect 25228 21812 25284 23662
rect 26012 23492 26068 23502
rect 25564 23156 25620 23166
rect 25676 23156 25732 23166
rect 25564 23154 25676 23156
rect 25564 23102 25566 23154
rect 25618 23102 25676 23154
rect 25564 23100 25676 23102
rect 25564 23090 25620 23100
rect 25564 22484 25620 22494
rect 24668 21810 25228 21812
rect 24668 21758 24670 21810
rect 24722 21758 25228 21810
rect 24668 21756 25228 21758
rect 24668 21746 24724 21756
rect 22876 20132 23044 20188
rect 23884 20132 24052 20188
rect 22652 18338 22708 18350
rect 22652 18286 22654 18338
rect 22706 18286 22708 18338
rect 22652 18228 22708 18286
rect 22876 18228 22932 20132
rect 23212 18564 23268 18574
rect 23212 18470 23268 18508
rect 23436 18564 23492 18574
rect 23436 18470 23492 18508
rect 22988 18452 23044 18462
rect 23548 18452 23604 18462
rect 22988 18450 23156 18452
rect 22988 18398 22990 18450
rect 23042 18398 23156 18450
rect 22988 18396 23156 18398
rect 22988 18386 23044 18396
rect 22876 18172 23044 18228
rect 22652 18162 22708 18172
rect 22876 18004 22932 18014
rect 22876 17778 22932 17948
rect 22876 17726 22878 17778
rect 22930 17726 22932 17778
rect 22876 17668 22932 17726
rect 22540 15026 22596 15036
rect 22764 17612 22876 17668
rect 21868 12982 21924 13020
rect 22652 12628 22708 12638
rect 22204 12404 22260 12414
rect 21084 12238 21086 12290
rect 21138 12238 21140 12290
rect 21084 12226 21140 12238
rect 21980 12348 22204 12404
rect 20524 12126 20526 12178
rect 20578 12126 20580 12178
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 20524 10724 20580 12126
rect 21644 12180 21700 12190
rect 21644 12066 21700 12124
rect 21644 12014 21646 12066
rect 21698 12014 21700 12066
rect 21644 12002 21700 12014
rect 21308 11956 21364 11966
rect 21308 11862 21364 11900
rect 21756 11396 21812 11406
rect 21756 11302 21812 11340
rect 21980 11394 22036 12348
rect 22204 12310 22260 12348
rect 22652 12292 22708 12572
rect 22540 12290 22708 12292
rect 22540 12238 22654 12290
rect 22706 12238 22708 12290
rect 22540 12236 22708 12238
rect 22092 12178 22148 12190
rect 22092 12126 22094 12178
rect 22146 12126 22148 12178
rect 22092 11956 22148 12126
rect 22428 12180 22484 12190
rect 22428 12086 22484 12124
rect 22092 11508 22148 11900
rect 22316 12066 22372 12078
rect 22316 12014 22318 12066
rect 22370 12014 22372 12066
rect 22204 11508 22260 11518
rect 22092 11506 22260 11508
rect 22092 11454 22206 11506
rect 22258 11454 22260 11506
rect 22092 11452 22260 11454
rect 22204 11442 22260 11452
rect 21980 11342 21982 11394
rect 22034 11342 22036 11394
rect 21980 11330 22036 11342
rect 20524 10658 20580 10668
rect 19740 10500 19796 10510
rect 19684 10498 19796 10500
rect 19684 10446 19742 10498
rect 19794 10446 19796 10498
rect 19684 10444 19796 10446
rect 19628 10052 19684 10444
rect 19740 10434 19796 10444
rect 19628 9826 19684 9996
rect 20412 10052 20468 10062
rect 20412 9958 20468 9996
rect 19628 9774 19630 9826
rect 19682 9774 19684 9826
rect 19628 9762 19684 9774
rect 20188 9602 20244 9614
rect 20188 9550 20190 9602
rect 20242 9550 20244 9602
rect 19516 9436 19684 9492
rect 19628 9380 19684 9436
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19516 9268 19572 9278
rect 19628 9268 19684 9324
rect 19852 9268 19908 9278
rect 19628 9266 19908 9268
rect 19628 9214 19854 9266
rect 19906 9214 19908 9266
rect 19628 9212 19908 9214
rect 19516 8428 19572 9212
rect 19852 9202 19908 9212
rect 20076 9268 20132 9278
rect 20076 9156 20132 9212
rect 20188 9156 20244 9550
rect 20300 9604 20356 9614
rect 20300 9510 20356 9548
rect 20076 9154 20244 9156
rect 20076 9102 20078 9154
rect 20130 9102 20244 9154
rect 20076 9100 20244 9102
rect 20076 9062 20132 9100
rect 19628 9042 19684 9054
rect 19628 8990 19630 9042
rect 19682 8990 19684 9042
rect 19628 8932 19684 8990
rect 19628 8866 19684 8876
rect 19740 8930 19796 8942
rect 19740 8878 19742 8930
rect 19794 8878 19796 8930
rect 19740 8428 19796 8878
rect 22316 8428 22372 12014
rect 22428 11396 22484 11406
rect 22540 11396 22596 12236
rect 22652 12226 22708 12236
rect 22428 11394 22596 11396
rect 22428 11342 22430 11394
rect 22482 11342 22596 11394
rect 22428 11340 22596 11342
rect 22652 11396 22708 11406
rect 22764 11396 22820 17612
rect 22876 17602 22932 17612
rect 22988 15876 23044 18172
rect 23100 16324 23156 18396
rect 23548 18358 23604 18396
rect 23884 18450 23940 20132
rect 24780 19348 24836 19358
rect 24108 19236 24164 19246
rect 24108 19234 24276 19236
rect 24108 19182 24110 19234
rect 24162 19182 24276 19234
rect 24108 19180 24276 19182
rect 24108 19170 24164 19180
rect 24220 18788 24276 19180
rect 24780 19234 24836 19292
rect 24780 19182 24782 19234
rect 24834 19182 24836 19234
rect 24780 19170 24836 19182
rect 24332 19124 24388 19134
rect 24332 19030 24388 19068
rect 24220 18732 24612 18788
rect 24556 18674 24612 18732
rect 24556 18622 24558 18674
rect 24610 18622 24612 18674
rect 24556 18610 24612 18622
rect 24444 18564 24500 18574
rect 23884 18398 23886 18450
rect 23938 18398 23940 18450
rect 23884 18228 23940 18398
rect 23884 18162 23940 18172
rect 23996 18450 24052 18462
rect 23996 18398 23998 18450
rect 24050 18398 24052 18450
rect 23996 18004 24052 18398
rect 24108 18452 24164 18462
rect 24108 18358 24164 18396
rect 23324 17948 24052 18004
rect 23324 17778 23380 17948
rect 23324 17726 23326 17778
rect 23378 17726 23380 17778
rect 23324 17714 23380 17726
rect 24444 17778 24500 18508
rect 24444 17726 24446 17778
rect 24498 17726 24500 17778
rect 24444 17714 24500 17726
rect 23436 17668 23492 17678
rect 23436 17574 23492 17612
rect 23884 17668 23940 17678
rect 24332 17668 24388 17678
rect 23884 17666 24388 17668
rect 23884 17614 23886 17666
rect 23938 17614 24334 17666
rect 24386 17614 24388 17666
rect 23884 17612 24388 17614
rect 23884 17602 23940 17612
rect 24332 17602 24388 17612
rect 23100 16258 23156 16268
rect 23212 17554 23268 17566
rect 23212 17502 23214 17554
rect 23266 17502 23268 17554
rect 23212 16100 23268 17502
rect 23436 16324 23492 16334
rect 23436 16230 23492 16268
rect 23996 16324 24052 16334
rect 23324 16100 23380 16110
rect 23212 16098 23604 16100
rect 23212 16046 23326 16098
rect 23378 16046 23604 16098
rect 23212 16044 23604 16046
rect 23324 16034 23380 16044
rect 23436 15876 23492 15886
rect 22876 15874 23492 15876
rect 22876 15822 22990 15874
rect 23042 15822 23438 15874
rect 23490 15822 23492 15874
rect 22876 15820 23492 15822
rect 22876 12740 22932 15820
rect 22988 15810 23044 15820
rect 23436 15810 23492 15820
rect 23548 15652 23604 16044
rect 23436 15596 23604 15652
rect 23212 15428 23268 15438
rect 23212 15334 23268 15372
rect 23324 15426 23380 15438
rect 23324 15374 23326 15426
rect 23378 15374 23380 15426
rect 23324 14980 23380 15374
rect 23212 14924 23380 14980
rect 23212 14644 23268 14924
rect 23324 14756 23380 14766
rect 23436 14756 23492 15596
rect 23548 15428 23604 15438
rect 23548 15426 23716 15428
rect 23548 15374 23550 15426
rect 23602 15374 23716 15426
rect 23548 15372 23716 15374
rect 23548 15362 23604 15372
rect 23660 15314 23716 15372
rect 23996 15426 24052 16268
rect 25004 15988 25060 21756
rect 25228 21718 25284 21756
rect 25340 22428 25564 22484
rect 25228 21474 25284 21486
rect 25228 21422 25230 21474
rect 25282 21422 25284 21474
rect 25228 21364 25284 21422
rect 25228 21298 25284 21308
rect 25228 20802 25284 20814
rect 25228 20750 25230 20802
rect 25282 20750 25284 20802
rect 25228 19012 25284 20750
rect 25228 18340 25284 18956
rect 25228 18274 25284 18284
rect 24220 15652 24276 15662
rect 23996 15374 23998 15426
rect 24050 15374 24052 15426
rect 23996 15362 24052 15374
rect 24108 15596 24220 15652
rect 23660 15262 23662 15314
rect 23714 15262 23716 15314
rect 23660 15250 23716 15262
rect 24108 14756 24164 15596
rect 24220 15586 24276 15596
rect 24220 15316 24276 15326
rect 24220 15222 24276 15260
rect 24668 15314 24724 15326
rect 24668 15262 24670 15314
rect 24722 15262 24724 15314
rect 24444 15204 24500 15214
rect 23324 14754 23492 14756
rect 23324 14702 23326 14754
rect 23378 14702 23492 14754
rect 23324 14700 23492 14702
rect 23548 14700 24164 14756
rect 23324 14690 23380 14700
rect 23212 14578 23268 14588
rect 22988 14532 23044 14542
rect 22988 14438 23044 14476
rect 23436 12964 23492 12974
rect 23100 12962 23492 12964
rect 23100 12910 23438 12962
rect 23490 12910 23492 12962
rect 23100 12908 23492 12910
rect 22988 12740 23044 12750
rect 22876 12684 22988 12740
rect 22988 12674 23044 12684
rect 23100 12404 23156 12908
rect 23436 12898 23492 12908
rect 23100 12178 23156 12348
rect 23100 12126 23102 12178
rect 23154 12126 23156 12178
rect 23100 12114 23156 12126
rect 23212 12740 23268 12750
rect 23212 12178 23268 12684
rect 23212 12126 23214 12178
rect 23266 12126 23268 12178
rect 23212 11508 23268 12126
rect 23212 11442 23268 11452
rect 23436 12628 23492 12638
rect 23436 12402 23492 12572
rect 23436 12350 23438 12402
rect 23490 12350 23492 12402
rect 22708 11340 22820 11396
rect 22428 11330 22484 11340
rect 22652 11302 22708 11340
rect 23436 11282 23492 12350
rect 23548 11396 23604 14700
rect 23660 14532 23716 14542
rect 23660 14530 24052 14532
rect 23660 14478 23662 14530
rect 23714 14478 24052 14530
rect 23660 14476 24052 14478
rect 23660 14466 23716 14476
rect 23996 12850 24052 14476
rect 24108 14420 24164 14700
rect 24332 15202 24500 15204
rect 24332 15150 24446 15202
rect 24498 15150 24500 15202
rect 24332 15148 24500 15150
rect 24220 14420 24276 14430
rect 24108 14418 24276 14420
rect 24108 14366 24222 14418
rect 24274 14366 24276 14418
rect 24108 14364 24276 14366
rect 24220 14354 24276 14364
rect 24332 13972 24388 15148
rect 24444 15138 24500 15148
rect 24556 15202 24612 15214
rect 24556 15150 24558 15202
rect 24610 15150 24612 15202
rect 24444 14644 24500 14654
rect 24444 14530 24500 14588
rect 24444 14478 24446 14530
rect 24498 14478 24500 14530
rect 24444 14466 24500 14478
rect 24108 13916 24388 13972
rect 24108 13186 24164 13916
rect 24556 13860 24612 15150
rect 24668 14756 24724 15262
rect 24668 14690 24724 14700
rect 25004 15316 25060 15932
rect 25340 15876 25396 22428
rect 25564 22418 25620 22428
rect 25676 20802 25732 23100
rect 26012 23154 26068 23436
rect 26012 23102 26014 23154
rect 26066 23102 26068 23154
rect 25788 21812 25844 21822
rect 25788 21718 25844 21756
rect 25676 20750 25678 20802
rect 25730 20750 25732 20802
rect 25676 20738 25732 20750
rect 25900 21364 25956 21374
rect 25452 19124 25508 19134
rect 25452 19030 25508 19068
rect 25340 15810 25396 15820
rect 25788 15652 25844 15662
rect 25340 15540 25396 15550
rect 25340 15446 25396 15484
rect 25788 15426 25844 15596
rect 25788 15374 25790 15426
rect 25842 15374 25844 15426
rect 25788 15362 25844 15374
rect 25004 14642 25060 15260
rect 25228 15316 25284 15326
rect 25228 15314 25732 15316
rect 25228 15262 25230 15314
rect 25282 15262 25732 15314
rect 25228 15260 25732 15262
rect 25228 15250 25284 15260
rect 25452 14756 25508 14766
rect 25452 14662 25508 14700
rect 25004 14590 25006 14642
rect 25058 14590 25060 14642
rect 25004 14578 25060 14590
rect 25564 14644 25620 14654
rect 25564 14550 25620 14588
rect 24556 13794 24612 13804
rect 24108 13134 24110 13186
rect 24162 13134 24164 13186
rect 24108 13122 24164 13134
rect 25676 12964 25732 15260
rect 23996 12798 23998 12850
rect 24050 12798 24052 12850
rect 23772 12738 23828 12750
rect 23772 12686 23774 12738
rect 23826 12686 23828 12738
rect 23772 12628 23828 12686
rect 23772 12562 23828 12572
rect 23884 12404 23940 12414
rect 23660 12348 23884 12404
rect 23996 12404 24052 12798
rect 25228 12962 25732 12964
rect 25228 12910 25678 12962
rect 25730 12910 25732 12962
rect 25228 12908 25732 12910
rect 24444 12740 24500 12750
rect 24444 12646 24500 12684
rect 24556 12404 24612 12414
rect 23996 12348 24164 12404
rect 23660 12290 23716 12348
rect 23884 12338 23940 12348
rect 23660 12238 23662 12290
rect 23714 12238 23716 12290
rect 23660 12226 23716 12238
rect 24108 12292 24164 12348
rect 24556 12310 24612 12348
rect 24108 12198 24164 12236
rect 24668 12292 24724 12302
rect 24668 12198 24724 12236
rect 23996 12180 24052 12190
rect 23996 12086 24052 12124
rect 24332 12178 24388 12190
rect 24332 12126 24334 12178
rect 24386 12126 24388 12178
rect 23772 12068 23828 12078
rect 23772 12066 23940 12068
rect 23772 12014 23774 12066
rect 23826 12014 23940 12066
rect 23772 12012 23940 12014
rect 23772 12002 23828 12012
rect 23660 11396 23716 11406
rect 23548 11394 23716 11396
rect 23548 11342 23662 11394
rect 23714 11342 23716 11394
rect 23548 11340 23716 11342
rect 23884 11396 23940 12012
rect 23996 11396 24052 11406
rect 23884 11394 24052 11396
rect 23884 11342 23998 11394
rect 24050 11342 24052 11394
rect 23884 11340 24052 11342
rect 23436 11230 23438 11282
rect 23490 11230 23492 11282
rect 23436 11218 23492 11230
rect 23660 8428 23716 11340
rect 23996 11330 24052 11340
rect 24332 11394 24388 12126
rect 25228 11506 25284 12908
rect 25676 12898 25732 12908
rect 25452 12738 25508 12750
rect 25452 12686 25454 12738
rect 25506 12686 25508 12738
rect 25452 12292 25508 12686
rect 25452 12226 25508 12236
rect 25900 11956 25956 21308
rect 26012 17556 26068 23102
rect 26236 22484 26292 29932
rect 28364 29650 28420 30158
rect 29372 30210 29428 30222
rect 29372 30158 29374 30210
rect 29426 30158 29428 30210
rect 28588 30100 28644 30110
rect 28588 30098 29204 30100
rect 28588 30046 28590 30098
rect 28642 30046 29204 30098
rect 28588 30044 29204 30046
rect 28588 30034 28644 30044
rect 28364 29598 28366 29650
rect 28418 29598 28420 29650
rect 26684 29316 26740 29326
rect 26348 27412 26404 27422
rect 26348 27188 26404 27356
rect 26348 27186 26516 27188
rect 26348 27134 26350 27186
rect 26402 27134 26516 27186
rect 26348 27132 26516 27134
rect 26348 27122 26404 27132
rect 26348 23156 26404 23166
rect 26348 23062 26404 23100
rect 26236 22390 26292 22428
rect 26236 21812 26292 21822
rect 26012 17490 26068 17500
rect 26124 21474 26180 21486
rect 26124 21422 26126 21474
rect 26178 21422 26180 21474
rect 26124 17780 26180 21422
rect 26236 20914 26292 21756
rect 26236 20862 26238 20914
rect 26290 20862 26292 20914
rect 26236 20850 26292 20862
rect 25228 11454 25230 11506
rect 25282 11454 25284 11506
rect 25228 11442 25284 11454
rect 25340 11900 25956 11956
rect 24332 11342 24334 11394
rect 24386 11342 24388 11394
rect 24332 11330 24388 11342
rect 24668 11396 24724 11406
rect 24668 11302 24724 11340
rect 25340 11396 25396 11900
rect 24220 11284 24276 11294
rect 24220 11190 24276 11228
rect 25340 10836 25396 11340
rect 25116 10834 25396 10836
rect 25116 10782 25342 10834
rect 25394 10782 25396 10834
rect 25116 10780 25396 10782
rect 19516 8372 19684 8428
rect 19740 8372 20132 8428
rect 19292 8206 19294 8258
rect 19346 8206 19348 8258
rect 19292 8194 19348 8206
rect 19180 8082 19236 8092
rect 19068 6066 19124 6076
rect 18620 5730 18676 5740
rect 17388 4274 17444 4284
rect 19628 5010 19684 8372
rect 19852 8260 19908 8270
rect 19852 8166 19908 8204
rect 20076 8258 20132 8372
rect 20076 8206 20078 8258
rect 20130 8206 20132 8258
rect 20076 8194 20132 8206
rect 20412 8372 20468 8382
rect 20412 8258 20468 8316
rect 21420 8372 21476 8382
rect 22316 8372 23156 8428
rect 23660 8372 24724 8428
rect 21420 8278 21476 8316
rect 23100 8370 23156 8372
rect 23100 8318 23102 8370
rect 23154 8318 23156 8370
rect 23100 8306 23156 8318
rect 20412 8206 20414 8258
rect 20466 8206 20468 8258
rect 20412 8194 20468 8206
rect 23436 8258 23492 8270
rect 23436 8206 23438 8258
rect 23490 8206 23492 8258
rect 20076 8036 20132 8046
rect 23212 8036 23268 8046
rect 20076 8034 20244 8036
rect 20076 7982 20078 8034
rect 20130 7982 20244 8034
rect 20076 7980 20244 7982
rect 20076 7970 20132 7980
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 20188 7700 20244 7980
rect 20076 7644 20244 7700
rect 22540 8034 23268 8036
rect 22540 7982 23214 8034
rect 23266 7982 23268 8034
rect 22540 7980 23268 7982
rect 20076 6468 20132 7644
rect 22540 7586 22596 7980
rect 23212 7970 23268 7980
rect 23436 8036 23492 8206
rect 23436 7970 23492 7980
rect 23884 8036 23940 8046
rect 23884 7942 23940 7980
rect 22540 7534 22542 7586
rect 22594 7534 22596 7586
rect 22540 7522 22596 7534
rect 24556 7700 24612 7710
rect 21868 7474 21924 7486
rect 21868 7422 21870 7474
rect 21922 7422 21924 7474
rect 21868 6804 21924 7422
rect 21868 6738 21924 6748
rect 22988 6804 23044 6814
rect 20076 6402 20132 6412
rect 21756 6468 21812 6478
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20748 6132 20804 6142
rect 20748 6038 20804 6076
rect 20300 5796 20356 5806
rect 19740 5124 19796 5134
rect 20300 5124 20356 5740
rect 19740 5122 20356 5124
rect 19740 5070 19742 5122
rect 19794 5070 20356 5122
rect 19740 5068 20356 5070
rect 19740 5058 19796 5068
rect 19628 4958 19630 5010
rect 19682 4958 19684 5010
rect 15260 4174 15262 4226
rect 15314 4174 15316 4226
rect 15260 4162 15316 4174
rect 19628 4226 19684 4958
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 21756 4450 21812 6412
rect 22988 4564 23044 6748
rect 24556 6804 24612 7644
rect 24668 7362 24724 8372
rect 25116 8372 25172 10780
rect 25340 10770 25396 10780
rect 26124 8428 26180 17724
rect 26460 9604 26516 27132
rect 26684 23378 26740 29260
rect 28252 28532 28308 28542
rect 27132 27076 27188 27086
rect 26796 26290 26852 26302
rect 26796 26238 26798 26290
rect 26850 26238 26852 26290
rect 26796 26180 26852 26238
rect 26796 26114 26852 26124
rect 27132 25618 27188 27020
rect 28252 27076 28308 28476
rect 27468 26180 27524 26190
rect 27468 26178 27636 26180
rect 27468 26126 27470 26178
rect 27522 26126 27636 26178
rect 27468 26124 27636 26126
rect 27468 26114 27524 26124
rect 27132 25566 27134 25618
rect 27186 25566 27188 25618
rect 27132 25554 27188 25566
rect 27580 25618 27636 26124
rect 27580 25566 27582 25618
rect 27634 25566 27636 25618
rect 27580 25554 27636 25566
rect 28252 25506 28308 27020
rect 28364 26964 28420 29598
rect 28588 29652 28644 29662
rect 28588 28868 28644 29596
rect 29148 29538 29204 30044
rect 29372 29988 29428 30158
rect 29372 29922 29428 29932
rect 29148 29486 29150 29538
rect 29202 29486 29204 29538
rect 29148 29474 29204 29486
rect 29372 29538 29428 29550
rect 29372 29486 29374 29538
rect 29426 29486 29428 29538
rect 28812 29316 28868 29326
rect 28812 29222 28868 29260
rect 29372 29316 29428 29486
rect 29372 29250 29428 29260
rect 29484 29314 29540 30830
rect 30268 30884 30324 30942
rect 32508 31666 33348 31668
rect 32508 31614 32958 31666
rect 33010 31614 33294 31666
rect 33346 31614 33348 31666
rect 32508 31612 33348 31614
rect 30716 30884 30772 30894
rect 30268 30882 30772 30884
rect 30268 30830 30718 30882
rect 30770 30830 30772 30882
rect 30268 30828 30772 30830
rect 29932 29988 29988 29998
rect 29932 29650 29988 29932
rect 29932 29598 29934 29650
rect 29986 29598 29988 29650
rect 29932 29586 29988 29598
rect 29484 29262 29486 29314
rect 29538 29262 29540 29314
rect 29484 29250 29540 29262
rect 28588 28802 28644 28812
rect 29372 28868 29428 28878
rect 28364 26898 28420 26908
rect 29372 26962 29428 28812
rect 30268 28644 30324 30828
rect 30716 30818 30772 30828
rect 31388 30098 31444 30110
rect 31388 30046 31390 30098
rect 31442 30046 31444 30098
rect 31052 28756 31108 28766
rect 31052 28662 31108 28700
rect 30156 28588 30268 28644
rect 29372 26910 29374 26962
rect 29426 26910 29428 26962
rect 29372 26898 29428 26910
rect 29484 26964 29540 26974
rect 28252 25454 28254 25506
rect 28306 25454 28308 25506
rect 28252 25442 28308 25454
rect 28924 25564 29428 25620
rect 27804 25396 27860 25406
rect 27804 25302 27860 25340
rect 27468 25284 27524 25294
rect 27468 25190 27524 25228
rect 27692 25282 27748 25294
rect 27692 25230 27694 25282
rect 27746 25230 27748 25282
rect 27692 24612 27748 25230
rect 28924 24946 28980 25564
rect 29372 25506 29428 25564
rect 29372 25454 29374 25506
rect 29426 25454 29428 25506
rect 29372 25442 29428 25454
rect 29260 25396 29316 25406
rect 29260 25302 29316 25340
rect 29148 25284 29204 25294
rect 28924 24894 28926 24946
rect 28978 24894 28980 24946
rect 27692 24546 27748 24556
rect 28476 24612 28532 24622
rect 28476 23716 28532 24556
rect 28476 23650 28532 23660
rect 26684 23326 26686 23378
rect 26738 23326 26740 23378
rect 26684 23314 26740 23326
rect 28924 23380 28980 24894
rect 28924 23314 28980 23324
rect 29036 25282 29204 25284
rect 29036 25230 29150 25282
rect 29202 25230 29204 25282
rect 29036 25228 29204 25230
rect 29036 23268 29092 25228
rect 29148 25218 29204 25228
rect 29484 24164 29540 26908
rect 29708 26964 29764 26974
rect 29820 26964 29876 26974
rect 29708 26962 29820 26964
rect 29708 26910 29710 26962
rect 29762 26910 29820 26962
rect 29708 26908 29820 26910
rect 29708 26898 29764 26908
rect 29596 26180 29652 26190
rect 29596 26178 29764 26180
rect 29596 26126 29598 26178
rect 29650 26126 29764 26178
rect 29596 26124 29764 26126
rect 29596 26114 29652 26124
rect 29708 25506 29764 26124
rect 29708 25454 29710 25506
rect 29762 25454 29764 25506
rect 29708 25284 29764 25454
rect 29708 25218 29764 25228
rect 29820 25508 29876 26908
rect 30044 26180 30100 26190
rect 30156 26180 30212 28588
rect 30268 28550 30324 28588
rect 31388 28644 31444 30046
rect 31388 28578 31444 28588
rect 32508 28532 32564 31612
rect 32956 31602 33012 31612
rect 33292 31602 33348 31612
rect 33516 31556 33572 31566
rect 33516 31462 33572 31500
rect 32620 30996 32676 31006
rect 33180 30996 33236 31006
rect 32620 30994 33236 30996
rect 32620 30942 32622 30994
rect 32674 30942 33182 30994
rect 33234 30942 33236 30994
rect 32620 30940 33236 30942
rect 32620 29988 32676 30940
rect 33180 30930 33236 30940
rect 32620 29922 32676 29932
rect 33068 30436 33124 30446
rect 32508 28466 32564 28476
rect 33068 29538 33124 30380
rect 33180 30324 33236 30334
rect 33180 29652 33236 30268
rect 33180 29650 33348 29652
rect 33180 29598 33182 29650
rect 33234 29598 33348 29650
rect 33180 29596 33348 29598
rect 33180 29586 33236 29596
rect 33068 29486 33070 29538
rect 33122 29486 33124 29538
rect 30268 26964 30324 26974
rect 30268 26870 30324 26908
rect 30100 26124 30212 26180
rect 30044 25508 30100 26124
rect 30044 25452 30324 25508
rect 29708 24164 29764 24174
rect 29484 24162 29764 24164
rect 29484 24110 29710 24162
rect 29762 24110 29764 24162
rect 29484 24108 29764 24110
rect 29260 23940 29316 23950
rect 29484 23940 29540 24108
rect 29708 24098 29764 24108
rect 29260 23938 29540 23940
rect 29260 23886 29262 23938
rect 29314 23886 29540 23938
rect 29260 23884 29540 23886
rect 29260 23874 29316 23884
rect 29484 23716 29540 23726
rect 29484 23622 29540 23660
rect 29148 23268 29204 23278
rect 29036 23212 29148 23268
rect 29148 23174 29204 23212
rect 28924 23154 28980 23166
rect 28924 23102 28926 23154
rect 28978 23102 28980 23154
rect 28924 23044 28980 23102
rect 29484 23154 29540 23166
rect 29484 23102 29486 23154
rect 29538 23102 29540 23154
rect 29484 23044 29540 23102
rect 28924 22988 29540 23044
rect 26572 21812 26628 21822
rect 26572 21700 26628 21756
rect 26684 21700 26740 21710
rect 26572 21698 26740 21700
rect 26572 21646 26686 21698
rect 26738 21646 26740 21698
rect 26572 21644 26740 21646
rect 26684 21634 26740 21644
rect 28924 21700 28980 22988
rect 28924 21606 28980 21644
rect 29596 21700 29652 21710
rect 29596 21606 29652 21644
rect 29820 21026 29876 25452
rect 30156 25284 30212 25294
rect 30156 25190 30212 25228
rect 29932 24162 29988 24174
rect 29932 24110 29934 24162
rect 29986 24110 29988 24162
rect 29932 24050 29988 24110
rect 29932 23998 29934 24050
rect 29986 23998 29988 24050
rect 29932 23380 29988 23998
rect 30268 23940 30324 25452
rect 32508 24724 32564 24734
rect 32732 24724 32788 24734
rect 32508 24722 32732 24724
rect 32508 24670 32510 24722
rect 32562 24670 32732 24722
rect 32508 24668 32732 24670
rect 32508 24658 32564 24668
rect 32732 24658 32788 24668
rect 31724 24612 31780 24622
rect 31724 24050 31780 24556
rect 31724 23998 31726 24050
rect 31778 23998 31780 24050
rect 31724 23986 31780 23998
rect 30268 23874 30324 23884
rect 31052 23940 31108 23950
rect 31052 23846 31108 23884
rect 29932 23042 29988 23324
rect 33068 23268 33124 29486
rect 33180 29204 33236 29214
rect 33180 29110 33236 29148
rect 33180 28756 33236 28766
rect 33292 28756 33348 29596
rect 33180 28754 33348 28756
rect 33180 28702 33182 28754
rect 33234 28702 33348 28754
rect 33180 28700 33348 28702
rect 33180 28690 33236 28700
rect 33516 28532 33572 28542
rect 33404 28530 33572 28532
rect 33404 28478 33518 28530
rect 33570 28478 33572 28530
rect 33404 28476 33572 28478
rect 33180 27748 33236 27758
rect 33404 27748 33460 28476
rect 33516 28466 33572 28476
rect 33628 28308 33684 31892
rect 33852 31780 33908 31790
rect 33852 31778 34020 31780
rect 33852 31726 33854 31778
rect 33906 31726 34020 31778
rect 33852 31724 34020 31726
rect 33852 31714 33908 31724
rect 33964 31666 34020 31724
rect 33964 31614 33966 31666
rect 34018 31614 34020 31666
rect 33964 31602 34020 31614
rect 33740 29204 33796 29214
rect 33740 28642 33796 29148
rect 33852 28756 33908 28766
rect 33908 28700 34020 28756
rect 33852 28690 33908 28700
rect 33740 28590 33742 28642
rect 33794 28590 33796 28642
rect 33740 28578 33796 28590
rect 33964 28642 34020 28700
rect 33964 28590 33966 28642
rect 34018 28590 34020 28642
rect 33964 28578 34020 28590
rect 33180 27746 33460 27748
rect 33180 27694 33182 27746
rect 33234 27694 33460 27746
rect 33180 27692 33460 27694
rect 33516 28252 33684 28308
rect 33180 24724 33236 27692
rect 33516 26852 33572 28252
rect 34076 27972 34132 31892
rect 34300 31778 34356 32620
rect 34300 31726 34302 31778
rect 34354 31726 34356 31778
rect 34300 31714 34356 31726
rect 34412 31780 34468 33182
rect 34412 31714 34468 31724
rect 34524 33740 34804 33796
rect 35196 33740 35460 33750
rect 34188 31554 34244 31566
rect 34188 31502 34190 31554
rect 34242 31502 34244 31554
rect 34188 30324 34244 31502
rect 34188 30258 34244 30268
rect 34524 29764 34580 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35532 32564 35588 36988
rect 36988 36978 37044 36988
rect 37436 36596 37492 36606
rect 37548 36596 37604 37886
rect 38668 37492 38724 39454
rect 39676 39396 39732 39406
rect 39564 39340 39676 39396
rect 39564 38276 39620 39340
rect 39676 39330 39732 39340
rect 39788 38668 39844 40908
rect 40460 40404 40516 40414
rect 41020 40404 41076 40414
rect 40516 40348 40740 40404
rect 40460 40310 40516 40348
rect 40348 40292 40404 40302
rect 39340 38220 39620 38276
rect 38444 37436 38724 37492
rect 39004 37492 39060 37502
rect 39340 37492 39396 38220
rect 39452 38052 39508 38062
rect 39452 37958 39508 37996
rect 39564 38050 39620 38220
rect 39564 37998 39566 38050
rect 39618 37998 39620 38050
rect 39564 37986 39620 37998
rect 39676 38612 39844 38668
rect 40236 40236 40348 40292
rect 39004 37490 39396 37492
rect 39004 37438 39006 37490
rect 39058 37438 39396 37490
rect 39004 37436 39396 37438
rect 38444 37154 38500 37436
rect 39004 37426 39060 37436
rect 38444 37102 38446 37154
rect 38498 37102 38500 37154
rect 38444 37090 38500 37102
rect 38556 37266 38612 37278
rect 38556 37214 38558 37266
rect 38610 37214 38612 37266
rect 38556 36932 38612 37214
rect 38556 36866 38612 36876
rect 38780 37266 38836 37278
rect 38780 37214 38782 37266
rect 38834 37214 38836 37266
rect 37436 36594 37604 36596
rect 37436 36542 37438 36594
rect 37490 36542 37604 36594
rect 37436 36540 37604 36542
rect 37436 36530 37492 36540
rect 36652 36372 36708 36382
rect 36652 35922 36708 36316
rect 36652 35870 36654 35922
rect 36706 35870 36708 35922
rect 36652 35858 36708 35870
rect 37100 36260 37156 36270
rect 36540 35700 36596 35710
rect 36540 35606 36596 35644
rect 36764 35698 36820 35710
rect 36764 35646 36766 35698
rect 36818 35646 36820 35698
rect 36204 35586 36260 35598
rect 36204 35534 36206 35586
rect 36258 35534 36260 35586
rect 36204 35476 36260 35534
rect 36764 35476 36820 35646
rect 37100 35700 37156 36204
rect 37324 36258 37380 36270
rect 37324 36206 37326 36258
rect 37378 36206 37380 36258
rect 37212 35700 37268 35710
rect 37100 35698 37268 35700
rect 37100 35646 37214 35698
rect 37266 35646 37268 35698
rect 37100 35644 37268 35646
rect 36204 35420 36820 35476
rect 35532 32498 35588 32508
rect 35644 34916 35700 34926
rect 36204 34916 36260 35420
rect 35644 34914 36260 34916
rect 35644 34862 35646 34914
rect 35698 34862 36260 34914
rect 35644 34860 36260 34862
rect 34748 32452 34804 32462
rect 34636 31666 34692 31678
rect 34636 31614 34638 31666
rect 34690 31614 34692 31666
rect 34636 30436 34692 31614
rect 34748 31666 34804 32396
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35644 31948 35700 34860
rect 37212 34244 37268 35644
rect 37324 35588 37380 36206
rect 37548 36258 37604 36270
rect 37548 36206 37550 36258
rect 37602 36206 37604 36258
rect 37324 35522 37380 35532
rect 37436 36036 37492 36046
rect 37436 35138 37492 35980
rect 37436 35086 37438 35138
rect 37490 35086 37492 35138
rect 37436 35074 37492 35086
rect 37548 35700 37604 36206
rect 38780 36036 38836 37214
rect 39228 37268 39284 37278
rect 39116 36260 39172 36270
rect 39116 36166 39172 36204
rect 38780 35970 38836 35980
rect 37548 34916 37604 35644
rect 37324 34860 37604 34916
rect 37324 34802 37380 34860
rect 37324 34750 37326 34802
rect 37378 34750 37380 34802
rect 37324 34468 37380 34750
rect 37436 34692 37492 34702
rect 37436 34690 37716 34692
rect 37436 34638 37438 34690
rect 37490 34638 37716 34690
rect 37436 34636 37716 34638
rect 37436 34626 37492 34636
rect 37324 34412 37604 34468
rect 37436 34244 37492 34254
rect 37212 34242 37492 34244
rect 37212 34190 37438 34242
rect 37490 34190 37492 34242
rect 37212 34188 37492 34190
rect 37100 34130 37156 34142
rect 37100 34078 37102 34130
rect 37154 34078 37156 34130
rect 36764 34020 36820 34030
rect 37100 34020 37156 34078
rect 36764 34018 37156 34020
rect 36764 33966 36766 34018
rect 36818 33966 37156 34018
rect 36764 33964 37156 33966
rect 36428 32564 36484 32574
rect 36428 32470 36484 32508
rect 35980 32452 36036 32462
rect 35980 32358 36036 32396
rect 35644 31892 35924 31948
rect 34748 31614 34750 31666
rect 34802 31614 34804 31666
rect 34748 31602 34804 31614
rect 34972 31556 35028 31566
rect 34972 31462 35028 31500
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34636 30370 34692 30380
rect 34524 29698 34580 29708
rect 35756 29764 35812 29774
rect 34188 29204 34244 29214
rect 34188 28642 34244 29148
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35084 28868 35140 28878
rect 35084 28756 35140 28812
rect 35084 28754 35476 28756
rect 35084 28702 35086 28754
rect 35138 28702 35476 28754
rect 35084 28700 35476 28702
rect 35084 28690 35140 28700
rect 34188 28590 34190 28642
rect 34242 28590 34244 28642
rect 34188 28578 34244 28590
rect 35420 28642 35476 28700
rect 35420 28590 35422 28642
rect 35474 28590 35476 28642
rect 35420 28578 35476 28590
rect 35756 28532 35812 29708
rect 35532 28530 35812 28532
rect 35532 28478 35758 28530
rect 35810 28478 35812 28530
rect 35532 28476 35812 28478
rect 34076 27916 35028 27972
rect 33628 27748 33684 27758
rect 33628 27746 34356 27748
rect 33628 27694 33630 27746
rect 33682 27694 34356 27746
rect 33628 27692 34356 27694
rect 33628 27682 33684 27692
rect 33516 26796 34020 26852
rect 33964 26290 34020 26796
rect 33964 26238 33966 26290
rect 34018 26238 34020 26290
rect 33964 25620 34020 26238
rect 33964 25554 34020 25564
rect 33852 25508 33908 25518
rect 33740 25452 33852 25508
rect 33236 24668 33348 24724
rect 33180 24630 33236 24668
rect 33292 23492 33348 24668
rect 33068 23174 33124 23212
rect 33180 23266 33236 23278
rect 33180 23214 33182 23266
rect 33234 23214 33236 23266
rect 33180 23156 33236 23214
rect 33292 23156 33348 23436
rect 33404 24722 33460 24734
rect 33404 24670 33406 24722
rect 33458 24670 33460 24722
rect 33404 23378 33460 24670
rect 33740 24722 33796 25452
rect 33852 25442 33908 25452
rect 33740 24670 33742 24722
rect 33794 24670 33796 24722
rect 33740 24658 33796 24670
rect 33516 24612 33572 24622
rect 33516 24518 33572 24556
rect 33404 23326 33406 23378
rect 33458 23326 33460 23378
rect 33404 23314 33460 23326
rect 33852 24050 33908 24062
rect 33852 23998 33854 24050
rect 33906 23998 33908 24050
rect 33852 23156 33908 23998
rect 34300 24052 34356 27692
rect 34748 26178 34804 26190
rect 34748 26126 34750 26178
rect 34802 26126 34804 26178
rect 34748 25732 34804 26126
rect 34748 25666 34804 25676
rect 34972 25618 35028 27916
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35420 27076 35476 27086
rect 35532 27076 35588 28476
rect 35756 28466 35812 28476
rect 35420 27074 35588 27076
rect 35420 27022 35422 27074
rect 35474 27022 35588 27074
rect 35420 27020 35588 27022
rect 35420 27010 35476 27020
rect 34972 25566 34974 25618
rect 35026 25566 35028 25618
rect 34972 25284 35028 25566
rect 35084 26850 35140 26862
rect 35084 26798 35086 26850
rect 35138 26798 35140 26850
rect 35084 25508 35140 26798
rect 35308 26852 35364 26862
rect 35308 26758 35364 26796
rect 35868 26404 35924 31892
rect 36540 31556 36596 31566
rect 36316 29428 36372 29438
rect 36540 29428 36596 31500
rect 36652 29540 36708 29550
rect 36652 29446 36708 29484
rect 36316 29426 36596 29428
rect 36316 29374 36318 29426
rect 36370 29374 36596 29426
rect 36316 29372 36596 29374
rect 35980 29316 36036 29326
rect 36316 29316 36372 29372
rect 35980 29314 36372 29316
rect 35980 29262 35982 29314
rect 36034 29262 36372 29314
rect 35980 29260 36372 29262
rect 35980 28868 36036 29260
rect 35980 28802 36036 28812
rect 36428 27188 36484 27198
rect 36428 27094 36484 27132
rect 36764 27188 36820 33964
rect 37436 33572 37492 34188
rect 37436 33506 37492 33516
rect 36876 32564 36932 32574
rect 36876 30882 36932 32508
rect 37548 31948 37604 34412
rect 37660 32452 37716 34636
rect 37660 32386 37716 32396
rect 39116 33572 39172 33582
rect 37324 31892 37604 31948
rect 37324 31666 37380 31892
rect 37324 31614 37326 31666
rect 37378 31614 37380 31666
rect 37324 31602 37380 31614
rect 38780 31666 38836 31678
rect 38780 31614 38782 31666
rect 38834 31614 38836 31666
rect 36988 31556 37044 31566
rect 36988 31462 37044 31500
rect 36876 30830 36878 30882
rect 36930 30830 36932 30882
rect 36876 30212 36932 30830
rect 37436 30322 37492 30334
rect 37436 30270 37438 30322
rect 37490 30270 37492 30322
rect 37100 30212 37156 30222
rect 36876 30156 37100 30212
rect 37100 30118 37156 30156
rect 37436 29652 37492 30270
rect 37660 29764 37716 29774
rect 37548 29652 37604 29662
rect 37436 29596 37548 29652
rect 37548 29558 37604 29596
rect 37212 29540 37268 29550
rect 36764 27122 36820 27132
rect 37100 27188 37156 27198
rect 37100 27074 37156 27132
rect 37100 27022 37102 27074
rect 37154 27022 37156 27074
rect 37100 27010 37156 27022
rect 36876 26852 36932 26862
rect 35868 26348 36036 26404
rect 35868 26180 35924 26190
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35420 25732 35476 25742
rect 35420 25618 35476 25676
rect 35420 25566 35422 25618
rect 35474 25566 35476 25618
rect 35420 25554 35476 25566
rect 35084 25442 35140 25452
rect 35196 25506 35252 25518
rect 35196 25454 35198 25506
rect 35250 25454 35252 25506
rect 35196 25396 35252 25454
rect 35868 25506 35924 26124
rect 35868 25454 35870 25506
rect 35922 25454 35924 25506
rect 35868 25442 35924 25454
rect 35196 25284 35252 25340
rect 34972 25228 35252 25284
rect 35644 25394 35700 25406
rect 35644 25342 35646 25394
rect 35698 25342 35700 25394
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35644 24164 35700 25342
rect 35756 24164 35812 24174
rect 35644 24162 35812 24164
rect 35644 24110 35758 24162
rect 35810 24110 35812 24162
rect 35644 24108 35812 24110
rect 34300 23958 34356 23996
rect 35532 24052 35588 24062
rect 35532 23958 35588 23996
rect 33292 23100 33684 23156
rect 33180 23090 33236 23100
rect 29932 22990 29934 23042
rect 29986 22990 29988 23042
rect 29932 22978 29988 22990
rect 30044 21756 30436 21812
rect 30044 21698 30100 21756
rect 30044 21646 30046 21698
rect 30098 21646 30100 21698
rect 30044 21634 30100 21646
rect 29820 20974 29822 21026
rect 29874 20974 29876 21026
rect 29820 20962 29876 20974
rect 30156 21588 30212 21598
rect 30156 20802 30212 21532
rect 30156 20750 30158 20802
rect 30210 20750 30212 20802
rect 30156 20738 30212 20750
rect 30380 20802 30436 21756
rect 30380 20750 30382 20802
rect 30434 20750 30436 20802
rect 28028 20020 28084 20030
rect 27580 19346 27636 19358
rect 27580 19294 27582 19346
rect 27634 19294 27636 19346
rect 27580 18564 27636 19294
rect 28028 19348 28084 19964
rect 29484 20020 29540 20030
rect 29484 19926 29540 19964
rect 30380 20020 30436 20750
rect 30604 21700 30660 21710
rect 30604 20802 30660 21644
rect 30604 20750 30606 20802
rect 30658 20750 30660 20802
rect 30492 20244 30548 20254
rect 30492 20020 30548 20188
rect 30604 20188 30660 20750
rect 31276 20244 31332 20254
rect 30604 20132 30772 20188
rect 30380 19964 30548 20020
rect 30156 19906 30212 19918
rect 30156 19854 30158 19906
rect 30210 19854 30212 19906
rect 30156 19458 30212 19854
rect 30156 19406 30158 19458
rect 30210 19406 30212 19458
rect 30156 19394 30212 19406
rect 30380 19460 30436 19964
rect 30492 19460 30548 19470
rect 30380 19458 30548 19460
rect 30380 19406 30494 19458
rect 30546 19406 30548 19458
rect 30380 19404 30548 19406
rect 30492 19394 30548 19404
rect 28028 19254 28084 19292
rect 30268 19234 30324 19246
rect 30268 19182 30270 19234
rect 30322 19182 30324 19234
rect 27580 15428 27636 18508
rect 29820 19012 29876 19022
rect 29596 16884 29652 16894
rect 28700 15876 28756 15886
rect 27804 15428 27860 15438
rect 27580 15426 27860 15428
rect 27580 15374 27806 15426
rect 27858 15374 27860 15426
rect 27580 15372 27860 15374
rect 27804 15362 27860 15372
rect 28700 14644 28756 15820
rect 29036 15314 29092 15326
rect 29036 15262 29038 15314
rect 29090 15262 29092 15314
rect 29036 14756 29092 15262
rect 29596 15202 29652 16828
rect 29596 15150 29598 15202
rect 29650 15150 29652 15202
rect 29596 15138 29652 15150
rect 29036 14700 29316 14756
rect 29260 14644 29316 14700
rect 28700 14642 29204 14644
rect 28700 14590 28702 14642
rect 28754 14590 29204 14642
rect 28700 14588 29204 14590
rect 28700 14578 28756 14588
rect 29148 14530 29204 14588
rect 29148 14478 29150 14530
rect 29202 14478 29204 14530
rect 29148 14466 29204 14478
rect 27244 13860 27300 13870
rect 27244 13766 27300 13804
rect 26572 13748 26628 13758
rect 26572 13654 26628 13692
rect 29260 13636 29316 14588
rect 29372 13636 29428 13646
rect 29260 13634 29428 13636
rect 29260 13582 29374 13634
rect 29426 13582 29428 13634
rect 29260 13580 29428 13582
rect 29372 13570 29428 13580
rect 28140 11394 28196 11406
rect 28140 11342 28142 11394
rect 28194 11342 28196 11394
rect 27356 11284 27412 11294
rect 27356 11190 27412 11228
rect 28140 10836 28196 11342
rect 28588 11170 28644 11182
rect 28588 11118 28590 11170
rect 28642 11118 28644 11170
rect 28588 10836 28644 11118
rect 28140 10780 28588 10836
rect 26460 9538 26516 9548
rect 25116 8306 25172 8316
rect 25676 8372 26180 8428
rect 25676 8036 25732 8372
rect 25340 7700 25396 7710
rect 25340 7606 25396 7644
rect 24668 7310 24670 7362
rect 24722 7310 24724 7362
rect 24668 7298 24724 7310
rect 24556 5122 24612 6748
rect 25452 6132 25508 6142
rect 25676 6132 25732 7980
rect 27804 7700 27860 7710
rect 27468 6692 27524 6702
rect 26236 6132 26292 6142
rect 25452 6130 26292 6132
rect 25452 6078 25454 6130
rect 25506 6078 26238 6130
rect 26290 6078 26292 6130
rect 25452 6076 26292 6078
rect 25452 6066 25508 6076
rect 26236 6066 26292 6076
rect 27468 5906 27524 6636
rect 27468 5854 27470 5906
rect 27522 5854 27524 5906
rect 25676 5796 25732 5806
rect 25676 5702 25732 5740
rect 26796 5796 26852 5806
rect 26796 5702 26852 5740
rect 25340 5684 25396 5694
rect 25228 5682 25396 5684
rect 25228 5630 25342 5682
rect 25394 5630 25396 5682
rect 25228 5628 25396 5630
rect 25228 5234 25284 5628
rect 25340 5618 25396 5628
rect 25228 5182 25230 5234
rect 25282 5182 25284 5234
rect 25228 5170 25284 5182
rect 27356 5236 27412 5246
rect 27468 5236 27524 5854
rect 27692 5796 27748 5806
rect 27692 5702 27748 5740
rect 27356 5234 27524 5236
rect 27356 5182 27358 5234
rect 27410 5182 27524 5234
rect 27356 5180 27524 5182
rect 27804 5234 27860 7644
rect 28364 7700 28420 10780
rect 28476 10610 28532 10780
rect 28588 10770 28644 10780
rect 28476 10558 28478 10610
rect 28530 10558 28532 10610
rect 28476 10546 28532 10558
rect 29148 10498 29204 10510
rect 29148 10446 29150 10498
rect 29202 10446 29204 10498
rect 29148 10052 29204 10446
rect 29596 10052 29652 10062
rect 29148 10050 29652 10052
rect 29148 9998 29598 10050
rect 29650 9998 29652 10050
rect 29148 9996 29652 9998
rect 29596 9986 29652 9996
rect 29708 10052 29764 10062
rect 29820 10052 29876 18956
rect 30268 19012 30324 19182
rect 30268 18946 30324 18956
rect 30604 19234 30660 19246
rect 30604 19182 30606 19234
rect 30658 19182 30660 19234
rect 30604 18788 30660 19182
rect 30604 18722 30660 18732
rect 30492 18228 30548 18238
rect 30492 17108 30548 18172
rect 30492 17014 30548 17052
rect 30044 14644 30100 14654
rect 30044 13970 30100 14588
rect 30044 13918 30046 13970
rect 30098 13918 30100 13970
rect 30044 13748 30100 13918
rect 30044 10836 30100 13692
rect 30044 10770 30100 10780
rect 29708 10050 29876 10052
rect 29708 9998 29710 10050
rect 29762 9998 29876 10050
rect 29708 9996 29876 9998
rect 30156 10052 30212 10062
rect 29372 9828 29428 9838
rect 29708 9828 29764 9996
rect 29372 9826 29764 9828
rect 29372 9774 29374 9826
rect 29426 9774 29764 9826
rect 29372 9772 29764 9774
rect 29932 9828 29988 9838
rect 29372 9762 29428 9772
rect 29932 9734 29988 9772
rect 30156 9826 30212 9996
rect 30156 9774 30158 9826
rect 30210 9774 30212 9826
rect 30156 8428 30212 9774
rect 30604 9828 30660 9838
rect 30604 9734 30660 9772
rect 30492 9714 30548 9726
rect 30492 9662 30494 9714
rect 30546 9662 30548 9714
rect 30492 9044 30548 9662
rect 30492 8978 30548 8988
rect 30604 9604 30660 9614
rect 28364 7634 28420 7644
rect 30044 8372 30212 8428
rect 29820 6692 29876 6702
rect 29820 6598 29876 6636
rect 30044 6132 30100 8372
rect 30380 6578 30436 6590
rect 30380 6526 30382 6578
rect 30434 6526 30436 6578
rect 29148 6130 30100 6132
rect 29148 6078 30046 6130
rect 30098 6078 30100 6130
rect 29148 6076 30100 6078
rect 28700 6020 28756 6030
rect 28700 5926 28756 5964
rect 28812 6020 28868 6030
rect 29148 6020 29204 6076
rect 30044 6066 30100 6076
rect 30268 6132 30324 6142
rect 30380 6132 30436 6526
rect 30268 6130 30436 6132
rect 30268 6078 30270 6130
rect 30322 6078 30436 6130
rect 30268 6076 30436 6078
rect 30604 6132 30660 9548
rect 30716 8428 30772 20132
rect 31276 19458 31332 20188
rect 33628 20188 33684 23100
rect 33852 23090 33908 23100
rect 34972 23156 35028 23166
rect 34972 23062 35028 23100
rect 35420 23156 35476 23166
rect 35644 23156 35700 24108
rect 35756 24098 35812 24108
rect 35868 24052 35924 24062
rect 35980 24052 36036 26348
rect 36876 26292 36932 26796
rect 37212 26516 37268 29484
rect 37660 29538 37716 29708
rect 38780 29650 38836 31614
rect 39004 31666 39060 31678
rect 39004 31614 39006 31666
rect 39058 31614 39060 31666
rect 39004 29988 39060 31614
rect 39004 29922 39060 29932
rect 38780 29598 38782 29650
rect 38834 29598 38836 29650
rect 38780 29586 38836 29598
rect 38892 29652 38948 29662
rect 38892 29558 38948 29596
rect 39116 29650 39172 33516
rect 39228 32676 39284 37212
rect 39564 37268 39620 37278
rect 39564 37174 39620 37212
rect 39452 36596 39508 36606
rect 39452 36502 39508 36540
rect 39340 36484 39396 36494
rect 39340 36390 39396 36428
rect 39564 36258 39620 36270
rect 39564 36206 39566 36258
rect 39618 36206 39620 36258
rect 39564 35700 39620 36206
rect 39564 35634 39620 35644
rect 39228 32610 39284 32620
rect 39340 31780 39396 31790
rect 39340 31686 39396 31724
rect 39228 31554 39284 31566
rect 39228 31502 39230 31554
rect 39282 31502 39284 31554
rect 39228 30884 39284 31502
rect 39228 30828 39620 30884
rect 39564 30322 39620 30828
rect 39564 30270 39566 30322
rect 39618 30270 39620 30322
rect 39564 30258 39620 30270
rect 39116 29598 39118 29650
rect 39170 29598 39172 29650
rect 39116 29586 39172 29598
rect 37660 29486 37662 29538
rect 37714 29486 37716 29538
rect 37660 29474 37716 29486
rect 38668 29540 38724 29550
rect 38668 29446 38724 29484
rect 37548 29204 37604 29214
rect 37548 29110 37604 29148
rect 37660 26964 37716 26974
rect 37436 26852 37492 26862
rect 37660 26852 37716 26908
rect 37436 26850 37716 26852
rect 37436 26798 37438 26850
rect 37490 26798 37716 26850
rect 37436 26796 37716 26798
rect 37436 26786 37492 26796
rect 37212 26422 37268 26460
rect 37660 26514 37716 26796
rect 38780 26964 38836 26974
rect 37660 26462 37662 26514
rect 37714 26462 37716 26514
rect 37660 26450 37716 26462
rect 38220 26516 38276 26526
rect 36876 26178 36932 26236
rect 37436 26292 37492 26302
rect 37436 26198 37492 26236
rect 36876 26126 36878 26178
rect 36930 26126 36932 26178
rect 36876 26114 36932 26126
rect 37324 26180 37380 26190
rect 37324 26086 37380 26124
rect 37212 25620 37268 25630
rect 37212 25526 37268 25564
rect 35924 23996 36036 24052
rect 36764 25396 36820 25406
rect 35868 23958 35924 23996
rect 36764 23492 36820 25340
rect 38220 25396 38276 26460
rect 38220 24946 38276 25340
rect 38220 24894 38222 24946
rect 38274 24894 38276 24946
rect 38220 24882 38276 24894
rect 38444 24722 38500 24734
rect 38444 24670 38446 24722
rect 38498 24670 38500 24722
rect 38332 24610 38388 24622
rect 38332 24558 38334 24610
rect 38386 24558 38388 24610
rect 38332 23940 38388 24558
rect 35868 23268 35924 23278
rect 36764 23268 36820 23436
rect 37324 23884 38388 23940
rect 35868 23266 36708 23268
rect 35868 23214 35870 23266
rect 35922 23214 36708 23266
rect 35868 23212 36708 23214
rect 35868 23202 35924 23212
rect 35420 23154 35700 23156
rect 35420 23102 35422 23154
rect 35474 23102 35700 23154
rect 35420 23100 35700 23102
rect 36652 23154 36708 23212
rect 36652 23102 36654 23154
rect 36706 23102 36708 23154
rect 35420 23090 35476 23100
rect 36652 23090 36708 23102
rect 36764 23212 37044 23268
rect 36540 23042 36596 23054
rect 36540 22990 36542 23042
rect 36594 22990 36596 23042
rect 36540 22932 36596 22990
rect 36764 22932 36820 23212
rect 36988 23154 37044 23212
rect 37324 23266 37380 23884
rect 37324 23214 37326 23266
rect 37378 23214 37380 23266
rect 37324 23202 37380 23214
rect 36988 23102 36990 23154
rect 37042 23102 37044 23154
rect 36988 23090 37044 23102
rect 38444 23156 38500 24670
rect 38780 24722 38836 26908
rect 39452 26964 39508 27002
rect 39452 26898 39508 26908
rect 39676 25284 39732 38612
rect 39900 37940 39956 37950
rect 39900 37846 39956 37884
rect 39788 37828 39844 37838
rect 39788 37734 39844 37772
rect 39788 37492 39844 37502
rect 40236 37492 40292 40236
rect 40348 40226 40404 40236
rect 40684 37828 40740 40348
rect 41020 40310 41076 40348
rect 41804 40292 41860 40302
rect 41804 40198 41860 40236
rect 42700 40292 42756 40302
rect 40796 39732 40852 39742
rect 41244 39732 41300 39742
rect 40796 39730 41300 39732
rect 40796 39678 40798 39730
rect 40850 39678 41246 39730
rect 41298 39678 41300 39730
rect 40796 39676 41300 39678
rect 40796 39666 40852 39676
rect 41244 39666 41300 39676
rect 42700 39730 42756 40236
rect 43932 40292 43988 41134
rect 43932 40198 43988 40236
rect 42700 39678 42702 39730
rect 42754 39678 42756 39730
rect 42700 39666 42756 39678
rect 41132 39396 41188 39406
rect 41132 39302 41188 39340
rect 42588 39394 42644 39406
rect 42588 39342 42590 39394
rect 42642 39342 42644 39394
rect 40796 37828 40852 37838
rect 40684 37826 40852 37828
rect 40684 37774 40798 37826
rect 40850 37774 40852 37826
rect 40684 37772 40852 37774
rect 40236 37436 40404 37492
rect 39788 37398 39844 37436
rect 39900 37380 39956 37390
rect 39900 37378 40180 37380
rect 39900 37326 39902 37378
rect 39954 37326 40180 37378
rect 39900 37324 40180 37326
rect 39900 37314 39956 37324
rect 39900 36932 39956 36942
rect 39900 36260 39956 36876
rect 40012 36260 40068 36270
rect 39900 36204 40012 36260
rect 39900 27300 39956 36204
rect 40012 36166 40068 36204
rect 40124 36036 40180 37324
rect 40236 37266 40292 37278
rect 40236 37214 40238 37266
rect 40290 37214 40292 37266
rect 40236 36932 40292 37214
rect 40348 37154 40404 37436
rect 40796 37268 40852 37772
rect 41916 37828 41972 37838
rect 41916 37378 41972 37772
rect 42588 37492 42644 39342
rect 42588 37426 42644 37436
rect 41916 37326 41918 37378
rect 41970 37326 41972 37378
rect 41916 37314 41972 37326
rect 41244 37268 41300 37278
rect 40796 37266 41300 37268
rect 40796 37214 41246 37266
rect 41298 37214 41300 37266
rect 40796 37212 41300 37214
rect 40348 37102 40350 37154
rect 40402 37102 40404 37154
rect 40348 37090 40404 37102
rect 40236 36866 40292 36876
rect 40124 35970 40180 35980
rect 40348 36484 40404 36494
rect 40236 34802 40292 34814
rect 40236 34750 40238 34802
rect 40290 34750 40292 34802
rect 40236 32676 40292 34750
rect 40348 34802 40404 36428
rect 40572 36260 40628 36270
rect 40572 36166 40628 36204
rect 40908 36036 40964 36046
rect 40908 35138 40964 35980
rect 40908 35086 40910 35138
rect 40962 35086 40964 35138
rect 40908 35074 40964 35086
rect 40348 34750 40350 34802
rect 40402 34750 40404 34802
rect 40348 34738 40404 34750
rect 40796 34802 40852 34814
rect 40796 34750 40798 34802
rect 40850 34750 40852 34802
rect 40572 34690 40628 34702
rect 40572 34638 40574 34690
rect 40626 34638 40628 34690
rect 40236 32610 40292 32620
rect 40348 34018 40404 34030
rect 40348 33966 40350 34018
rect 40402 33966 40404 34018
rect 40348 30212 40404 33966
rect 40572 33346 40628 34638
rect 40572 33294 40574 33346
rect 40626 33294 40628 33346
rect 40572 33282 40628 33294
rect 40460 33122 40516 33134
rect 40460 33070 40462 33122
rect 40514 33070 40516 33122
rect 40460 31892 40516 33070
rect 40460 31826 40516 31836
rect 40348 29652 40404 30156
rect 40796 29764 40852 34750
rect 40908 34690 40964 34702
rect 40908 34638 40910 34690
rect 40962 34638 40964 34690
rect 40908 33796 40964 34638
rect 41244 34130 41300 37212
rect 44044 37154 44100 37166
rect 44044 37102 44046 37154
rect 44098 37102 44100 37154
rect 44044 36484 44100 37102
rect 44044 36418 44100 36428
rect 41244 34078 41246 34130
rect 41298 34078 41300 34130
rect 41244 34066 41300 34078
rect 41916 34020 41972 34030
rect 40908 33730 40964 33740
rect 41356 34018 41972 34020
rect 41356 33966 41918 34018
rect 41970 33966 41972 34018
rect 41356 33964 41972 33966
rect 41244 33572 41300 33582
rect 41356 33572 41412 33964
rect 41916 33954 41972 33964
rect 44044 34018 44100 34030
rect 44044 33966 44046 34018
rect 44098 33966 44100 34018
rect 41244 33570 41412 33572
rect 41244 33518 41246 33570
rect 41298 33518 41412 33570
rect 41244 33516 41412 33518
rect 41580 33796 41636 33806
rect 41244 33506 41300 33516
rect 40908 33348 40964 33358
rect 41356 33348 41412 33358
rect 40908 33346 41412 33348
rect 40908 33294 40910 33346
rect 40962 33294 41358 33346
rect 41410 33294 41412 33346
rect 40908 33292 41412 33294
rect 40908 33282 40964 33292
rect 41356 33282 41412 33292
rect 41580 33234 41636 33740
rect 44044 33796 44100 33966
rect 44044 33730 44100 33740
rect 41580 33182 41582 33234
rect 41634 33182 41636 33234
rect 41580 33170 41636 33182
rect 41692 33236 41748 33246
rect 42140 33236 42196 33246
rect 41692 33234 42196 33236
rect 41692 33182 41694 33234
rect 41746 33182 42142 33234
rect 42194 33182 42196 33234
rect 41692 33180 42196 33182
rect 41132 33122 41188 33134
rect 41132 33070 41134 33122
rect 41186 33070 41188 33122
rect 41132 31892 41188 33070
rect 41132 31826 41188 31836
rect 40796 29698 40852 29708
rect 41468 29988 41524 29998
rect 40348 29558 40404 29596
rect 41132 29652 41188 29662
rect 41132 29426 41188 29596
rect 41132 29374 41134 29426
rect 41186 29374 41188 29426
rect 41132 29362 41188 29374
rect 40460 29316 40516 29326
rect 40012 28756 40068 28766
rect 40012 28662 40068 28700
rect 40460 28754 40516 29260
rect 40460 28702 40462 28754
rect 40514 28702 40516 28754
rect 40460 28644 40516 28702
rect 41244 28866 41300 28878
rect 41244 28814 41246 28866
rect 41298 28814 41300 28866
rect 40460 28578 40516 28588
rect 41132 28644 41188 28654
rect 41132 28084 41188 28588
rect 41244 28196 41300 28814
rect 41468 28642 41524 29932
rect 41692 29428 41748 33180
rect 42140 33170 42196 33180
rect 42700 30100 42756 30110
rect 42700 30006 42756 30044
rect 44044 30100 44100 30110
rect 42588 29988 42644 29998
rect 42588 29894 42644 29932
rect 41468 28590 41470 28642
rect 41522 28590 41524 28642
rect 41468 28578 41524 28590
rect 41580 29372 41748 29428
rect 41580 28756 41636 29372
rect 41916 29314 41972 29326
rect 41916 29262 41918 29314
rect 41970 29262 41972 29314
rect 41580 28532 41636 28700
rect 41692 28756 41748 28766
rect 41916 28756 41972 29262
rect 44044 29314 44100 30044
rect 44044 29262 44046 29314
rect 44098 29262 44100 29314
rect 44044 29250 44100 29262
rect 41692 28754 41972 28756
rect 41692 28702 41694 28754
rect 41746 28702 41972 28754
rect 41692 28700 41972 28702
rect 41692 28690 41748 28700
rect 41804 28532 41860 28542
rect 41580 28530 41860 28532
rect 41580 28478 41806 28530
rect 41858 28478 41860 28530
rect 41580 28476 41860 28478
rect 41244 28140 41412 28196
rect 41132 28028 41300 28084
rect 39900 27186 39956 27244
rect 39900 27134 39902 27186
rect 39954 27134 39956 27186
rect 39900 27122 39956 27134
rect 40348 27860 40404 27870
rect 41132 27860 41188 27870
rect 40348 27858 41188 27860
rect 40348 27806 40350 27858
rect 40402 27806 41134 27858
rect 41186 27806 41188 27858
rect 40348 27804 41188 27806
rect 40236 27076 40292 27086
rect 40124 26964 40180 26974
rect 40124 26404 40180 26908
rect 40012 26348 40180 26404
rect 39900 25620 39956 25630
rect 39900 25526 39956 25564
rect 40012 25506 40068 26348
rect 40012 25454 40014 25506
rect 40066 25454 40068 25506
rect 40012 25442 40068 25454
rect 40124 26180 40180 26190
rect 40236 26180 40292 27020
rect 40124 26178 40292 26180
rect 40124 26126 40126 26178
rect 40178 26126 40292 26178
rect 40124 26124 40292 26126
rect 39676 25218 39732 25228
rect 38780 24670 38782 24722
rect 38834 24670 38836 24722
rect 38780 24658 38836 24670
rect 39116 24052 39172 24062
rect 39116 23380 39172 23996
rect 40124 24052 40180 26124
rect 40348 24836 40404 27804
rect 41132 27794 41188 27804
rect 41020 27186 41076 27198
rect 41020 27134 41022 27186
rect 41074 27134 41076 27186
rect 40796 27076 40852 27114
rect 40796 27010 40852 27020
rect 41020 26908 41076 27134
rect 40572 26852 41076 26908
rect 40460 25508 40516 25518
rect 40572 25508 40628 26852
rect 40516 25452 40628 25508
rect 41132 25620 41188 25630
rect 41132 25506 41188 25564
rect 41132 25454 41134 25506
rect 41186 25454 41188 25506
rect 40460 25414 40516 25452
rect 41132 25442 41188 25454
rect 40684 25396 40740 25406
rect 40684 25302 40740 25340
rect 40572 25282 40628 25294
rect 41244 25284 41300 28028
rect 41356 28082 41412 28140
rect 41356 28030 41358 28082
rect 41410 28030 41412 28082
rect 41356 28018 41412 28030
rect 41468 27634 41524 27646
rect 41468 27582 41470 27634
rect 41522 27582 41524 27634
rect 41468 27186 41524 27582
rect 41468 27134 41470 27186
rect 41522 27134 41524 27186
rect 41468 27122 41524 27134
rect 41804 25620 41860 28476
rect 44044 25620 44100 25630
rect 41804 25564 42084 25620
rect 40572 25230 40574 25282
rect 40626 25230 40628 25282
rect 40572 24948 40628 25230
rect 41132 25228 41300 25284
rect 41916 25394 41972 25406
rect 41916 25342 41918 25394
rect 41970 25342 41972 25394
rect 40572 24892 40964 24948
rect 40348 24780 40516 24836
rect 40124 23986 40180 23996
rect 40348 24610 40404 24622
rect 40348 24558 40350 24610
rect 40402 24558 40404 24610
rect 40348 23604 40404 24558
rect 40348 23538 40404 23548
rect 40012 23380 40068 23390
rect 40460 23380 40516 24780
rect 40908 24834 40964 24892
rect 40908 24782 40910 24834
rect 40962 24782 40964 24834
rect 40908 24770 40964 24782
rect 40684 23716 40740 23726
rect 40684 23622 40740 23660
rect 39116 23378 39732 23380
rect 39116 23326 39118 23378
rect 39170 23326 39732 23378
rect 39116 23324 39732 23326
rect 39116 23314 39172 23324
rect 39452 23156 39508 23166
rect 38444 23090 38500 23100
rect 39228 23100 39452 23156
rect 36540 22876 36820 22932
rect 36876 23042 36932 23054
rect 36876 22990 36878 23042
rect 36930 22990 36932 23042
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 36876 21812 36932 22990
rect 36876 21756 37156 21812
rect 37100 21698 37156 21756
rect 37100 21646 37102 21698
rect 37154 21646 37156 21698
rect 37100 21634 37156 21646
rect 35980 21588 36036 21598
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 33628 20132 34020 20188
rect 31276 19406 31278 19458
rect 31330 19406 31332 19458
rect 31276 19394 31332 19406
rect 32284 19906 32340 19918
rect 32284 19854 32286 19906
rect 32338 19854 32340 19906
rect 31724 19236 31780 19246
rect 31724 19142 31780 19180
rect 31948 19234 32004 19246
rect 31948 19182 31950 19234
rect 32002 19182 32004 19234
rect 31612 18788 31668 18798
rect 31668 18732 31892 18788
rect 31612 18722 31668 18732
rect 31836 18674 31892 18732
rect 31836 18622 31838 18674
rect 31890 18622 31892 18674
rect 31052 17444 31108 17454
rect 30940 17108 30996 17118
rect 30940 17014 30996 17052
rect 31052 16994 31108 17388
rect 31052 16942 31054 16994
rect 31106 16942 31108 16994
rect 31052 16930 31108 16942
rect 31612 16884 31668 16922
rect 31612 16818 31668 16828
rect 31836 16772 31892 18622
rect 31948 18452 32004 19182
rect 32284 19236 32340 19854
rect 33180 19908 33236 19918
rect 32396 19236 32452 19246
rect 32284 19180 32396 19236
rect 32172 18452 32228 18462
rect 31948 18396 32172 18452
rect 32172 18358 32228 18396
rect 32396 18338 32452 19180
rect 32396 18286 32398 18338
rect 32450 18286 32452 18338
rect 32396 17554 32452 18286
rect 32396 17502 32398 17554
rect 32450 17502 32452 17554
rect 32396 17490 32452 17502
rect 32844 18452 32900 18462
rect 32844 17554 32900 18396
rect 32844 17502 32846 17554
rect 32898 17502 32900 17554
rect 32844 17490 32900 17502
rect 32956 17668 33012 17678
rect 32284 17444 32340 17454
rect 32284 17350 32340 17388
rect 32956 17108 33012 17612
rect 32956 17042 33012 17052
rect 32508 16884 32564 16894
rect 33068 16884 33124 16894
rect 32508 16882 33124 16884
rect 32508 16830 32510 16882
rect 32562 16830 33070 16882
rect 33122 16830 33124 16882
rect 32508 16828 33124 16830
rect 31948 16772 32004 16782
rect 31836 16770 32004 16772
rect 31836 16718 31950 16770
rect 32002 16718 32004 16770
rect 31836 16716 32004 16718
rect 31948 16706 32004 16716
rect 30940 16658 30996 16670
rect 31612 16660 31668 16670
rect 30940 16606 30942 16658
rect 30994 16606 30996 16658
rect 30940 16324 30996 16606
rect 31388 16658 31668 16660
rect 31388 16606 31614 16658
rect 31666 16606 31668 16658
rect 31388 16604 31668 16606
rect 31052 16324 31108 16334
rect 30940 16322 31108 16324
rect 30940 16270 31054 16322
rect 31106 16270 31108 16322
rect 30940 16268 31108 16270
rect 31052 16258 31108 16268
rect 31276 16210 31332 16222
rect 31276 16158 31278 16210
rect 31330 16158 31332 16210
rect 31276 15540 31332 16158
rect 31388 16098 31444 16604
rect 31612 16594 31668 16604
rect 31388 16046 31390 16098
rect 31442 16046 31444 16098
rect 31388 16034 31444 16046
rect 32508 15876 32564 16828
rect 33068 16818 33124 16828
rect 33180 16660 33236 19852
rect 33516 19346 33572 19358
rect 33516 19294 33518 19346
rect 33570 19294 33572 19346
rect 33516 18452 33572 19294
rect 33516 18386 33572 18396
rect 33964 18452 34020 20132
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 34636 19124 34692 19134
rect 34524 18562 34580 18574
rect 34524 18510 34526 18562
rect 34578 18510 34580 18562
rect 34300 18452 34356 18462
rect 33964 18450 34356 18452
rect 33964 18398 33966 18450
rect 34018 18398 34302 18450
rect 34354 18398 34356 18450
rect 33964 18396 34356 18398
rect 33964 18386 34020 18396
rect 34300 18386 34356 18396
rect 34524 18452 34580 18510
rect 34524 18386 34580 18396
rect 34636 18338 34692 19068
rect 35644 19124 35700 19134
rect 35644 19030 35700 19068
rect 34636 18286 34638 18338
rect 34690 18286 34692 18338
rect 34636 18274 34692 18286
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 33068 16604 33236 16660
rect 34188 17668 34244 17678
rect 35756 17668 35812 17678
rect 32732 15876 32788 15886
rect 32508 15810 32564 15820
rect 32620 15820 32732 15876
rect 31276 15484 31780 15540
rect 31724 15426 31780 15484
rect 31724 15374 31726 15426
rect 31778 15374 31780 15426
rect 31724 15362 31780 15374
rect 32508 15316 32564 15326
rect 32620 15316 32676 15820
rect 32732 15810 32788 15820
rect 32508 15314 32676 15316
rect 32508 15262 32510 15314
rect 32562 15262 32676 15314
rect 32508 15260 32676 15262
rect 32508 15250 32564 15260
rect 31948 14644 32004 14654
rect 31948 14550 32004 14588
rect 32956 14644 33012 14654
rect 33068 14644 33124 16604
rect 33852 15988 33908 15998
rect 33852 15894 33908 15932
rect 33180 15876 33236 15886
rect 33180 15538 33236 15820
rect 33180 15486 33182 15538
rect 33234 15486 33236 15538
rect 33180 15474 33236 15486
rect 34188 15314 34244 17612
rect 35308 17666 35812 17668
rect 35308 17614 35758 17666
rect 35810 17614 35812 17666
rect 35308 17612 35812 17614
rect 35196 17556 35252 17566
rect 34972 17554 35252 17556
rect 34972 17502 35198 17554
rect 35250 17502 35252 17554
rect 34972 17500 35252 17502
rect 34972 17444 35028 17500
rect 35196 17490 35252 17500
rect 35308 17554 35364 17612
rect 35756 17602 35812 17612
rect 35308 17502 35310 17554
rect 35362 17502 35364 17554
rect 34860 16324 34916 16334
rect 34972 16324 35028 17388
rect 35308 16884 35364 17502
rect 35868 17554 35924 17566
rect 35868 17502 35870 17554
rect 35922 17502 35924 17554
rect 35532 17442 35588 17454
rect 35532 17390 35534 17442
rect 35586 17390 35588 17442
rect 35532 16996 35588 17390
rect 35868 16996 35924 17502
rect 35532 16930 35588 16940
rect 35644 16940 35924 16996
rect 34860 16322 35028 16324
rect 34860 16270 34862 16322
rect 34914 16270 35028 16322
rect 34860 16268 35028 16270
rect 35084 16828 35364 16884
rect 34860 16258 34916 16268
rect 34412 16100 34468 16110
rect 34412 16006 34468 16044
rect 34300 15988 34356 15998
rect 34300 15894 34356 15932
rect 34524 15988 34580 15998
rect 34972 15988 35028 15998
rect 34524 15986 35028 15988
rect 34524 15934 34526 15986
rect 34578 15934 34974 15986
rect 35026 15934 35028 15986
rect 34524 15932 35028 15934
rect 34524 15922 34580 15932
rect 34188 15262 34190 15314
rect 34242 15262 34244 15314
rect 34188 15250 34244 15262
rect 34972 14756 35028 15932
rect 35084 15986 35140 16828
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35084 15934 35086 15986
rect 35138 15934 35140 15986
rect 35084 15922 35140 15934
rect 35644 16324 35700 16940
rect 35420 15428 35476 15438
rect 35644 15428 35700 16268
rect 35868 16660 35924 16670
rect 35868 16210 35924 16604
rect 35868 16158 35870 16210
rect 35922 16158 35924 16210
rect 35868 16146 35924 16158
rect 35980 15538 36036 21532
rect 36428 21586 36484 21598
rect 36428 21534 36430 21586
rect 36482 21534 36484 21586
rect 36428 19234 36484 21534
rect 39228 21474 39284 23100
rect 39452 23062 39508 23100
rect 39676 23154 39732 23324
rect 39676 23102 39678 23154
rect 39730 23102 39732 23154
rect 39676 23090 39732 23102
rect 40068 23324 40516 23380
rect 40012 22484 40068 23324
rect 41132 23156 41188 25228
rect 41916 25060 41972 25342
rect 41356 25004 41972 25060
rect 41356 24946 41412 25004
rect 41356 24894 41358 24946
rect 41410 24894 41412 24946
rect 41356 24882 41412 24894
rect 42028 24836 42084 25564
rect 44044 25526 44100 25564
rect 41804 24780 42084 24836
rect 41244 24722 41300 24734
rect 41244 24670 41246 24722
rect 41298 24670 41300 24722
rect 41244 23604 41300 24670
rect 41580 24724 41636 24734
rect 41580 24722 41748 24724
rect 41580 24670 41582 24722
rect 41634 24670 41748 24722
rect 41580 24668 41748 24670
rect 41580 24658 41636 24668
rect 41244 23548 41636 23604
rect 40908 23154 41188 23156
rect 40908 23102 41134 23154
rect 41186 23102 41188 23154
rect 40908 23100 41188 23102
rect 40348 23044 40404 23054
rect 40348 23042 40852 23044
rect 40348 22990 40350 23042
rect 40402 22990 40852 23042
rect 40348 22988 40852 22990
rect 40348 22978 40404 22988
rect 40796 22594 40852 22988
rect 40796 22542 40798 22594
rect 40850 22542 40852 22594
rect 40796 22530 40852 22542
rect 40012 22390 40068 22428
rect 40572 22372 40628 22382
rect 40908 22372 40964 23100
rect 41132 23090 41188 23100
rect 41468 23378 41524 23390
rect 41468 23326 41470 23378
rect 41522 23326 41524 23378
rect 41244 22930 41300 22942
rect 41244 22878 41246 22930
rect 41298 22878 41300 22930
rect 41132 22596 41188 22606
rect 41244 22596 41300 22878
rect 41132 22594 41300 22596
rect 41132 22542 41134 22594
rect 41186 22542 41300 22594
rect 41132 22540 41300 22542
rect 41132 22530 41188 22540
rect 40572 22370 40964 22372
rect 40572 22318 40574 22370
rect 40626 22318 40964 22370
rect 40572 22316 40964 22318
rect 41020 22484 41076 22494
rect 40572 22306 40628 22316
rect 41020 22258 41076 22428
rect 41020 22206 41022 22258
rect 41074 22206 41076 22258
rect 41020 22194 41076 22206
rect 39228 21422 39230 21474
rect 39282 21422 39284 21474
rect 39228 21410 39284 21422
rect 39788 21474 39844 21486
rect 39788 21422 39790 21474
rect 39842 21422 39844 21474
rect 36428 19182 36430 19234
rect 36482 19182 36484 19234
rect 36428 19012 36484 19182
rect 37100 20244 37156 20254
rect 37100 19012 37156 20188
rect 39788 20244 39844 21422
rect 41468 20914 41524 23326
rect 41580 23154 41636 23548
rect 41692 23492 41748 24668
rect 41692 23426 41748 23436
rect 41804 23716 41860 24780
rect 41804 23266 41860 23660
rect 41804 23214 41806 23266
rect 41858 23214 41860 23266
rect 41804 23202 41860 23214
rect 41580 23102 41582 23154
rect 41634 23102 41636 23154
rect 41580 21812 41636 23102
rect 41580 21746 41636 21756
rect 42588 21812 42644 21822
rect 42588 21718 42644 21756
rect 42700 21476 42756 21486
rect 42700 21474 43652 21476
rect 42700 21422 42702 21474
rect 42754 21422 43652 21474
rect 42700 21420 43652 21422
rect 42700 21410 42756 21420
rect 41468 20862 41470 20914
rect 41522 20862 41524 20914
rect 41468 20850 41524 20862
rect 43596 20914 43652 21420
rect 43596 20862 43598 20914
rect 43650 20862 43652 20914
rect 43596 20850 43652 20862
rect 40684 20802 40740 20814
rect 40684 20750 40686 20802
rect 40738 20750 40740 20802
rect 39788 20178 39844 20188
rect 40348 20580 40404 20590
rect 40684 20580 40740 20750
rect 40348 20578 40740 20580
rect 40348 20526 40350 20578
rect 40402 20526 40740 20578
rect 40348 20524 40740 20526
rect 40348 20244 40404 20524
rect 40348 20178 40404 20188
rect 36428 19010 37156 19012
rect 36428 18958 37102 19010
rect 37154 18958 37156 19010
rect 36428 18956 37156 18958
rect 36428 17556 36484 17566
rect 36428 16322 36484 17500
rect 36876 16772 36932 18956
rect 37100 18946 37156 18956
rect 36988 17556 37044 17566
rect 36988 17462 37044 17500
rect 37324 17442 37380 17454
rect 37324 17390 37326 17442
rect 37378 17390 37380 17442
rect 37100 16772 37156 16782
rect 36876 16770 37156 16772
rect 36876 16718 37102 16770
rect 37154 16718 37156 16770
rect 36876 16716 37156 16718
rect 36428 16270 36430 16322
rect 36482 16270 36484 16322
rect 36428 16258 36484 16270
rect 36092 16100 36148 16110
rect 36092 16006 36148 16044
rect 35980 15486 35982 15538
rect 36034 15486 36036 15538
rect 35980 15474 36036 15486
rect 37100 15876 37156 16716
rect 37324 16212 37380 17390
rect 37324 16146 37380 16156
rect 37436 16324 37492 16334
rect 37436 16210 37492 16268
rect 37436 16158 37438 16210
rect 37490 16158 37492 16210
rect 37436 16146 37492 16158
rect 39564 16212 39620 16222
rect 39564 16118 39620 16156
rect 36876 15428 36932 15438
rect 35420 15426 35700 15428
rect 35420 15374 35422 15426
rect 35474 15374 35700 15426
rect 35420 15372 35700 15374
rect 36764 15426 36932 15428
rect 36764 15374 36878 15426
rect 36930 15374 36932 15426
rect 36764 15372 36932 15374
rect 35420 15362 35476 15372
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 34972 14700 35700 14756
rect 33012 14588 33124 14644
rect 32956 14578 33012 14588
rect 35420 13972 35476 13982
rect 35420 13878 35476 13916
rect 35644 13970 35700 14700
rect 35644 13918 35646 13970
rect 35698 13918 35700 13970
rect 34972 13746 35028 13758
rect 34972 13694 34974 13746
rect 35026 13694 35028 13746
rect 34748 13636 34804 13646
rect 34972 13636 35028 13694
rect 35644 13748 35700 13918
rect 36540 13972 36596 13982
rect 36764 13972 36820 15372
rect 36876 15362 36932 15372
rect 36596 13916 37044 13972
rect 35644 13682 35700 13692
rect 36316 13748 36372 13758
rect 36316 13654 36372 13692
rect 36540 13746 36596 13916
rect 36540 13694 36542 13746
rect 36594 13694 36596 13746
rect 36540 13682 36596 13694
rect 34804 13580 35028 13636
rect 35532 13634 35588 13646
rect 35532 13582 35534 13634
rect 35586 13582 35588 13634
rect 34524 11508 34580 11518
rect 34748 11508 34804 13580
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35532 13300 35588 13582
rect 35980 13522 36036 13534
rect 35980 13470 35982 13522
rect 36034 13470 36036 13522
rect 35532 13244 35924 13300
rect 35868 13186 35924 13244
rect 35868 13134 35870 13186
rect 35922 13134 35924 13186
rect 35868 13122 35924 13134
rect 35980 12852 36036 13470
rect 36092 13076 36148 13086
rect 36092 12982 36148 13020
rect 36988 13074 37044 13916
rect 36988 13022 36990 13074
rect 37042 13022 37044 13074
rect 36988 13010 37044 13022
rect 36092 12852 36148 12862
rect 35532 12850 36148 12852
rect 35532 12798 36094 12850
rect 36146 12798 36148 12850
rect 35532 12796 36148 12798
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 34524 11506 34804 11508
rect 34524 11454 34526 11506
rect 34578 11454 34804 11506
rect 34524 11452 34804 11454
rect 34524 11442 34580 11452
rect 34748 11394 34804 11452
rect 35420 11396 35476 11406
rect 35532 11396 35588 12796
rect 36092 12786 36148 12796
rect 36652 12066 36708 12078
rect 36652 12014 36654 12066
rect 36706 12014 36708 12066
rect 36652 11956 36708 12014
rect 36988 11956 37044 11966
rect 37100 11956 37156 15820
rect 40348 16098 40404 16110
rect 40348 16046 40350 16098
rect 40402 16046 40404 16098
rect 40348 15876 40404 16046
rect 40348 15810 40404 15820
rect 36652 11900 36988 11956
rect 37044 11900 37156 11956
rect 37996 15314 38052 15326
rect 37996 15262 37998 15314
rect 38050 15262 38052 15314
rect 34748 11342 34750 11394
rect 34802 11342 34804 11394
rect 34748 11330 34804 11342
rect 34860 11394 35588 11396
rect 34860 11342 35422 11394
rect 35474 11342 35588 11394
rect 34860 11340 35588 11342
rect 31724 10836 31780 10846
rect 31724 10742 31780 10780
rect 34860 10610 34916 11340
rect 35420 11330 35476 11340
rect 35196 11172 35252 11182
rect 34860 10558 34862 10610
rect 34914 10558 34916 10610
rect 34860 10546 34916 10558
rect 35084 11116 35196 11172
rect 35084 10610 35140 11116
rect 35196 11078 35252 11116
rect 35308 11170 35364 11182
rect 35308 11118 35310 11170
rect 35362 11118 35364 11170
rect 35308 10724 35364 11118
rect 35420 10724 35476 10734
rect 35308 10722 35476 10724
rect 35308 10670 35422 10722
rect 35474 10670 35476 10722
rect 35308 10668 35476 10670
rect 35420 10658 35476 10668
rect 35644 10722 35700 10734
rect 35644 10670 35646 10722
rect 35698 10670 35700 10722
rect 35084 10558 35086 10610
rect 35138 10558 35140 10610
rect 35084 10546 35140 10558
rect 31276 10498 31332 10510
rect 31276 10446 31278 10498
rect 31330 10446 31332 10498
rect 31052 9940 31108 9950
rect 31276 9940 31332 10446
rect 35532 10498 35588 10510
rect 35532 10446 35534 10498
rect 35586 10446 35588 10498
rect 34524 10386 34580 10398
rect 34524 10334 34526 10386
rect 34578 10334 34580 10386
rect 31388 10052 31444 10062
rect 31388 9958 31444 9996
rect 31108 9884 31332 9940
rect 32060 9940 32116 9950
rect 31052 9826 31108 9884
rect 31052 9774 31054 9826
rect 31106 9774 31108 9826
rect 31052 9762 31108 9774
rect 31836 9828 31892 9838
rect 31836 9734 31892 9772
rect 32060 9828 32116 9884
rect 33964 9828 34020 9838
rect 32060 9826 32340 9828
rect 32060 9774 32062 9826
rect 32114 9774 32340 9826
rect 32060 9772 32340 9774
rect 32060 9762 32116 9772
rect 30828 9716 30884 9726
rect 30828 9622 30884 9660
rect 31948 9716 32004 9726
rect 31948 9622 32004 9660
rect 31388 9604 31444 9614
rect 31388 9268 31444 9548
rect 32284 9380 32340 9772
rect 33964 9734 34020 9772
rect 34524 9828 34580 10334
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 34524 9762 34580 9772
rect 33740 9716 33796 9726
rect 32284 9324 32452 9380
rect 31388 9266 31668 9268
rect 31388 9214 31390 9266
rect 31442 9214 31668 9266
rect 31388 9212 31668 9214
rect 31388 9202 31444 9212
rect 31612 9042 31668 9212
rect 31612 8990 31614 9042
rect 31666 8990 31668 9042
rect 31612 8978 31668 8990
rect 32060 9156 32116 9166
rect 30716 8372 30884 8428
rect 30828 6466 30884 8372
rect 32060 7698 32116 9100
rect 32284 9044 32340 9054
rect 32284 8950 32340 8988
rect 32172 8932 32228 8942
rect 32172 8838 32228 8876
rect 32396 8428 32452 9324
rect 33292 9156 33348 9166
rect 33292 9062 33348 9100
rect 33068 9042 33124 9054
rect 33068 8990 33070 9042
rect 33122 8990 33124 9042
rect 32844 8932 32900 8942
rect 33068 8932 33124 8990
rect 33740 9044 33796 9660
rect 35532 9154 35588 10446
rect 35644 9716 35700 10670
rect 35644 9650 35700 9660
rect 35532 9102 35534 9154
rect 35586 9102 35588 9154
rect 35532 9090 35588 9102
rect 33740 8950 33796 8988
rect 34860 9042 34916 9054
rect 34860 8990 34862 9042
rect 34914 8990 34916 9042
rect 32900 8876 33124 8932
rect 33516 8930 33572 8942
rect 33516 8878 33518 8930
rect 33570 8878 33572 8930
rect 32844 8866 32900 8876
rect 32060 7646 32062 7698
rect 32114 7646 32116 7698
rect 32060 7634 32116 7646
rect 32284 8372 32452 8428
rect 32284 6580 32340 8372
rect 32396 7474 32452 7486
rect 32396 7422 32398 7474
rect 32450 7422 32452 7474
rect 32396 6916 32452 7422
rect 33516 6916 33572 8878
rect 32396 6860 32788 6916
rect 32620 6692 32676 6702
rect 32396 6580 32452 6590
rect 32284 6578 32452 6580
rect 32284 6526 32398 6578
rect 32450 6526 32452 6578
rect 32284 6524 32452 6526
rect 32396 6514 32452 6524
rect 30828 6414 30830 6466
rect 30882 6414 30884 6466
rect 30828 6402 30884 6414
rect 31164 6132 31220 6142
rect 30604 6130 31220 6132
rect 30604 6078 31166 6130
rect 31218 6078 31220 6130
rect 30604 6076 31220 6078
rect 28812 6018 29204 6020
rect 28812 5966 28814 6018
rect 28866 5966 29150 6018
rect 29202 5966 29204 6018
rect 28812 5964 29204 5966
rect 28812 5954 28868 5964
rect 29148 5954 29204 5964
rect 30268 6020 30324 6076
rect 30268 5954 30324 5964
rect 28476 5906 28532 5918
rect 28476 5854 28478 5906
rect 28530 5854 28532 5906
rect 28476 5796 28532 5854
rect 29372 5908 29428 5918
rect 28476 5730 28532 5740
rect 29260 5796 29316 5806
rect 29260 5702 29316 5740
rect 29372 5572 29428 5852
rect 29596 5908 29652 5918
rect 29596 5814 29652 5852
rect 30156 5908 30212 5918
rect 30156 5814 30212 5852
rect 30604 5906 30660 6076
rect 31164 6066 31220 6076
rect 30604 5854 30606 5906
rect 30658 5854 30660 5906
rect 30604 5842 30660 5854
rect 27804 5182 27806 5234
rect 27858 5182 27860 5234
rect 27356 5170 27412 5180
rect 27804 5170 27860 5182
rect 29148 5516 29428 5572
rect 31276 5796 31332 5806
rect 29148 5234 29204 5516
rect 29148 5182 29150 5234
rect 29202 5182 29204 5234
rect 29148 5170 29204 5182
rect 31276 5234 31332 5740
rect 31276 5182 31278 5234
rect 31330 5182 31332 5234
rect 31276 5170 31332 5182
rect 32620 5234 32676 6636
rect 32732 5796 32788 6860
rect 33516 6850 33572 6860
rect 34860 8484 34916 8990
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 33516 6690 33572 6702
rect 33516 6638 33518 6690
rect 33570 6638 33572 6690
rect 33068 5796 33124 5806
rect 33516 5796 33572 6638
rect 34860 6692 34916 8428
rect 36428 8484 36484 8494
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 34860 6626 34916 6636
rect 35196 6916 35252 6926
rect 35196 6018 35252 6860
rect 36428 6132 36484 8428
rect 36988 8484 37044 11900
rect 37660 11172 37716 11182
rect 37660 8930 37716 11116
rect 37996 11172 38052 15262
rect 39116 13076 39172 13086
rect 39116 12982 39172 13020
rect 39788 12962 39844 12974
rect 39788 12910 39790 12962
rect 39842 12910 39844 12962
rect 39788 11956 39844 12910
rect 39788 11890 39844 11900
rect 37996 11106 38052 11116
rect 37660 8878 37662 8930
rect 37714 8878 37716 8930
rect 37660 8866 37716 8878
rect 38108 8930 38164 8942
rect 38108 8878 38110 8930
rect 38162 8878 38164 8930
rect 36988 8418 37044 8428
rect 38108 8484 38164 8878
rect 38108 8418 38164 8428
rect 35196 5966 35198 6018
rect 35250 5966 35252 6018
rect 35196 5954 35252 5966
rect 35980 6130 36484 6132
rect 35980 6078 36430 6130
rect 36482 6078 36484 6130
rect 35980 6076 36484 6078
rect 35980 5906 36036 6076
rect 36428 6066 36484 6076
rect 35980 5854 35982 5906
rect 36034 5854 36036 5906
rect 35980 5842 36036 5854
rect 32732 5794 33572 5796
rect 32732 5742 33070 5794
rect 33122 5742 33572 5794
rect 32732 5740 33572 5742
rect 33068 5730 33124 5740
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 32620 5182 32622 5234
rect 32674 5182 32676 5234
rect 24556 5070 24558 5122
rect 24610 5070 24612 5122
rect 24556 5058 24612 5070
rect 31948 5124 32004 5134
rect 31948 5030 32004 5068
rect 32620 5124 32676 5182
rect 32620 5058 32676 5068
rect 21756 4398 21758 4450
rect 21810 4398 21812 4450
rect 21756 4386 21812 4398
rect 22540 4562 23044 4564
rect 22540 4510 22990 4562
rect 23042 4510 23044 4562
rect 22540 4508 23044 4510
rect 22540 4338 22596 4508
rect 22988 4498 23044 4508
rect 22540 4286 22542 4338
rect 22594 4286 22596 4338
rect 22540 4274 22596 4286
rect 19628 4174 19630 4226
rect 19682 4174 19684 4226
rect 19628 4162 19684 4174
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
<< via2 >>
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 2940 40402 2996 40404
rect 2940 40350 2942 40402
rect 2942 40350 2994 40402
rect 2994 40350 2996 40402
rect 2940 40348 2996 40350
rect 5068 40290 5124 40292
rect 5068 40238 5070 40290
rect 5070 40238 5122 40290
rect 5122 40238 5124 40290
rect 5068 40236 5124 40238
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 2716 38892 2772 38948
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 2268 37772 2324 37828
rect 3052 37772 3108 37828
rect 3724 37378 3780 37380
rect 3724 37326 3726 37378
rect 3726 37326 3778 37378
rect 3778 37326 3780 37378
rect 3724 37324 3780 37326
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 5740 37826 5796 37828
rect 5740 37774 5742 37826
rect 5742 37774 5794 37826
rect 5794 37774 5796 37826
rect 5740 37772 5796 37774
rect 6300 37772 6356 37828
rect 5852 36540 5908 36596
rect 4844 35756 4900 35812
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 2268 31778 2324 31780
rect 2268 31726 2270 31778
rect 2270 31726 2322 31778
rect 2322 31726 2324 31778
rect 2268 31724 2324 31726
rect 2716 31724 2772 31780
rect 8988 40012 9044 40068
rect 8316 39506 8372 39508
rect 8316 39454 8318 39506
rect 8318 39454 8370 39506
rect 8370 39454 8372 39506
rect 8316 39452 8372 39454
rect 7196 39228 7252 39284
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 13244 41804 13300 41860
rect 11564 40514 11620 40516
rect 11564 40462 11566 40514
rect 11566 40462 11618 40514
rect 11618 40462 11620 40514
rect 11564 40460 11620 40462
rect 9772 37826 9828 37828
rect 9772 37774 9774 37826
rect 9774 37774 9826 37826
rect 9826 37774 9828 37826
rect 9772 37772 9828 37774
rect 10332 38780 10388 38836
rect 10332 37378 10388 37380
rect 10332 37326 10334 37378
rect 10334 37326 10386 37378
rect 10386 37326 10388 37378
rect 10332 37324 10388 37326
rect 6524 36764 6580 36820
rect 6972 36594 7028 36596
rect 6972 36542 6974 36594
rect 6974 36542 7026 36594
rect 7026 36542 7028 36594
rect 6972 36540 7028 36542
rect 9996 36540 10052 36596
rect 7084 36258 7140 36260
rect 7084 36206 7086 36258
rect 7086 36206 7138 36258
rect 7138 36206 7140 36258
rect 7084 36204 7140 36206
rect 10220 36204 10276 36260
rect 10332 35308 10388 35364
rect 6636 33458 6692 33460
rect 6636 33406 6638 33458
rect 6638 33406 6690 33458
rect 6690 33406 6692 33458
rect 6636 33404 6692 33406
rect 8988 33404 9044 33460
rect 11340 40402 11396 40404
rect 11340 40350 11342 40402
rect 11342 40350 11394 40402
rect 11394 40350 11396 40402
rect 11340 40348 11396 40350
rect 12012 40460 12068 40516
rect 11676 40402 11732 40404
rect 11676 40350 11678 40402
rect 11678 40350 11730 40402
rect 11730 40350 11732 40402
rect 11676 40348 11732 40350
rect 12348 40514 12404 40516
rect 12348 40462 12350 40514
rect 12350 40462 12402 40514
rect 12402 40462 12404 40514
rect 12348 40460 12404 40462
rect 12124 40348 12180 40404
rect 12460 40290 12516 40292
rect 12460 40238 12462 40290
rect 12462 40238 12514 40290
rect 12514 40238 12516 40290
rect 12460 40236 12516 40238
rect 11004 39618 11060 39620
rect 11004 39566 11006 39618
rect 11006 39566 11058 39618
rect 11058 39566 11060 39618
rect 11004 39564 11060 39566
rect 14476 41858 14532 41860
rect 14476 41806 14478 41858
rect 14478 41806 14530 41858
rect 14530 41806 14532 41858
rect 14476 41804 14532 41806
rect 13468 40124 13524 40180
rect 13916 40348 13972 40404
rect 12572 39564 12628 39620
rect 12684 39452 12740 39508
rect 10668 39394 10724 39396
rect 10668 39342 10670 39394
rect 10670 39342 10722 39394
rect 10722 39342 10724 39394
rect 10668 39340 10724 39342
rect 11900 39228 11956 39284
rect 11676 38892 11732 38948
rect 12012 39004 12068 39060
rect 12572 38946 12628 38948
rect 12572 38894 12574 38946
rect 12574 38894 12626 38946
rect 12626 38894 12628 38946
rect 12572 38892 12628 38894
rect 14252 39618 14308 39620
rect 14252 39566 14254 39618
rect 14254 39566 14306 39618
rect 14306 39566 14308 39618
rect 14252 39564 14308 39566
rect 14028 39506 14084 39508
rect 14028 39454 14030 39506
rect 14030 39454 14082 39506
rect 14082 39454 14084 39506
rect 14028 39452 14084 39454
rect 13804 38834 13860 38836
rect 13804 38782 13806 38834
rect 13806 38782 13858 38834
rect 13858 38782 13860 38834
rect 13804 38780 13860 38782
rect 14028 38834 14084 38836
rect 14028 38782 14030 38834
rect 14030 38782 14082 38834
rect 14082 38782 14084 38834
rect 14028 38780 14084 38782
rect 11004 36988 11060 37044
rect 11228 37266 11284 37268
rect 11228 37214 11230 37266
rect 11230 37214 11282 37266
rect 11282 37214 11284 37266
rect 11228 37212 11284 37214
rect 11564 37100 11620 37156
rect 11788 37212 11844 37268
rect 12236 37212 12292 37268
rect 11676 36988 11732 37044
rect 12460 37100 12516 37156
rect 12348 36988 12404 37044
rect 12012 36764 12068 36820
rect 13468 36764 13524 36820
rect 12348 36594 12404 36596
rect 12348 36542 12350 36594
rect 12350 36542 12402 36594
rect 12402 36542 12404 36594
rect 12348 36540 12404 36542
rect 12908 36594 12964 36596
rect 12908 36542 12910 36594
rect 12910 36542 12962 36594
rect 12962 36542 12964 36594
rect 12908 36540 12964 36542
rect 12572 36482 12628 36484
rect 12572 36430 12574 36482
rect 12574 36430 12626 36482
rect 12626 36430 12628 36482
rect 12572 36428 12628 36430
rect 13244 36428 13300 36484
rect 13020 35810 13076 35812
rect 13020 35758 13022 35810
rect 13022 35758 13074 35810
rect 13074 35758 13076 35810
rect 13020 35756 13076 35758
rect 14364 39452 14420 39508
rect 14700 40124 14756 40180
rect 16940 40514 16996 40516
rect 16940 40462 16942 40514
rect 16942 40462 16994 40514
rect 16994 40462 16996 40514
rect 16940 40460 16996 40462
rect 15484 40124 15540 40180
rect 16044 39730 16100 39732
rect 16044 39678 16046 39730
rect 16046 39678 16098 39730
rect 16098 39678 16100 39730
rect 16044 39676 16100 39678
rect 15596 39618 15652 39620
rect 15596 39566 15598 39618
rect 15598 39566 15650 39618
rect 15650 39566 15652 39618
rect 15596 39564 15652 39566
rect 14812 39452 14868 39508
rect 14588 39394 14644 39396
rect 14588 39342 14590 39394
rect 14590 39342 14642 39394
rect 14642 39342 14644 39394
rect 14588 39340 14644 39342
rect 14476 37100 14532 37156
rect 14588 36988 14644 37044
rect 13468 36482 13524 36484
rect 13468 36430 13470 36482
rect 13470 36430 13522 36482
rect 13522 36430 13524 36482
rect 13468 36428 13524 36430
rect 13804 36540 13860 36596
rect 13692 36370 13748 36372
rect 13692 36318 13694 36370
rect 13694 36318 13746 36370
rect 13746 36318 13748 36370
rect 13692 36316 13748 36318
rect 15148 39228 15204 39284
rect 14924 38892 14980 38948
rect 15820 39452 15876 39508
rect 15036 38834 15092 38836
rect 15036 38782 15038 38834
rect 15038 38782 15090 38834
rect 15090 38782 15092 38834
rect 15036 38780 15092 38782
rect 15708 39058 15764 39060
rect 15708 39006 15710 39058
rect 15710 39006 15762 39058
rect 15762 39006 15764 39058
rect 15708 39004 15764 39006
rect 15596 38780 15652 38836
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 17276 40012 17332 40068
rect 17836 40348 17892 40404
rect 20076 40402 20132 40404
rect 20076 40350 20078 40402
rect 20078 40350 20130 40402
rect 20130 40350 20132 40402
rect 20076 40348 20132 40350
rect 23212 41916 23268 41972
rect 21420 40348 21476 40404
rect 21084 40290 21140 40292
rect 21084 40238 21086 40290
rect 21086 40238 21138 40290
rect 21138 40238 21140 40290
rect 21084 40236 21140 40238
rect 28476 42140 28532 42196
rect 24892 41970 24948 41972
rect 24892 41918 24894 41970
rect 24894 41918 24946 41970
rect 24946 41918 24948 41970
rect 24892 41916 24948 41918
rect 24668 41804 24724 41860
rect 25900 41858 25956 41860
rect 25900 41806 25902 41858
rect 25902 41806 25954 41858
rect 25954 41806 25956 41858
rect 25900 41804 25956 41806
rect 25340 40402 25396 40404
rect 25340 40350 25342 40402
rect 25342 40350 25394 40402
rect 25394 40350 25396 40402
rect 25340 40348 25396 40350
rect 16828 39506 16884 39508
rect 16828 39454 16830 39506
rect 16830 39454 16882 39506
rect 16882 39454 16884 39506
rect 16828 39452 16884 39454
rect 16380 39394 16436 39396
rect 16380 39342 16382 39394
rect 16382 39342 16434 39394
rect 16434 39342 16436 39394
rect 16380 39340 16436 39342
rect 16940 39394 16996 39396
rect 16940 39342 16942 39394
rect 16942 39342 16994 39394
rect 16994 39342 16996 39394
rect 16940 39340 16996 39342
rect 16156 39228 16212 39284
rect 17052 39228 17108 39284
rect 15932 39004 15988 39060
rect 18620 39618 18676 39620
rect 18620 39566 18622 39618
rect 18622 39566 18674 39618
rect 18674 39566 18676 39618
rect 18620 39564 18676 39566
rect 30380 41970 30436 41972
rect 30380 41918 30382 41970
rect 30382 41918 30434 41970
rect 30434 41918 30436 41970
rect 30380 41916 30436 41918
rect 31388 41916 31444 41972
rect 28588 40402 28644 40404
rect 28588 40350 28590 40402
rect 28590 40350 28642 40402
rect 28642 40350 28644 40402
rect 28588 40348 28644 40350
rect 26012 39340 26068 39396
rect 32508 41970 32564 41972
rect 32508 41918 32510 41970
rect 32510 41918 32562 41970
rect 32562 41918 32564 41970
rect 32508 41916 32564 41918
rect 33740 41916 33796 41972
rect 31612 40460 31668 40516
rect 29260 39676 29316 39732
rect 28364 39618 28420 39620
rect 28364 39566 28366 39618
rect 28366 39566 28418 39618
rect 28418 39566 28420 39618
rect 28364 39564 28420 39566
rect 30268 39564 30324 39620
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 15596 36540 15652 36596
rect 15036 36428 15092 36484
rect 15484 36482 15540 36484
rect 15484 36430 15486 36482
rect 15486 36430 15538 36482
rect 15538 36430 15540 36482
rect 15484 36428 15540 36430
rect 16716 37154 16772 37156
rect 16716 37102 16718 37154
rect 16718 37102 16770 37154
rect 16770 37102 16772 37154
rect 16716 37100 16772 37102
rect 16268 36316 16324 36372
rect 13244 35698 13300 35700
rect 13244 35646 13246 35698
rect 13246 35646 13298 35698
rect 13298 35646 13300 35698
rect 13244 35644 13300 35646
rect 13916 35644 13972 35700
rect 14252 35308 14308 35364
rect 14700 35308 14756 35364
rect 15036 35532 15092 35588
rect 16716 35420 16772 35476
rect 14812 34802 14868 34804
rect 14812 34750 14814 34802
rect 14814 34750 14866 34802
rect 14866 34750 14868 34802
rect 14812 34748 14868 34750
rect 8988 32732 9044 32788
rect 8428 32674 8484 32676
rect 8428 32622 8430 32674
rect 8430 32622 8482 32674
rect 8482 32622 8484 32674
rect 8428 32620 8484 32622
rect 9772 32786 9828 32788
rect 9772 32734 9774 32786
rect 9774 32734 9826 32786
rect 9826 32734 9828 32786
rect 9772 32732 9828 32734
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 3388 30828 3444 30884
rect 4956 30828 5012 30884
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 3388 29372 3444 29428
rect 3276 28924 3332 28980
rect 3164 28642 3220 28644
rect 3164 28590 3166 28642
rect 3166 28590 3218 28642
rect 3218 28590 3220 28642
rect 3164 28588 3220 28590
rect 3612 28588 3668 28644
rect 3500 28530 3556 28532
rect 3500 28478 3502 28530
rect 3502 28478 3554 28530
rect 3554 28478 3556 28530
rect 3500 28476 3556 28478
rect 2940 25228 2996 25284
rect 3164 24444 3220 24500
rect 2268 23938 2324 23940
rect 2268 23886 2270 23938
rect 2270 23886 2322 23938
rect 2322 23886 2324 23938
rect 2268 23884 2324 23886
rect 2492 23154 2548 23156
rect 2492 23102 2494 23154
rect 2494 23102 2546 23154
rect 2546 23102 2548 23154
rect 2492 23100 2548 23102
rect 1820 22092 1876 22148
rect 1820 18508 1876 18564
rect 3836 28924 3892 28980
rect 4620 29426 4676 29428
rect 4620 29374 4622 29426
rect 4622 29374 4674 29426
rect 4674 29374 4676 29426
rect 4620 29372 4676 29374
rect 4396 29148 4452 29204
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4060 28700 4116 28756
rect 4284 28476 4340 28532
rect 4396 28812 4452 28868
rect 4508 28642 4564 28644
rect 4508 28590 4510 28642
rect 4510 28590 4562 28642
rect 4562 28590 4564 28642
rect 4508 28588 4564 28590
rect 4732 28642 4788 28644
rect 4732 28590 4734 28642
rect 4734 28590 4786 28642
rect 4786 28590 4788 28642
rect 4732 28588 4788 28590
rect 4508 28364 4564 28420
rect 3724 27804 3780 27860
rect 5068 28924 5124 28980
rect 5628 29372 5684 29428
rect 5740 31052 5796 31108
rect 5068 28476 5124 28532
rect 4956 28364 5012 28420
rect 5628 28418 5684 28420
rect 5628 28366 5630 28418
rect 5630 28366 5682 28418
rect 5682 28366 5684 28418
rect 5628 28364 5684 28366
rect 4732 27858 4788 27860
rect 4732 27806 4734 27858
rect 4734 27806 4786 27858
rect 4786 27806 4788 27858
rect 4732 27804 4788 27806
rect 4284 27692 4340 27748
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 5292 27692 5348 27748
rect 3836 26684 3892 26740
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 3724 24444 3780 24500
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 5068 24050 5124 24052
rect 5068 23998 5070 24050
rect 5070 23998 5122 24050
rect 5122 23998 5124 24050
rect 5068 23996 5124 23998
rect 5292 23100 5348 23156
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 5964 31724 6020 31780
rect 5964 31052 6020 31108
rect 5852 30156 5908 30212
rect 6636 30380 6692 30436
rect 6076 29314 6132 29316
rect 6076 29262 6078 29314
rect 6078 29262 6130 29314
rect 6130 29262 6132 29314
rect 6076 29260 6132 29262
rect 6300 28924 6356 28980
rect 5964 28642 6020 28644
rect 5964 28590 5966 28642
rect 5966 28590 6018 28642
rect 6018 28590 6020 28642
rect 5964 28588 6020 28590
rect 6412 28866 6468 28868
rect 6412 28814 6414 28866
rect 6414 28814 6466 28866
rect 6466 28814 6468 28866
rect 6412 28812 6468 28814
rect 6524 28530 6580 28532
rect 6524 28478 6526 28530
rect 6526 28478 6578 28530
rect 6578 28478 6580 28530
rect 6524 28476 6580 28478
rect 5964 28364 6020 28420
rect 5964 27804 6020 27860
rect 5740 25282 5796 25284
rect 5740 25230 5742 25282
rect 5742 25230 5794 25282
rect 5794 25230 5796 25282
rect 5740 25228 5796 25230
rect 8092 30380 8148 30436
rect 8764 30434 8820 30436
rect 8764 30382 8766 30434
rect 8766 30382 8818 30434
rect 8818 30382 8820 30434
rect 8764 30380 8820 30382
rect 10444 32620 10500 32676
rect 9996 31836 10052 31892
rect 9100 30322 9156 30324
rect 9100 30270 9102 30322
rect 9102 30270 9154 30322
rect 9154 30270 9156 30322
rect 9100 30268 9156 30270
rect 6972 29596 7028 29652
rect 7980 28642 8036 28644
rect 7980 28590 7982 28642
rect 7982 28590 8034 28642
rect 8034 28590 8036 28642
rect 7980 28588 8036 28590
rect 6972 28476 7028 28532
rect 8316 28530 8372 28532
rect 8316 28478 8318 28530
rect 8318 28478 8370 28530
rect 8370 28478 8372 28530
rect 8316 28476 8372 28478
rect 8204 28028 8260 28084
rect 6412 26402 6468 26404
rect 6412 26350 6414 26402
rect 6414 26350 6466 26402
rect 6466 26350 6468 26402
rect 6412 26348 6468 26350
rect 6188 25228 6244 25284
rect 8876 28700 8932 28756
rect 8764 28642 8820 28644
rect 8764 28590 8766 28642
rect 8766 28590 8818 28642
rect 8818 28590 8820 28642
rect 8764 28588 8820 28590
rect 10108 30210 10164 30212
rect 10108 30158 10110 30210
rect 10110 30158 10162 30210
rect 10162 30158 10164 30210
rect 10108 30156 10164 30158
rect 9996 29426 10052 29428
rect 9996 29374 9998 29426
rect 9998 29374 10050 29426
rect 10050 29374 10052 29426
rect 9996 29372 10052 29374
rect 9660 28866 9716 28868
rect 9660 28814 9662 28866
rect 9662 28814 9714 28866
rect 9714 28814 9716 28866
rect 9660 28812 9716 28814
rect 9548 28700 9604 28756
rect 9212 28476 9268 28532
rect 9884 29148 9940 29204
rect 9884 28642 9940 28644
rect 9884 28590 9886 28642
rect 9886 28590 9938 28642
rect 9938 28590 9940 28642
rect 9884 28588 9940 28590
rect 10108 28476 10164 28532
rect 9996 28028 10052 28084
rect 8988 26572 9044 26628
rect 10444 31106 10500 31108
rect 10444 31054 10446 31106
rect 10446 31054 10498 31106
rect 10498 31054 10500 31106
rect 10444 31052 10500 31054
rect 10780 28924 10836 28980
rect 10892 28700 10948 28756
rect 10668 27132 10724 27188
rect 12012 30268 12068 30324
rect 11900 30156 11956 30212
rect 11452 29426 11508 29428
rect 11452 29374 11454 29426
rect 11454 29374 11506 29426
rect 11506 29374 11508 29426
rect 11452 29372 11508 29374
rect 11228 28642 11284 28644
rect 11228 28590 11230 28642
rect 11230 28590 11282 28642
rect 11282 28590 11284 28642
rect 11228 28588 11284 28590
rect 11564 29260 11620 29316
rect 11676 29202 11732 29204
rect 11676 29150 11678 29202
rect 11678 29150 11730 29202
rect 11730 29150 11732 29202
rect 11676 29148 11732 29150
rect 16380 31836 16436 31892
rect 22764 38108 22820 38164
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 18396 36482 18452 36484
rect 18396 36430 18398 36482
rect 18398 36430 18450 36482
rect 18450 36430 18452 36482
rect 18396 36428 18452 36430
rect 19068 36482 19124 36484
rect 19068 36430 19070 36482
rect 19070 36430 19122 36482
rect 19122 36430 19124 36482
rect 19068 36428 19124 36430
rect 17724 36316 17780 36372
rect 17276 35698 17332 35700
rect 17276 35646 17278 35698
rect 17278 35646 17330 35698
rect 17330 35646 17332 35698
rect 17276 35644 17332 35646
rect 18060 35532 18116 35588
rect 18396 35644 18452 35700
rect 20300 37100 20356 37156
rect 19628 36316 19684 36372
rect 19964 36370 20020 36372
rect 19964 36318 19966 36370
rect 19966 36318 20018 36370
rect 20018 36318 20020 36370
rect 19964 36316 20020 36318
rect 20972 36428 21028 36484
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 18844 35474 18900 35476
rect 18844 35422 18846 35474
rect 18846 35422 18898 35474
rect 18898 35422 18900 35474
rect 18844 35420 18900 35422
rect 18620 35138 18676 35140
rect 18620 35086 18622 35138
rect 18622 35086 18674 35138
rect 18674 35086 18676 35138
rect 18620 35084 18676 35086
rect 18396 34802 18452 34804
rect 18396 34750 18398 34802
rect 18398 34750 18450 34802
rect 18450 34750 18452 34802
rect 18396 34748 18452 34750
rect 18956 34690 19012 34692
rect 18956 34638 18958 34690
rect 18958 34638 19010 34690
rect 19010 34638 19012 34690
rect 18956 34636 19012 34638
rect 20300 35756 20356 35812
rect 19180 35084 19236 35140
rect 20076 35698 20132 35700
rect 20076 35646 20078 35698
rect 20078 35646 20130 35698
rect 20130 35646 20132 35698
rect 20076 35644 20132 35646
rect 19852 35084 19908 35140
rect 19516 34802 19572 34804
rect 19516 34750 19518 34802
rect 19518 34750 19570 34802
rect 19570 34750 19572 34802
rect 19516 34748 19572 34750
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19180 34300 19236 34356
rect 20076 34300 20132 34356
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 16828 31890 16884 31892
rect 16828 31838 16830 31890
rect 16830 31838 16882 31890
rect 16882 31838 16884 31890
rect 16828 31836 16884 31838
rect 15484 30994 15540 30996
rect 15484 30942 15486 30994
rect 15486 30942 15538 30994
rect 15538 30942 15540 30994
rect 15484 30940 15540 30942
rect 16492 30940 16548 30996
rect 12124 29484 12180 29540
rect 12012 28530 12068 28532
rect 12012 28478 12014 28530
rect 12014 28478 12066 28530
rect 12066 28478 12068 28530
rect 12012 28476 12068 28478
rect 12572 28642 12628 28644
rect 12572 28590 12574 28642
rect 12574 28590 12626 28642
rect 12626 28590 12628 28642
rect 12572 28588 12628 28590
rect 10892 28082 10948 28084
rect 10892 28030 10894 28082
rect 10894 28030 10946 28082
rect 10946 28030 10948 28082
rect 10892 28028 10948 28030
rect 10780 26684 10836 26740
rect 12124 27804 12180 27860
rect 10108 26348 10164 26404
rect 9772 26236 9828 26292
rect 8316 25564 8372 25620
rect 6748 25282 6804 25284
rect 6748 25230 6750 25282
rect 6750 25230 6802 25282
rect 6802 25230 6804 25282
rect 6748 25228 6804 25230
rect 5852 23938 5908 23940
rect 5852 23886 5854 23938
rect 5854 23886 5906 23938
rect 5906 23886 5908 23938
rect 5852 23884 5908 23886
rect 5404 22316 5460 22372
rect 5852 23042 5908 23044
rect 5852 22990 5854 23042
rect 5854 22990 5906 23042
rect 5906 22990 5908 23042
rect 5852 22988 5908 22990
rect 3612 21868 3668 21924
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 5068 19852 5124 19908
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4732 19346 4788 19348
rect 4732 19294 4734 19346
rect 4734 19294 4786 19346
rect 4786 19294 4788 19346
rect 4732 19292 4788 19294
rect 2604 18396 2660 18452
rect 3948 18338 4004 18340
rect 3948 18286 3950 18338
rect 3950 18286 4002 18338
rect 4002 18286 4004 18338
rect 3948 18284 4004 18286
rect 5852 19852 5908 19908
rect 6412 22876 6468 22932
rect 6412 21868 6468 21924
rect 5068 18508 5124 18564
rect 4844 18338 4900 18340
rect 4844 18286 4846 18338
rect 4846 18286 4898 18338
rect 4898 18286 4900 18338
rect 4844 18284 4900 18286
rect 4284 18226 4340 18228
rect 4284 18174 4286 18226
rect 4286 18174 4338 18226
rect 4338 18174 4340 18226
rect 4284 18172 4340 18174
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4508 17836 4564 17892
rect 5292 18508 5348 18564
rect 6076 19292 6132 19348
rect 5740 18508 5796 18564
rect 6076 18508 6132 18564
rect 5964 18172 6020 18228
rect 5068 16940 5124 16996
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 5852 15932 5908 15988
rect 6076 16940 6132 16996
rect 6188 16828 6244 16884
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 1932 13468 1988 13524
rect 4844 14306 4900 14308
rect 4844 14254 4846 14306
rect 4846 14254 4898 14306
rect 4898 14254 4900 14306
rect 4844 14252 4900 14254
rect 5180 13468 5236 13524
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 2604 13020 2660 13076
rect 5068 12850 5124 12852
rect 5068 12798 5070 12850
rect 5070 12798 5122 12850
rect 5122 12798 5124 12850
rect 5068 12796 5124 12798
rect 4956 12684 5012 12740
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 5068 11788 5124 11844
rect 4684 11732 4740 11734
rect 4844 11676 4900 11732
rect 4396 11394 4452 11396
rect 4396 11342 4398 11394
rect 4398 11342 4450 11394
rect 4450 11342 4452 11394
rect 4396 11340 4452 11342
rect 4172 11282 4228 11284
rect 4172 11230 4174 11282
rect 4174 11230 4226 11282
rect 4226 11230 4228 11282
rect 4172 11228 4228 11230
rect 2604 11116 2660 11172
rect 4284 11170 4340 11172
rect 4284 11118 4286 11170
rect 4286 11118 4338 11170
rect 4338 11118 4340 11170
rect 4284 11116 4340 11118
rect 6188 14306 6244 14308
rect 6188 14254 6190 14306
rect 6190 14254 6242 14306
rect 6242 14254 6244 14306
rect 6188 14252 6244 14254
rect 5964 13468 6020 13524
rect 5740 13074 5796 13076
rect 5740 13022 5742 13074
rect 5742 13022 5794 13074
rect 5794 13022 5796 13074
rect 5740 13020 5796 13022
rect 5852 12850 5908 12852
rect 5852 12798 5854 12850
rect 5854 12798 5906 12850
rect 5906 12798 5908 12850
rect 5852 12796 5908 12798
rect 6076 12962 6132 12964
rect 6076 12910 6078 12962
rect 6078 12910 6130 12962
rect 6130 12910 6132 12962
rect 6076 12908 6132 12910
rect 8204 24780 8260 24836
rect 6860 23996 6916 24052
rect 7308 24050 7364 24052
rect 7308 23998 7310 24050
rect 7310 23998 7362 24050
rect 7362 23998 7364 24050
rect 7308 23996 7364 23998
rect 7420 23714 7476 23716
rect 7420 23662 7422 23714
rect 7422 23662 7474 23714
rect 7474 23662 7476 23714
rect 7420 23660 7476 23662
rect 6860 23100 6916 23156
rect 7644 23100 7700 23156
rect 8876 25618 8932 25620
rect 8876 25566 8878 25618
rect 8878 25566 8930 25618
rect 8930 25566 8932 25618
rect 8876 25564 8932 25566
rect 8988 24332 9044 24388
rect 8428 23660 8484 23716
rect 6748 21308 6804 21364
rect 6748 17388 6804 17444
rect 7420 21586 7476 21588
rect 7420 21534 7422 21586
rect 7422 21534 7474 21586
rect 7474 21534 7476 21586
rect 7420 21532 7476 21534
rect 11116 26236 11172 26292
rect 10780 25676 10836 25732
rect 10556 24332 10612 24388
rect 9324 20578 9380 20580
rect 9324 20526 9326 20578
rect 9326 20526 9378 20578
rect 9378 20526 9380 20578
rect 9324 20524 9380 20526
rect 8540 20130 8596 20132
rect 8540 20078 8542 20130
rect 8542 20078 8594 20130
rect 8594 20078 8596 20130
rect 8540 20076 8596 20078
rect 8876 20018 8932 20020
rect 8876 19966 8878 20018
rect 8878 19966 8930 20018
rect 8930 19966 8932 20018
rect 8876 19964 8932 19966
rect 8428 19292 8484 19348
rect 9996 20748 10052 20804
rect 10220 20076 10276 20132
rect 10892 20802 10948 20804
rect 10892 20750 10894 20802
rect 10894 20750 10946 20802
rect 10946 20750 10948 20802
rect 10892 20748 10948 20750
rect 11788 25506 11844 25508
rect 11788 25454 11790 25506
rect 11790 25454 11842 25506
rect 11842 25454 11844 25506
rect 11788 25452 11844 25454
rect 12572 27356 12628 27412
rect 12684 26796 12740 26852
rect 12796 28476 12852 28532
rect 12236 26348 12292 26404
rect 12236 25730 12292 25732
rect 12236 25678 12238 25730
rect 12238 25678 12290 25730
rect 12290 25678 12292 25730
rect 12236 25676 12292 25678
rect 12684 26290 12740 26292
rect 12684 26238 12686 26290
rect 12686 26238 12738 26290
rect 12738 26238 12740 26290
rect 12684 26236 12740 26238
rect 13916 29372 13972 29428
rect 15932 30044 15988 30100
rect 16044 29932 16100 29988
rect 16828 30828 16884 30884
rect 20748 36316 20804 36372
rect 21756 36316 21812 36372
rect 21756 35756 21812 35812
rect 26012 38162 26068 38164
rect 26012 38110 26014 38162
rect 26014 38110 26066 38162
rect 26066 38110 26068 38162
rect 26012 38108 26068 38110
rect 28364 38108 28420 38164
rect 24556 36652 24612 36708
rect 25564 36706 25620 36708
rect 25564 36654 25566 36706
rect 25566 36654 25618 36706
rect 25618 36654 25620 36706
rect 25564 36652 25620 36654
rect 26460 36652 26516 36708
rect 24108 36370 24164 36372
rect 24108 36318 24110 36370
rect 24110 36318 24162 36370
rect 24162 36318 24164 36370
rect 24108 36316 24164 36318
rect 25228 35698 25284 35700
rect 25228 35646 25230 35698
rect 25230 35646 25282 35698
rect 25282 35646 25284 35698
rect 25228 35644 25284 35646
rect 23436 35420 23492 35476
rect 24220 35420 24276 35476
rect 21644 34860 21700 34916
rect 16492 29932 16548 29988
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 18284 30882 18340 30884
rect 18284 30830 18286 30882
rect 18286 30830 18338 30882
rect 18338 30830 18340 30882
rect 18284 30828 18340 30830
rect 17500 30044 17556 30100
rect 14476 29538 14532 29540
rect 14476 29486 14478 29538
rect 14478 29486 14530 29538
rect 14530 29486 14532 29538
rect 14476 29484 14532 29486
rect 14364 29426 14420 29428
rect 14364 29374 14366 29426
rect 14366 29374 14418 29426
rect 14418 29374 14420 29426
rect 14364 29372 14420 29374
rect 15484 29372 15540 29428
rect 16156 29538 16212 29540
rect 16156 29486 16158 29538
rect 16158 29486 16210 29538
rect 16210 29486 16212 29538
rect 16156 29484 16212 29486
rect 15596 29314 15652 29316
rect 15596 29262 15598 29314
rect 15598 29262 15650 29314
rect 15650 29262 15652 29314
rect 15596 29260 15652 29262
rect 15484 29148 15540 29204
rect 15708 28924 15764 28980
rect 15932 29036 15988 29092
rect 16268 29036 16324 29092
rect 16380 28924 16436 28980
rect 15932 28700 15988 28756
rect 14028 28588 14084 28644
rect 15148 28588 15204 28644
rect 13580 28476 13636 28532
rect 13468 27804 13524 27860
rect 14140 27186 14196 27188
rect 14140 27134 14142 27186
rect 14142 27134 14194 27186
rect 14194 27134 14196 27186
rect 14140 27132 14196 27134
rect 14364 26514 14420 26516
rect 14364 26462 14366 26514
rect 14366 26462 14418 26514
rect 14418 26462 14420 26514
rect 14364 26460 14420 26462
rect 14476 26572 14532 26628
rect 12460 24834 12516 24836
rect 12460 24782 12462 24834
rect 12462 24782 12514 24834
rect 12514 24782 12516 24834
rect 12460 24780 12516 24782
rect 11340 23100 11396 23156
rect 12684 23154 12740 23156
rect 12684 23102 12686 23154
rect 12686 23102 12738 23154
rect 12738 23102 12740 23154
rect 12684 23100 12740 23102
rect 14364 25506 14420 25508
rect 14364 25454 14366 25506
rect 14366 25454 14418 25506
rect 14418 25454 14420 25506
rect 14364 25452 14420 25454
rect 14476 24722 14532 24724
rect 14476 24670 14478 24722
rect 14478 24670 14530 24722
rect 14530 24670 14532 24722
rect 14476 24668 14532 24670
rect 13020 22204 13076 22260
rect 11340 21586 11396 21588
rect 11340 21534 11342 21586
rect 11342 21534 11394 21586
rect 11394 21534 11396 21586
rect 11340 21532 11396 21534
rect 13468 22370 13524 22372
rect 13468 22318 13470 22370
rect 13470 22318 13522 22370
rect 13522 22318 13524 22370
rect 13468 22316 13524 22318
rect 13580 21810 13636 21812
rect 13580 21758 13582 21810
rect 13582 21758 13634 21810
rect 13634 21758 13636 21810
rect 13580 21756 13636 21758
rect 11340 20636 11396 20692
rect 10220 19852 10276 19908
rect 9436 18396 9492 18452
rect 10892 19906 10948 19908
rect 10892 19854 10894 19906
rect 10894 19854 10946 19906
rect 10946 19854 10948 19906
rect 10892 19852 10948 19854
rect 11228 20188 11284 20244
rect 10220 18620 10276 18676
rect 10108 18562 10164 18564
rect 10108 18510 10110 18562
rect 10110 18510 10162 18562
rect 10162 18510 10164 18562
rect 10108 18508 10164 18510
rect 10556 18508 10612 18564
rect 10444 18396 10500 18452
rect 10444 17836 10500 17892
rect 9660 16994 9716 16996
rect 9660 16942 9662 16994
rect 9662 16942 9714 16994
rect 9714 16942 9716 16994
rect 9660 16940 9716 16942
rect 10668 18620 10724 18676
rect 11452 19852 11508 19908
rect 11452 19292 11508 19348
rect 11228 18620 11284 18676
rect 11004 18284 11060 18340
rect 11116 17442 11172 17444
rect 11116 17390 11118 17442
rect 11118 17390 11170 17442
rect 11170 17390 11172 17442
rect 11116 17388 11172 17390
rect 11004 15986 11060 15988
rect 11004 15934 11006 15986
rect 11006 15934 11058 15986
rect 11058 15934 11060 15986
rect 11004 15932 11060 15934
rect 11452 17724 11508 17780
rect 12012 17778 12068 17780
rect 12012 17726 12014 17778
rect 12014 17726 12066 17778
rect 12066 17726 12068 17778
rect 12012 17724 12068 17726
rect 11564 16828 11620 16884
rect 12908 16098 12964 16100
rect 12908 16046 12910 16098
rect 12910 16046 12962 16098
rect 12962 16046 12964 16098
rect 12908 16044 12964 16046
rect 11900 15932 11956 15988
rect 8540 13916 8596 13972
rect 7308 13356 7364 13412
rect 6972 13020 7028 13076
rect 5964 12684 6020 12740
rect 6636 12460 6692 12516
rect 5628 12178 5684 12180
rect 5628 12126 5630 12178
rect 5630 12126 5682 12178
rect 5682 12126 5684 12178
rect 5628 12124 5684 12126
rect 5516 11788 5572 11844
rect 6748 12124 6804 12180
rect 6076 11788 6132 11844
rect 6860 11788 6916 11844
rect 6748 11394 6804 11396
rect 6748 11342 6750 11394
rect 6750 11342 6802 11394
rect 6802 11342 6804 11394
rect 6748 11340 6804 11342
rect 8428 13356 8484 13412
rect 7420 12850 7476 12852
rect 7420 12798 7422 12850
rect 7422 12798 7474 12850
rect 7474 12798 7476 12850
rect 7420 12796 7476 12798
rect 10668 14252 10724 14308
rect 9996 13970 10052 13972
rect 9996 13918 9998 13970
rect 9998 13918 10050 13970
rect 10050 13918 10052 13970
rect 9996 13916 10052 13918
rect 8764 13020 8820 13076
rect 8652 12908 8708 12964
rect 8988 12908 9044 12964
rect 8876 12796 8932 12852
rect 7532 12236 7588 12292
rect 8316 12290 8372 12292
rect 8316 12238 8318 12290
rect 8318 12238 8370 12290
rect 8370 12238 8372 12290
rect 8316 12236 8372 12238
rect 9548 12908 9604 12964
rect 10220 13746 10276 13748
rect 10220 13694 10222 13746
rect 10222 13694 10274 13746
rect 10274 13694 10276 13746
rect 10220 13692 10276 13694
rect 9436 12348 9492 12404
rect 7308 11676 7364 11732
rect 5964 11282 6020 11284
rect 5964 11230 5966 11282
rect 5966 11230 6018 11282
rect 6018 11230 6020 11282
rect 5964 11228 6020 11230
rect 5852 11170 5908 11172
rect 5852 11118 5854 11170
rect 5854 11118 5906 11170
rect 5906 11118 5908 11170
rect 5852 11116 5908 11118
rect 7084 11004 7140 11060
rect 7644 11004 7700 11060
rect 6188 10780 6244 10836
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 7756 9884 7812 9940
rect 9548 12290 9604 12292
rect 9548 12238 9550 12290
rect 9550 12238 9602 12290
rect 9602 12238 9604 12290
rect 9548 12236 9604 12238
rect 9436 9884 9492 9940
rect 9884 12796 9940 12852
rect 9772 12402 9828 12404
rect 9772 12350 9774 12402
rect 9774 12350 9826 12402
rect 9826 12350 9828 12402
rect 9772 12348 9828 12350
rect 9660 12124 9716 12180
rect 10108 12460 10164 12516
rect 11452 12460 11508 12516
rect 11004 12348 11060 12404
rect 10668 12178 10724 12180
rect 10668 12126 10670 12178
rect 10670 12126 10722 12178
rect 10722 12126 10724 12178
rect 10668 12124 10724 12126
rect 9772 12012 9828 12068
rect 11004 12012 11060 12068
rect 12572 15986 12628 15988
rect 12572 15934 12574 15986
rect 12574 15934 12626 15986
rect 12626 15934 12628 15986
rect 12572 15932 12628 15934
rect 12460 15036 12516 15092
rect 12460 12850 12516 12852
rect 12460 12798 12462 12850
rect 12462 12798 12514 12850
rect 12514 12798 12516 12850
rect 12460 12796 12516 12798
rect 13244 12460 13300 12516
rect 12012 11116 12068 11172
rect 11676 10834 11732 10836
rect 11676 10782 11678 10834
rect 11678 10782 11730 10834
rect 11730 10782 11732 10834
rect 11676 10780 11732 10782
rect 12908 11116 12964 11172
rect 11788 10610 11844 10612
rect 11788 10558 11790 10610
rect 11790 10558 11842 10610
rect 11842 10558 11844 10610
rect 11788 10556 11844 10558
rect 5180 7980 5236 8036
rect 7084 7980 7140 8036
rect 10556 8034 10612 8036
rect 10556 7982 10558 8034
rect 10558 7982 10610 8034
rect 10610 7982 10612 8034
rect 10556 7980 10612 7982
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 10220 5906 10276 5908
rect 10220 5854 10222 5906
rect 10222 5854 10274 5906
rect 10274 5854 10276 5906
rect 10220 5852 10276 5854
rect 12012 10108 12068 10164
rect 11564 9714 11620 9716
rect 11564 9662 11566 9714
rect 11566 9662 11618 9714
rect 11618 9662 11620 9714
rect 11564 9660 11620 9662
rect 12124 9884 12180 9940
rect 12236 10556 12292 10612
rect 14028 20524 14084 20580
rect 13692 20188 13748 20244
rect 14028 17666 14084 17668
rect 14028 17614 14030 17666
rect 14030 17614 14082 17666
rect 14082 17614 14084 17666
rect 14028 17612 14084 17614
rect 13804 16098 13860 16100
rect 13804 16046 13806 16098
rect 13806 16046 13858 16098
rect 13858 16046 13860 16098
rect 13804 16044 13860 16046
rect 14476 22258 14532 22260
rect 14476 22206 14478 22258
rect 14478 22206 14530 22258
rect 14530 22206 14532 22258
rect 14476 22204 14532 22206
rect 14924 26236 14980 26292
rect 16044 28642 16100 28644
rect 16044 28590 16046 28642
rect 16046 28590 16098 28642
rect 16098 28590 16100 28642
rect 16044 28588 16100 28590
rect 17500 29372 17556 29428
rect 17388 28924 17444 28980
rect 17276 28754 17332 28756
rect 17276 28702 17278 28754
rect 17278 28702 17330 28754
rect 17330 28702 17332 28754
rect 17276 28700 17332 28702
rect 15260 27132 15316 27188
rect 16156 27186 16212 27188
rect 16156 27134 16158 27186
rect 16158 27134 16210 27186
rect 16210 27134 16212 27186
rect 16156 27132 16212 27134
rect 15596 26796 15652 26852
rect 15260 26460 15316 26516
rect 16044 26290 16100 26292
rect 16044 26238 16046 26290
rect 16046 26238 16098 26290
rect 16098 26238 16100 26290
rect 16044 26236 16100 26238
rect 16268 26236 16324 26292
rect 16156 26178 16212 26180
rect 16156 26126 16158 26178
rect 16158 26126 16210 26178
rect 16210 26126 16212 26178
rect 16156 26124 16212 26126
rect 15148 24668 15204 24724
rect 16380 25228 16436 25284
rect 15036 23324 15092 23380
rect 15148 22428 15204 22484
rect 15372 23324 15428 23380
rect 15932 22652 15988 22708
rect 17612 28588 17668 28644
rect 17276 26850 17332 26852
rect 17276 26798 17278 26850
rect 17278 26798 17330 26850
rect 17330 26798 17332 26850
rect 17276 26796 17332 26798
rect 17724 26908 17780 26964
rect 17836 27132 17892 27188
rect 17388 26290 17444 26292
rect 17388 26238 17390 26290
rect 17390 26238 17442 26290
rect 17442 26238 17444 26290
rect 17388 26236 17444 26238
rect 18060 28700 18116 28756
rect 18172 29372 18228 29428
rect 18060 27970 18116 27972
rect 18060 27918 18062 27970
rect 18062 27918 18114 27970
rect 18114 27918 18116 27970
rect 18060 27916 18116 27918
rect 17948 26796 18004 26852
rect 18060 26908 18116 26964
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 20300 29986 20356 29988
rect 20300 29934 20302 29986
rect 20302 29934 20354 29986
rect 20354 29934 20356 29986
rect 20300 29932 20356 29934
rect 18620 29484 18676 29540
rect 18396 28754 18452 28756
rect 18396 28702 18398 28754
rect 18398 28702 18450 28754
rect 18450 28702 18452 28754
rect 18396 28700 18452 28702
rect 18508 28588 18564 28644
rect 18284 26460 18340 26516
rect 18508 26796 18564 26852
rect 18060 26348 18116 26404
rect 18172 26290 18228 26292
rect 18172 26238 18174 26290
rect 18174 26238 18226 26290
rect 18226 26238 18228 26290
rect 18172 26236 18228 26238
rect 17164 25394 17220 25396
rect 17164 25342 17166 25394
rect 17166 25342 17218 25394
rect 17218 25342 17220 25394
rect 17164 25340 17220 25342
rect 15372 22316 15428 22372
rect 15708 22540 15764 22596
rect 15932 22482 15988 22484
rect 15932 22430 15934 22482
rect 15934 22430 15986 22482
rect 15986 22430 15988 22482
rect 15932 22428 15988 22430
rect 15036 20690 15092 20692
rect 15036 20638 15038 20690
rect 15038 20638 15090 20690
rect 15090 20638 15092 20690
rect 15036 20636 15092 20638
rect 14588 20018 14644 20020
rect 14588 19966 14590 20018
rect 14590 19966 14642 20018
rect 14642 19966 14644 20018
rect 14588 19964 14644 19966
rect 14252 18674 14308 18676
rect 14252 18622 14254 18674
rect 14254 18622 14306 18674
rect 14306 18622 14308 18674
rect 14252 18620 14308 18622
rect 14476 18562 14532 18564
rect 14476 18510 14478 18562
rect 14478 18510 14530 18562
rect 14530 18510 14532 18562
rect 14476 18508 14532 18510
rect 14364 18450 14420 18452
rect 14364 18398 14366 18450
rect 14366 18398 14418 18450
rect 14418 18398 14420 18450
rect 14364 18396 14420 18398
rect 14476 17948 14532 18004
rect 14476 17724 14532 17780
rect 18172 25394 18228 25396
rect 18172 25342 18174 25394
rect 18174 25342 18226 25394
rect 18226 25342 18228 25394
rect 18172 25340 18228 25342
rect 19292 29426 19348 29428
rect 19292 29374 19294 29426
rect 19294 29374 19346 29426
rect 19346 29374 19348 29426
rect 19292 29372 19348 29374
rect 19068 29260 19124 29316
rect 18844 28476 18900 28532
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 18844 26908 18900 26964
rect 18956 26290 19012 26292
rect 18956 26238 18958 26290
rect 18958 26238 19010 26290
rect 19010 26238 19012 26290
rect 18956 26236 19012 26238
rect 18732 26012 18788 26068
rect 18732 25228 18788 25284
rect 18956 23884 19012 23940
rect 17164 22540 17220 22596
rect 17276 22988 17332 23044
rect 17164 22370 17220 22372
rect 17164 22318 17166 22370
rect 17166 22318 17218 22370
rect 17218 22318 17220 22370
rect 17164 22316 17220 22318
rect 17052 22258 17108 22260
rect 17052 22206 17054 22258
rect 17054 22206 17106 22258
rect 17106 22206 17108 22258
rect 17052 22204 17108 22206
rect 17052 21756 17108 21812
rect 14812 18620 14868 18676
rect 15036 18508 15092 18564
rect 15260 18226 15316 18228
rect 15260 18174 15262 18226
rect 15262 18174 15314 18226
rect 15314 18174 15316 18226
rect 15260 18172 15316 18174
rect 15036 17836 15092 17892
rect 15708 18450 15764 18452
rect 15708 18398 15710 18450
rect 15710 18398 15762 18450
rect 15762 18398 15764 18450
rect 15708 18396 15764 18398
rect 15484 17612 15540 17668
rect 15708 15820 15764 15876
rect 13692 13916 13748 13972
rect 15484 14418 15540 14420
rect 15484 14366 15486 14418
rect 15486 14366 15538 14418
rect 15538 14366 15540 14418
rect 15484 14364 15540 14366
rect 14364 13746 14420 13748
rect 14364 13694 14366 13746
rect 14366 13694 14418 13746
rect 14418 13694 14420 13746
rect 14364 13692 14420 13694
rect 15036 13692 15092 13748
rect 14140 13580 14196 13636
rect 14924 13580 14980 13636
rect 15372 13468 15428 13524
rect 15596 13580 15652 13636
rect 15484 13020 15540 13076
rect 15820 14364 15876 14420
rect 16156 18172 16212 18228
rect 16828 17836 16884 17892
rect 16044 13468 16100 13524
rect 14028 12796 14084 12852
rect 13356 12348 13412 12404
rect 13244 10780 13300 10836
rect 13468 10556 13524 10612
rect 12908 10108 12964 10164
rect 12348 9714 12404 9716
rect 12348 9662 12350 9714
rect 12350 9662 12402 9714
rect 12402 9662 12404 9714
rect 12348 9660 12404 9662
rect 12572 9660 12628 9716
rect 12796 9660 12852 9716
rect 13916 11282 13972 11284
rect 13916 11230 13918 11282
rect 13918 11230 13970 11282
rect 13970 11230 13972 11282
rect 13916 11228 13972 11230
rect 14364 11452 14420 11508
rect 14140 11228 14196 11284
rect 13804 9884 13860 9940
rect 14028 9884 14084 9940
rect 14924 11506 14980 11508
rect 14924 11454 14926 11506
rect 14926 11454 14978 11506
rect 14978 11454 14980 11506
rect 14924 11452 14980 11454
rect 14588 10610 14644 10612
rect 14588 10558 14590 10610
rect 14590 10558 14642 10610
rect 14642 10558 14644 10610
rect 14588 10556 14644 10558
rect 15260 10834 15316 10836
rect 15260 10782 15262 10834
rect 15262 10782 15314 10834
rect 15314 10782 15316 10834
rect 15260 10780 15316 10782
rect 14924 10332 14980 10388
rect 13020 6748 13076 6804
rect 10556 5852 10612 5908
rect 13468 5906 13524 5908
rect 13468 5854 13470 5906
rect 13470 5854 13522 5906
rect 13522 5854 13524 5906
rect 13468 5852 13524 5854
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 15820 9772 15876 9828
rect 14588 8092 14644 8148
rect 13804 6748 13860 6804
rect 15484 6748 15540 6804
rect 16044 6748 16100 6804
rect 15260 5068 15316 5124
rect 12460 4338 12516 4340
rect 12460 4286 12462 4338
rect 12462 4286 12514 4338
rect 12514 4286 12516 4338
rect 12460 4284 12516 4286
rect 15932 5122 15988 5124
rect 15932 5070 15934 5122
rect 15934 5070 15986 5122
rect 15986 5070 15988 5122
rect 15932 5068 15988 5070
rect 17836 19346 17892 19348
rect 17836 19294 17838 19346
rect 17838 19294 17890 19346
rect 17890 19294 17892 19346
rect 17836 19292 17892 19294
rect 18844 22540 18900 22596
rect 20636 27244 20692 27300
rect 20188 27020 20244 27076
rect 20524 26962 20580 26964
rect 20524 26910 20526 26962
rect 20526 26910 20578 26962
rect 20578 26910 20580 26962
rect 20524 26908 20580 26910
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19852 26514 19908 26516
rect 19852 26462 19854 26514
rect 19854 26462 19906 26514
rect 19906 26462 19908 26514
rect 19852 26460 19908 26462
rect 19180 26348 19236 26404
rect 20188 26290 20244 26292
rect 20188 26238 20190 26290
rect 20190 26238 20242 26290
rect 20242 26238 20244 26290
rect 20188 26236 20244 26238
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 21420 30994 21476 30996
rect 21420 30942 21422 30994
rect 21422 30942 21474 30994
rect 21474 30942 21476 30994
rect 21420 30940 21476 30942
rect 28700 36652 28756 36708
rect 26012 34914 26068 34916
rect 26012 34862 26014 34914
rect 26014 34862 26066 34914
rect 26066 34862 26068 34914
rect 26012 34860 26068 34862
rect 24220 32508 24276 32564
rect 24668 32620 24724 32676
rect 24108 31666 24164 31668
rect 24108 31614 24110 31666
rect 24110 31614 24162 31666
rect 24162 31614 24164 31666
rect 24108 31612 24164 31614
rect 25228 32674 25284 32676
rect 25228 32622 25230 32674
rect 25230 32622 25282 32674
rect 25282 32622 25284 32674
rect 25228 32620 25284 32622
rect 25340 32562 25396 32564
rect 25340 32510 25342 32562
rect 25342 32510 25394 32562
rect 25394 32510 25396 32562
rect 25340 32508 25396 32510
rect 25452 32284 25508 32340
rect 23548 29260 23604 29316
rect 24780 31666 24836 31668
rect 24780 31614 24782 31666
rect 24782 31614 24834 31666
rect 24834 31614 24836 31666
rect 24780 31612 24836 31614
rect 23996 28924 24052 28980
rect 22876 28642 22932 28644
rect 22876 28590 22878 28642
rect 22878 28590 22930 28642
rect 22930 28590 22932 28642
rect 22876 28588 22932 28590
rect 21980 27132 22036 27188
rect 22540 27132 22596 27188
rect 21756 27020 21812 27076
rect 21084 23996 21140 24052
rect 21308 26962 21364 26964
rect 21308 26910 21310 26962
rect 21310 26910 21362 26962
rect 21362 26910 21364 26962
rect 21308 26908 21364 26910
rect 19292 23938 19348 23940
rect 19292 23886 19294 23938
rect 19294 23886 19346 23938
rect 19346 23886 19348 23938
rect 19292 23884 19348 23886
rect 19180 22764 19236 22820
rect 19404 22594 19460 22596
rect 19404 22542 19406 22594
rect 19406 22542 19458 22594
rect 19458 22542 19460 22594
rect 19404 22540 19460 22542
rect 18844 22204 18900 22260
rect 19068 21698 19124 21700
rect 19068 21646 19070 21698
rect 19070 21646 19122 21698
rect 19122 21646 19124 21698
rect 19068 21644 19124 21646
rect 17948 17948 18004 18004
rect 17500 17836 17556 17892
rect 17276 17612 17332 17668
rect 17276 17442 17332 17444
rect 17276 17390 17278 17442
rect 17278 17390 17330 17442
rect 17330 17390 17332 17442
rect 17276 17388 17332 17390
rect 17276 16828 17332 16884
rect 17612 15484 17668 15540
rect 18060 15148 18116 15204
rect 18396 16828 18452 16884
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20188 23436 20244 23492
rect 19852 23154 19908 23156
rect 19852 23102 19854 23154
rect 19854 23102 19906 23154
rect 19906 23102 19908 23154
rect 19852 23100 19908 23102
rect 20412 23324 20468 23380
rect 20748 23154 20804 23156
rect 20748 23102 20750 23154
rect 20750 23102 20802 23154
rect 20802 23102 20804 23154
rect 20748 23100 20804 23102
rect 19740 22764 19796 22820
rect 21084 22764 21140 22820
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 22204 26962 22260 26964
rect 22204 26910 22206 26962
rect 22206 26910 22258 26962
rect 22258 26910 22260 26962
rect 22204 26908 22260 26910
rect 22876 26124 22932 26180
rect 21532 25452 21588 25508
rect 22764 25340 22820 25396
rect 21532 23378 21588 23380
rect 21532 23326 21534 23378
rect 21534 23326 21586 23378
rect 21586 23326 21588 23378
rect 21532 23324 21588 23326
rect 21532 22092 21588 22148
rect 19068 19964 19124 20020
rect 19068 18562 19124 18564
rect 19068 18510 19070 18562
rect 19070 18510 19122 18562
rect 19122 18510 19124 18562
rect 19068 18508 19124 18510
rect 19740 20018 19796 20020
rect 19740 19966 19742 20018
rect 19742 19966 19794 20018
rect 19794 19966 19796 20018
rect 19740 19964 19796 19966
rect 20188 19292 20244 19348
rect 19292 18450 19348 18452
rect 19292 18398 19294 18450
rect 19294 18398 19346 18450
rect 19346 18398 19348 18450
rect 19292 18396 19348 18398
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 20188 18396 20244 18452
rect 20300 18172 20356 18228
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20748 18450 20804 18452
rect 20748 18398 20750 18450
rect 20750 18398 20802 18450
rect 20802 18398 20804 18450
rect 20748 18396 20804 18398
rect 20636 16828 20692 16884
rect 18956 16044 19012 16100
rect 19964 15874 20020 15876
rect 19964 15822 19966 15874
rect 19966 15822 20018 15874
rect 20018 15822 20020 15874
rect 19964 15820 20020 15822
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19516 15484 19572 15540
rect 17836 13074 17892 13076
rect 17836 13022 17838 13074
rect 17838 13022 17890 13074
rect 17890 13022 17892 13074
rect 17836 13020 17892 13022
rect 17276 10668 17332 10724
rect 18284 10498 18340 10500
rect 18284 10446 18286 10498
rect 18286 10446 18338 10498
rect 18338 10446 18340 10498
rect 18284 10444 18340 10446
rect 17836 9996 17892 10052
rect 17500 9826 17556 9828
rect 17500 9774 17502 9826
rect 17502 9774 17554 9826
rect 17554 9774 17556 9826
rect 17500 9772 17556 9774
rect 17836 9042 17892 9044
rect 17836 8990 17838 9042
rect 17838 8990 17890 9042
rect 17890 8990 17892 9042
rect 17836 8988 17892 8990
rect 17836 8034 17892 8036
rect 17836 7982 17838 8034
rect 17838 7982 17890 8034
rect 17890 7982 17892 8034
rect 17836 7980 17892 7982
rect 17388 6076 17444 6132
rect 18284 9212 18340 9268
rect 18732 9324 18788 9380
rect 18508 9042 18564 9044
rect 18508 8990 18510 9042
rect 18510 8990 18562 9042
rect 18562 8990 18564 9042
rect 18508 8988 18564 8990
rect 18396 8876 18452 8932
rect 18284 8146 18340 8148
rect 18284 8094 18286 8146
rect 18286 8094 18338 8146
rect 18338 8094 18340 8146
rect 18284 8092 18340 8094
rect 18956 8204 19012 8260
rect 18844 8092 18900 8148
rect 15708 4338 15764 4340
rect 15708 4286 15710 4338
rect 15710 4286 15762 4338
rect 15762 4286 15764 4338
rect 15708 4284 15764 4286
rect 19292 9548 19348 9604
rect 19852 15538 19908 15540
rect 19852 15486 19854 15538
rect 19854 15486 19906 15538
rect 19906 15486 19908 15538
rect 19852 15484 19908 15486
rect 19628 15036 19684 15092
rect 20076 15036 20132 15092
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 21868 15036 21924 15092
rect 20412 13580 20468 13636
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19628 11340 19684 11396
rect 20412 11116 20468 11172
rect 20524 14476 20580 14532
rect 21084 13020 21140 13076
rect 20748 12402 20804 12404
rect 20748 12350 20750 12402
rect 20750 12350 20802 12402
rect 20802 12350 20804 12402
rect 20748 12348 20804 12350
rect 22652 23378 22708 23380
rect 22652 23326 22654 23378
rect 22654 23326 22706 23378
rect 22706 23326 22708 23378
rect 22652 23324 22708 23326
rect 23100 26012 23156 26068
rect 22876 25228 22932 25284
rect 23436 24050 23492 24052
rect 23436 23998 23438 24050
rect 23438 23998 23490 24050
rect 23490 23998 23492 24050
rect 23436 23996 23492 23998
rect 23884 24050 23940 24052
rect 23884 23998 23886 24050
rect 23886 23998 23938 24050
rect 23938 23998 23940 24050
rect 23884 23996 23940 23998
rect 22876 23436 22932 23492
rect 23548 23324 23604 23380
rect 23884 23042 23940 23044
rect 23884 22990 23886 23042
rect 23886 22990 23938 23042
rect 23938 22990 23940 23042
rect 23884 22988 23940 22990
rect 24220 25506 24276 25508
rect 24220 25454 24222 25506
rect 24222 25454 24274 25506
rect 24274 25454 24276 25506
rect 24220 25452 24276 25454
rect 24892 30210 24948 30212
rect 24892 30158 24894 30210
rect 24894 30158 24946 30210
rect 24946 30158 24948 30210
rect 24892 30156 24948 30158
rect 25676 30156 25732 30212
rect 25340 29314 25396 29316
rect 25340 29262 25342 29314
rect 25342 29262 25394 29314
rect 25394 29262 25396 29314
rect 25340 29260 25396 29262
rect 25564 29260 25620 29316
rect 27356 35586 27412 35588
rect 27356 35534 27358 35586
rect 27358 35534 27410 35586
rect 27410 35534 27412 35586
rect 27356 35532 27412 35534
rect 29036 34972 29092 35028
rect 27468 33964 27524 34020
rect 27356 33068 27412 33124
rect 28364 34914 28420 34916
rect 28364 34862 28366 34914
rect 28366 34862 28418 34914
rect 28418 34862 28420 34914
rect 28364 34860 28420 34862
rect 29372 34914 29428 34916
rect 29372 34862 29374 34914
rect 29374 34862 29426 34914
rect 29426 34862 29428 34914
rect 29372 34860 29428 34862
rect 28140 32284 28196 32340
rect 26908 30156 26964 30212
rect 29372 33068 29428 33124
rect 29148 32284 29204 32340
rect 30940 39618 30996 39620
rect 30940 39566 30942 39618
rect 30942 39566 30994 39618
rect 30994 39566 30996 39618
rect 30940 39564 30996 39566
rect 36316 41970 36372 41972
rect 36316 41918 36318 41970
rect 36318 41918 36370 41970
rect 36370 41918 36372 41970
rect 36316 41916 36372 41918
rect 36092 41804 36148 41860
rect 37324 41858 37380 41860
rect 37324 41806 37326 41858
rect 37326 41806 37378 41858
rect 37378 41806 37380 41858
rect 37324 41804 37380 41806
rect 39900 41804 39956 41860
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 41132 41858 41188 41860
rect 41132 41806 41134 41858
rect 41134 41806 41186 41858
rect 41186 41806 41188 41858
rect 41132 41804 41188 41806
rect 31948 39564 32004 39620
rect 34188 39618 34244 39620
rect 34188 39566 34190 39618
rect 34190 39566 34242 39618
rect 34242 39566 34244 39618
rect 34188 39564 34244 39566
rect 31612 37266 31668 37268
rect 31612 37214 31614 37266
rect 31614 37214 31666 37266
rect 31666 37214 31668 37266
rect 31612 37212 31668 37214
rect 30828 36540 30884 36596
rect 32060 37266 32116 37268
rect 32060 37214 32062 37266
rect 32062 37214 32114 37266
rect 32114 37214 32116 37266
rect 32060 37212 32116 37214
rect 32284 36652 32340 36708
rect 33516 36652 33572 36708
rect 32396 36258 32452 36260
rect 32396 36206 32398 36258
rect 32398 36206 32450 36258
rect 32450 36206 32452 36258
rect 32396 36204 32452 36206
rect 31948 34860 32004 34916
rect 33852 36594 33908 36596
rect 33852 36542 33854 36594
rect 33854 36542 33906 36594
rect 33906 36542 33908 36594
rect 33852 36540 33908 36542
rect 34412 36876 34468 36932
rect 33852 36258 33908 36260
rect 33852 36206 33854 36258
rect 33854 36206 33906 36258
rect 33906 36206 33908 36258
rect 33852 36204 33908 36206
rect 34636 36204 34692 36260
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 38108 40348 38164 40404
rect 36988 37938 37044 37940
rect 36988 37886 36990 37938
rect 36990 37886 37042 37938
rect 37042 37886 37044 37938
rect 36988 37884 37044 37886
rect 35308 37826 35364 37828
rect 35308 37774 35310 37826
rect 35310 37774 35362 37826
rect 35362 37774 35364 37826
rect 35308 37772 35364 37774
rect 35308 37212 35364 37268
rect 37436 37772 37492 37828
rect 37324 37436 37380 37492
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35420 36652 35476 36708
rect 34972 36370 35028 36372
rect 34972 36318 34974 36370
rect 34974 36318 35026 36370
rect 35026 36318 35028 36370
rect 34972 36316 35028 36318
rect 34636 35532 34692 35588
rect 32284 33292 32340 33348
rect 33180 33346 33236 33348
rect 33180 33294 33182 33346
rect 33182 33294 33234 33346
rect 33234 33294 33236 33346
rect 33180 33292 33236 33294
rect 32284 32620 32340 32676
rect 32508 32674 32564 32676
rect 32508 32622 32510 32674
rect 32510 32622 32562 32674
rect 32562 32622 32564 32674
rect 32508 32620 32564 32622
rect 33516 32508 33572 32564
rect 33404 32172 33460 32228
rect 33292 31836 33348 31892
rect 33852 32172 33908 32228
rect 34076 33346 34132 33348
rect 34076 33294 34078 33346
rect 34078 33294 34130 33346
rect 34130 33294 34132 33346
rect 34076 33292 34132 33294
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35084 34914 35140 34916
rect 35084 34862 35086 34914
rect 35086 34862 35138 34914
rect 35138 34862 35140 34914
rect 35084 34860 35140 34862
rect 34300 32620 34356 32676
rect 26236 29932 26292 29988
rect 26012 29314 26068 29316
rect 26012 29262 26014 29314
rect 26014 29262 26066 29314
rect 26066 29262 26068 29314
rect 26012 29260 26068 29262
rect 26124 28642 26180 28644
rect 26124 28590 26126 28642
rect 26126 28590 26178 28642
rect 26178 28590 26180 28642
rect 26124 28588 26180 28590
rect 25452 27186 25508 27188
rect 25452 27134 25454 27186
rect 25454 27134 25506 27186
rect 25506 27134 25508 27186
rect 25452 27132 25508 27134
rect 25900 27132 25956 27188
rect 24892 25506 24948 25508
rect 24892 25454 24894 25506
rect 24894 25454 24946 25506
rect 24946 25454 24948 25506
rect 24892 25452 24948 25454
rect 24444 25394 24500 25396
rect 24444 25342 24446 25394
rect 24446 25342 24498 25394
rect 24498 25342 24500 25394
rect 24444 25340 24500 25342
rect 24332 23996 24388 24052
rect 24892 23996 24948 24052
rect 24444 23154 24500 23156
rect 24444 23102 24446 23154
rect 24446 23102 24498 23154
rect 24498 23102 24500 23154
rect 24444 23100 24500 23102
rect 26012 23436 26068 23492
rect 25676 23100 25732 23156
rect 25228 21756 25284 21812
rect 22652 18172 22708 18228
rect 23212 18562 23268 18564
rect 23212 18510 23214 18562
rect 23214 18510 23266 18562
rect 23266 18510 23268 18562
rect 23212 18508 23268 18510
rect 23436 18562 23492 18564
rect 23436 18510 23438 18562
rect 23438 18510 23490 18562
rect 23490 18510 23492 18562
rect 23436 18508 23492 18510
rect 22876 17948 22932 18004
rect 22540 15036 22596 15092
rect 22876 17612 22932 17668
rect 21868 13074 21924 13076
rect 21868 13022 21870 13074
rect 21870 13022 21922 13074
rect 21922 13022 21924 13074
rect 21868 13020 21924 13022
rect 22652 12572 22708 12628
rect 22204 12402 22260 12404
rect 22204 12350 22206 12402
rect 22206 12350 22258 12402
rect 22258 12350 22260 12402
rect 22204 12348 22260 12350
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 21644 12124 21700 12180
rect 21308 11954 21364 11956
rect 21308 11902 21310 11954
rect 21310 11902 21362 11954
rect 21362 11902 21364 11954
rect 21308 11900 21364 11902
rect 21756 11394 21812 11396
rect 21756 11342 21758 11394
rect 21758 11342 21810 11394
rect 21810 11342 21812 11394
rect 21756 11340 21812 11342
rect 22428 12178 22484 12180
rect 22428 12126 22430 12178
rect 22430 12126 22482 12178
rect 22482 12126 22484 12178
rect 22428 12124 22484 12126
rect 22092 11900 22148 11956
rect 20524 10668 20580 10724
rect 19628 10444 19684 10500
rect 19628 9996 19684 10052
rect 20412 10050 20468 10052
rect 20412 9998 20414 10050
rect 20414 9998 20466 10050
rect 20466 9998 20468 10050
rect 20412 9996 20468 9998
rect 19628 9324 19684 9380
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19516 9212 19572 9268
rect 20076 9212 20132 9268
rect 20300 9602 20356 9604
rect 20300 9550 20302 9602
rect 20302 9550 20354 9602
rect 20354 9550 20356 9602
rect 20300 9548 20356 9550
rect 19628 8876 19684 8932
rect 23548 18450 23604 18452
rect 23548 18398 23550 18450
rect 23550 18398 23602 18450
rect 23602 18398 23604 18450
rect 23548 18396 23604 18398
rect 24780 19292 24836 19348
rect 24332 19122 24388 19124
rect 24332 19070 24334 19122
rect 24334 19070 24386 19122
rect 24386 19070 24388 19122
rect 24332 19068 24388 19070
rect 24444 18508 24500 18564
rect 23884 18172 23940 18228
rect 24108 18450 24164 18452
rect 24108 18398 24110 18450
rect 24110 18398 24162 18450
rect 24162 18398 24164 18450
rect 24108 18396 24164 18398
rect 23436 17666 23492 17668
rect 23436 17614 23438 17666
rect 23438 17614 23490 17666
rect 23490 17614 23492 17666
rect 23436 17612 23492 17614
rect 23100 16268 23156 16324
rect 23436 16322 23492 16324
rect 23436 16270 23438 16322
rect 23438 16270 23490 16322
rect 23490 16270 23492 16322
rect 23436 16268 23492 16270
rect 23996 16268 24052 16324
rect 23212 15426 23268 15428
rect 23212 15374 23214 15426
rect 23214 15374 23266 15426
rect 23266 15374 23268 15426
rect 23212 15372 23268 15374
rect 25564 22428 25620 22484
rect 25228 21308 25284 21364
rect 25228 18956 25284 19012
rect 25228 18284 25284 18340
rect 25004 15932 25060 15988
rect 24220 15596 24276 15652
rect 24220 15314 24276 15316
rect 24220 15262 24222 15314
rect 24222 15262 24274 15314
rect 24274 15262 24276 15314
rect 24220 15260 24276 15262
rect 23212 14588 23268 14644
rect 22988 14530 23044 14532
rect 22988 14478 22990 14530
rect 22990 14478 23042 14530
rect 23042 14478 23044 14530
rect 22988 14476 23044 14478
rect 22988 12684 23044 12740
rect 23100 12348 23156 12404
rect 23212 12684 23268 12740
rect 23212 11452 23268 11508
rect 23436 12572 23492 12628
rect 22652 11394 22708 11396
rect 22652 11342 22654 11394
rect 22654 11342 22706 11394
rect 22706 11342 22708 11394
rect 22652 11340 22708 11342
rect 24444 14588 24500 14644
rect 24668 14700 24724 14756
rect 25788 21810 25844 21812
rect 25788 21758 25790 21810
rect 25790 21758 25842 21810
rect 25842 21758 25844 21810
rect 25788 21756 25844 21758
rect 25900 21308 25956 21364
rect 25452 19122 25508 19124
rect 25452 19070 25454 19122
rect 25454 19070 25506 19122
rect 25506 19070 25508 19122
rect 25452 19068 25508 19070
rect 25340 15820 25396 15876
rect 25788 15596 25844 15652
rect 25340 15538 25396 15540
rect 25340 15486 25342 15538
rect 25342 15486 25394 15538
rect 25394 15486 25396 15538
rect 25340 15484 25396 15486
rect 25004 15260 25060 15316
rect 25452 14754 25508 14756
rect 25452 14702 25454 14754
rect 25454 14702 25506 14754
rect 25506 14702 25508 14754
rect 25452 14700 25508 14702
rect 25564 14642 25620 14644
rect 25564 14590 25566 14642
rect 25566 14590 25618 14642
rect 25618 14590 25620 14642
rect 25564 14588 25620 14590
rect 24556 13804 24612 13860
rect 23772 12572 23828 12628
rect 23884 12348 23940 12404
rect 24444 12738 24500 12740
rect 24444 12686 24446 12738
rect 24446 12686 24498 12738
rect 24498 12686 24500 12738
rect 24444 12684 24500 12686
rect 24556 12402 24612 12404
rect 24556 12350 24558 12402
rect 24558 12350 24610 12402
rect 24610 12350 24612 12402
rect 24556 12348 24612 12350
rect 24108 12290 24164 12292
rect 24108 12238 24110 12290
rect 24110 12238 24162 12290
rect 24162 12238 24164 12290
rect 24108 12236 24164 12238
rect 24668 12290 24724 12292
rect 24668 12238 24670 12290
rect 24670 12238 24722 12290
rect 24722 12238 24724 12290
rect 24668 12236 24724 12238
rect 23996 12178 24052 12180
rect 23996 12126 23998 12178
rect 23998 12126 24050 12178
rect 24050 12126 24052 12178
rect 23996 12124 24052 12126
rect 25452 12236 25508 12292
rect 26684 29260 26740 29316
rect 26348 27356 26404 27412
rect 26348 23154 26404 23156
rect 26348 23102 26350 23154
rect 26350 23102 26402 23154
rect 26402 23102 26404 23154
rect 26348 23100 26404 23102
rect 26236 22482 26292 22484
rect 26236 22430 26238 22482
rect 26238 22430 26290 22482
rect 26290 22430 26292 22482
rect 26236 22428 26292 22430
rect 26236 21756 26292 21812
rect 26012 17500 26068 17556
rect 26124 17724 26180 17780
rect 24668 11394 24724 11396
rect 24668 11342 24670 11394
rect 24670 11342 24722 11394
rect 24722 11342 24724 11394
rect 24668 11340 24724 11342
rect 25340 11340 25396 11396
rect 24220 11282 24276 11284
rect 24220 11230 24222 11282
rect 24222 11230 24274 11282
rect 24274 11230 24276 11282
rect 24220 11228 24276 11230
rect 19180 8092 19236 8148
rect 19068 6076 19124 6132
rect 18620 5740 18676 5796
rect 17388 4284 17444 4340
rect 19852 8258 19908 8260
rect 19852 8206 19854 8258
rect 19854 8206 19906 8258
rect 19906 8206 19908 8258
rect 19852 8204 19908 8206
rect 20412 8316 20468 8372
rect 21420 8370 21476 8372
rect 21420 8318 21422 8370
rect 21422 8318 21474 8370
rect 21474 8318 21476 8370
rect 21420 8316 21476 8318
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 23436 7980 23492 8036
rect 23884 8034 23940 8036
rect 23884 7982 23886 8034
rect 23886 7982 23938 8034
rect 23938 7982 23940 8034
rect 23884 7980 23940 7982
rect 24556 7644 24612 7700
rect 21868 6748 21924 6804
rect 22988 6748 23044 6804
rect 20076 6412 20132 6468
rect 21756 6412 21812 6468
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 20748 6130 20804 6132
rect 20748 6078 20750 6130
rect 20750 6078 20802 6130
rect 20802 6078 20804 6130
rect 20748 6076 20804 6078
rect 20300 5794 20356 5796
rect 20300 5742 20302 5794
rect 20302 5742 20354 5794
rect 20354 5742 20356 5794
rect 20300 5740 20356 5742
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 28252 28476 28308 28532
rect 27132 27020 27188 27076
rect 26796 26124 26852 26180
rect 28252 27020 28308 27076
rect 28588 29596 28644 29652
rect 29372 29932 29428 29988
rect 28812 29314 28868 29316
rect 28812 29262 28814 29314
rect 28814 29262 28866 29314
rect 28866 29262 28868 29314
rect 28812 29260 28868 29262
rect 29372 29260 29428 29316
rect 29932 29932 29988 29988
rect 28588 28812 28644 28868
rect 29372 28812 29428 28868
rect 28364 26908 28420 26964
rect 31052 28754 31108 28756
rect 31052 28702 31054 28754
rect 31054 28702 31106 28754
rect 31106 28702 31108 28754
rect 31052 28700 31108 28702
rect 30268 28642 30324 28644
rect 30268 28590 30270 28642
rect 30270 28590 30322 28642
rect 30322 28590 30324 28642
rect 30268 28588 30324 28590
rect 29484 26908 29540 26964
rect 27804 25394 27860 25396
rect 27804 25342 27806 25394
rect 27806 25342 27858 25394
rect 27858 25342 27860 25394
rect 27804 25340 27860 25342
rect 27468 25282 27524 25284
rect 27468 25230 27470 25282
rect 27470 25230 27522 25282
rect 27522 25230 27524 25282
rect 27468 25228 27524 25230
rect 29260 25394 29316 25396
rect 29260 25342 29262 25394
rect 29262 25342 29314 25394
rect 29314 25342 29316 25394
rect 29260 25340 29316 25342
rect 27692 24556 27748 24612
rect 28476 24610 28532 24612
rect 28476 24558 28478 24610
rect 28478 24558 28530 24610
rect 28530 24558 28532 24610
rect 28476 24556 28532 24558
rect 28476 23660 28532 23716
rect 28924 23324 28980 23380
rect 29820 26908 29876 26964
rect 29708 25228 29764 25284
rect 29820 25452 29876 25508
rect 31388 28588 31444 28644
rect 33516 31554 33572 31556
rect 33516 31502 33518 31554
rect 33518 31502 33570 31554
rect 33570 31502 33572 31554
rect 33516 31500 33572 31502
rect 32620 29932 32676 29988
rect 33068 30380 33124 30436
rect 32508 28476 32564 28532
rect 33180 30268 33236 30324
rect 30268 26962 30324 26964
rect 30268 26910 30270 26962
rect 30270 26910 30322 26962
rect 30322 26910 30324 26962
rect 30268 26908 30324 26910
rect 30044 26178 30100 26180
rect 30044 26126 30046 26178
rect 30046 26126 30098 26178
rect 30098 26126 30100 26178
rect 30044 26124 30100 26126
rect 29484 23714 29540 23716
rect 29484 23662 29486 23714
rect 29486 23662 29538 23714
rect 29538 23662 29540 23714
rect 29484 23660 29540 23662
rect 29148 23266 29204 23268
rect 29148 23214 29150 23266
rect 29150 23214 29202 23266
rect 29202 23214 29204 23266
rect 29148 23212 29204 23214
rect 26572 21756 26628 21812
rect 28924 21698 28980 21700
rect 28924 21646 28926 21698
rect 28926 21646 28978 21698
rect 28978 21646 28980 21698
rect 28924 21644 28980 21646
rect 29596 21698 29652 21700
rect 29596 21646 29598 21698
rect 29598 21646 29650 21698
rect 29650 21646 29652 21698
rect 29596 21644 29652 21646
rect 30156 25282 30212 25284
rect 30156 25230 30158 25282
rect 30158 25230 30210 25282
rect 30210 25230 30212 25282
rect 30156 25228 30212 25230
rect 32732 24668 32788 24724
rect 31724 24556 31780 24612
rect 30268 23884 30324 23940
rect 31052 23938 31108 23940
rect 31052 23886 31054 23938
rect 31054 23886 31106 23938
rect 31106 23886 31108 23938
rect 31052 23884 31108 23886
rect 29932 23324 29988 23380
rect 33180 29202 33236 29204
rect 33180 29150 33182 29202
rect 33182 29150 33234 29202
rect 33234 29150 33236 29202
rect 33180 29148 33236 29150
rect 33740 29148 33796 29204
rect 33852 28700 33908 28756
rect 34412 31724 34468 31780
rect 34188 30268 34244 30324
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 36988 36988 37044 37044
rect 39676 39340 39732 39396
rect 40460 40402 40516 40404
rect 40460 40350 40462 40402
rect 40462 40350 40514 40402
rect 40514 40350 40516 40402
rect 40460 40348 40516 40350
rect 39452 38050 39508 38052
rect 39452 37998 39454 38050
rect 39454 37998 39506 38050
rect 39506 37998 39508 38050
rect 39452 37996 39508 37998
rect 40348 40236 40404 40292
rect 38556 36876 38612 36932
rect 36652 36316 36708 36372
rect 37100 36258 37156 36260
rect 37100 36206 37102 36258
rect 37102 36206 37154 36258
rect 37154 36206 37156 36258
rect 37100 36204 37156 36206
rect 36540 35698 36596 35700
rect 36540 35646 36542 35698
rect 36542 35646 36594 35698
rect 36594 35646 36596 35698
rect 36540 35644 36596 35646
rect 35532 32508 35588 32564
rect 34748 32396 34804 32452
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 37324 35532 37380 35588
rect 37436 35980 37492 36036
rect 39228 37266 39284 37268
rect 39228 37214 39230 37266
rect 39230 37214 39282 37266
rect 39282 37214 39284 37266
rect 39228 37212 39284 37214
rect 39116 36258 39172 36260
rect 39116 36206 39118 36258
rect 39118 36206 39170 36258
rect 39170 36206 39172 36258
rect 39116 36204 39172 36206
rect 38780 35980 38836 36036
rect 37548 35644 37604 35700
rect 36428 32562 36484 32564
rect 36428 32510 36430 32562
rect 36430 32510 36482 32562
rect 36482 32510 36484 32562
rect 36428 32508 36484 32510
rect 35980 32450 36036 32452
rect 35980 32398 35982 32450
rect 35982 32398 36034 32450
rect 36034 32398 36036 32450
rect 35980 32396 36036 32398
rect 34972 31554 35028 31556
rect 34972 31502 34974 31554
rect 34974 31502 35026 31554
rect 35026 31502 35028 31554
rect 34972 31500 35028 31502
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34636 30380 34692 30436
rect 34524 29708 34580 29764
rect 35756 29708 35812 29764
rect 34188 29148 34244 29204
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35084 28812 35140 28868
rect 33964 25564 34020 25620
rect 33852 25452 33908 25508
rect 33180 24722 33236 24724
rect 33180 24670 33182 24722
rect 33182 24670 33234 24722
rect 33234 24670 33236 24722
rect 33180 24668 33236 24670
rect 33292 23436 33348 23492
rect 33068 23266 33124 23268
rect 33068 23214 33070 23266
rect 33070 23214 33122 23266
rect 33122 23214 33124 23266
rect 33068 23212 33124 23214
rect 33180 23100 33236 23156
rect 33516 24610 33572 24612
rect 33516 24558 33518 24610
rect 33518 24558 33570 24610
rect 33570 24558 33572 24610
rect 33516 24556 33572 24558
rect 34748 25676 34804 25732
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35308 26850 35364 26852
rect 35308 26798 35310 26850
rect 35310 26798 35362 26850
rect 35362 26798 35364 26850
rect 35308 26796 35364 26798
rect 36540 31554 36596 31556
rect 36540 31502 36542 31554
rect 36542 31502 36594 31554
rect 36594 31502 36596 31554
rect 36540 31500 36596 31502
rect 36652 29538 36708 29540
rect 36652 29486 36654 29538
rect 36654 29486 36706 29538
rect 36706 29486 36708 29538
rect 36652 29484 36708 29486
rect 35980 28812 36036 28868
rect 36428 27186 36484 27188
rect 36428 27134 36430 27186
rect 36430 27134 36482 27186
rect 36482 27134 36484 27186
rect 36428 27132 36484 27134
rect 37436 33516 37492 33572
rect 36876 32508 36932 32564
rect 37660 32396 37716 32452
rect 39116 33516 39172 33572
rect 36988 31554 37044 31556
rect 36988 31502 36990 31554
rect 36990 31502 37042 31554
rect 37042 31502 37044 31554
rect 36988 31500 37044 31502
rect 37100 30210 37156 30212
rect 37100 30158 37102 30210
rect 37102 30158 37154 30210
rect 37154 30158 37156 30210
rect 37100 30156 37156 30158
rect 37660 29708 37716 29764
rect 37548 29650 37604 29652
rect 37548 29598 37550 29650
rect 37550 29598 37602 29650
rect 37602 29598 37604 29650
rect 37548 29596 37604 29598
rect 37212 29484 37268 29540
rect 36764 27132 36820 27188
rect 37100 27132 37156 27188
rect 36876 26796 36932 26852
rect 35868 26124 35924 26180
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35420 25676 35476 25732
rect 35084 25452 35140 25508
rect 35196 25340 35252 25396
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 34300 24050 34356 24052
rect 34300 23998 34302 24050
rect 34302 23998 34354 24050
rect 34354 23998 34356 24050
rect 34300 23996 34356 23998
rect 35532 24050 35588 24052
rect 35532 23998 35534 24050
rect 35534 23998 35586 24050
rect 35586 23998 35588 24050
rect 35532 23996 35588 23998
rect 30156 21586 30212 21588
rect 30156 21534 30158 21586
rect 30158 21534 30210 21586
rect 30210 21534 30212 21586
rect 30156 21532 30212 21534
rect 28028 19964 28084 20020
rect 29484 20018 29540 20020
rect 29484 19966 29486 20018
rect 29486 19966 29538 20018
rect 29538 19966 29540 20018
rect 29484 19964 29540 19966
rect 30604 21644 30660 21700
rect 30492 20188 30548 20244
rect 31276 20188 31332 20244
rect 28028 19346 28084 19348
rect 28028 19294 28030 19346
rect 28030 19294 28082 19346
rect 28082 19294 28084 19346
rect 28028 19292 28084 19294
rect 27580 18508 27636 18564
rect 29820 19010 29876 19012
rect 29820 18958 29822 19010
rect 29822 18958 29874 19010
rect 29874 18958 29876 19010
rect 29820 18956 29876 18958
rect 29596 16828 29652 16884
rect 28700 15820 28756 15876
rect 29260 14588 29316 14644
rect 27244 13858 27300 13860
rect 27244 13806 27246 13858
rect 27246 13806 27298 13858
rect 27298 13806 27300 13858
rect 27244 13804 27300 13806
rect 26572 13746 26628 13748
rect 26572 13694 26574 13746
rect 26574 13694 26626 13746
rect 26626 13694 26628 13746
rect 26572 13692 26628 13694
rect 27356 11282 27412 11284
rect 27356 11230 27358 11282
rect 27358 11230 27410 11282
rect 27410 11230 27412 11282
rect 27356 11228 27412 11230
rect 28588 10780 28644 10836
rect 26460 9548 26516 9604
rect 25116 8316 25172 8372
rect 25676 7980 25732 8036
rect 25340 7698 25396 7700
rect 25340 7646 25342 7698
rect 25342 7646 25394 7698
rect 25394 7646 25396 7698
rect 25340 7644 25396 7646
rect 24556 6748 24612 6804
rect 27804 7644 27860 7700
rect 27468 6636 27524 6692
rect 25676 5794 25732 5796
rect 25676 5742 25678 5794
rect 25678 5742 25730 5794
rect 25730 5742 25732 5794
rect 25676 5740 25732 5742
rect 26796 5794 26852 5796
rect 26796 5742 26798 5794
rect 26798 5742 26850 5794
rect 26850 5742 26852 5794
rect 26796 5740 26852 5742
rect 27692 5794 27748 5796
rect 27692 5742 27694 5794
rect 27694 5742 27746 5794
rect 27746 5742 27748 5794
rect 27692 5740 27748 5742
rect 30268 18956 30324 19012
rect 30604 18732 30660 18788
rect 30492 18172 30548 18228
rect 30492 17106 30548 17108
rect 30492 17054 30494 17106
rect 30494 17054 30546 17106
rect 30546 17054 30548 17106
rect 30492 17052 30548 17054
rect 30044 14588 30100 14644
rect 30044 13692 30100 13748
rect 30044 10780 30100 10836
rect 30156 9996 30212 10052
rect 29932 9826 29988 9828
rect 29932 9774 29934 9826
rect 29934 9774 29986 9826
rect 29986 9774 29988 9826
rect 29932 9772 29988 9774
rect 30604 9826 30660 9828
rect 30604 9774 30606 9826
rect 30606 9774 30658 9826
rect 30658 9774 30660 9826
rect 30604 9772 30660 9774
rect 30492 8988 30548 9044
rect 30604 9548 30660 9604
rect 28364 7644 28420 7700
rect 29820 6690 29876 6692
rect 29820 6638 29822 6690
rect 29822 6638 29874 6690
rect 29874 6638 29876 6690
rect 29820 6636 29876 6638
rect 28700 6018 28756 6020
rect 28700 5966 28702 6018
rect 28702 5966 28754 6018
rect 28754 5966 28756 6018
rect 28700 5964 28756 5966
rect 33852 23100 33908 23156
rect 34972 23154 35028 23156
rect 34972 23102 34974 23154
rect 34974 23102 35026 23154
rect 35026 23102 35028 23154
rect 34972 23100 35028 23102
rect 39004 29932 39060 29988
rect 38892 29650 38948 29652
rect 38892 29598 38894 29650
rect 38894 29598 38946 29650
rect 38946 29598 38948 29650
rect 38892 29596 38948 29598
rect 39564 37266 39620 37268
rect 39564 37214 39566 37266
rect 39566 37214 39618 37266
rect 39618 37214 39620 37266
rect 39564 37212 39620 37214
rect 39452 36594 39508 36596
rect 39452 36542 39454 36594
rect 39454 36542 39506 36594
rect 39506 36542 39508 36594
rect 39452 36540 39508 36542
rect 39340 36482 39396 36484
rect 39340 36430 39342 36482
rect 39342 36430 39394 36482
rect 39394 36430 39396 36482
rect 39340 36428 39396 36430
rect 39564 35644 39620 35700
rect 39228 32620 39284 32676
rect 39340 31778 39396 31780
rect 39340 31726 39342 31778
rect 39342 31726 39394 31778
rect 39394 31726 39396 31778
rect 39340 31724 39396 31726
rect 38668 29538 38724 29540
rect 38668 29486 38670 29538
rect 38670 29486 38722 29538
rect 38722 29486 38724 29538
rect 38668 29484 38724 29486
rect 37548 29202 37604 29204
rect 37548 29150 37550 29202
rect 37550 29150 37602 29202
rect 37602 29150 37604 29202
rect 37548 29148 37604 29150
rect 37660 26908 37716 26964
rect 37212 26514 37268 26516
rect 37212 26462 37214 26514
rect 37214 26462 37266 26514
rect 37266 26462 37268 26514
rect 37212 26460 37268 26462
rect 38780 26908 38836 26964
rect 38220 26460 38276 26516
rect 36876 26236 36932 26292
rect 37436 26290 37492 26292
rect 37436 26238 37438 26290
rect 37438 26238 37490 26290
rect 37490 26238 37492 26290
rect 37436 26236 37492 26238
rect 37324 26178 37380 26180
rect 37324 26126 37326 26178
rect 37326 26126 37378 26178
rect 37378 26126 37380 26178
rect 37324 26124 37380 26126
rect 37212 25618 37268 25620
rect 37212 25566 37214 25618
rect 37214 25566 37266 25618
rect 37266 25566 37268 25618
rect 37212 25564 37268 25566
rect 35868 24050 35924 24052
rect 35868 23998 35870 24050
rect 35870 23998 35922 24050
rect 35922 23998 35924 24050
rect 35868 23996 35924 23998
rect 36764 25340 36820 25396
rect 38220 25340 38276 25396
rect 36764 23436 36820 23492
rect 39452 26962 39508 26964
rect 39452 26910 39454 26962
rect 39454 26910 39506 26962
rect 39506 26910 39508 26962
rect 39452 26908 39508 26910
rect 39900 37938 39956 37940
rect 39900 37886 39902 37938
rect 39902 37886 39954 37938
rect 39954 37886 39956 37938
rect 39900 37884 39956 37886
rect 39788 37826 39844 37828
rect 39788 37774 39790 37826
rect 39790 37774 39842 37826
rect 39842 37774 39844 37826
rect 39788 37772 39844 37774
rect 39788 37490 39844 37492
rect 39788 37438 39790 37490
rect 39790 37438 39842 37490
rect 39842 37438 39844 37490
rect 39788 37436 39844 37438
rect 41020 40402 41076 40404
rect 41020 40350 41022 40402
rect 41022 40350 41074 40402
rect 41074 40350 41076 40402
rect 41020 40348 41076 40350
rect 41804 40290 41860 40292
rect 41804 40238 41806 40290
rect 41806 40238 41858 40290
rect 41858 40238 41860 40290
rect 41804 40236 41860 40238
rect 42700 40236 42756 40292
rect 43932 40290 43988 40292
rect 43932 40238 43934 40290
rect 43934 40238 43986 40290
rect 43986 40238 43988 40290
rect 43932 40236 43988 40238
rect 41132 39394 41188 39396
rect 41132 39342 41134 39394
rect 41134 39342 41186 39394
rect 41186 39342 41188 39394
rect 41132 39340 41188 39342
rect 39900 36876 39956 36932
rect 40012 36258 40068 36260
rect 40012 36206 40014 36258
rect 40014 36206 40066 36258
rect 40066 36206 40068 36258
rect 40012 36204 40068 36206
rect 41916 37772 41972 37828
rect 42588 37436 42644 37492
rect 40236 36876 40292 36932
rect 40124 35980 40180 36036
rect 40348 36428 40404 36484
rect 40572 36258 40628 36260
rect 40572 36206 40574 36258
rect 40574 36206 40626 36258
rect 40626 36206 40628 36258
rect 40572 36204 40628 36206
rect 40908 35980 40964 36036
rect 40236 32620 40292 32676
rect 40460 31836 40516 31892
rect 40348 30210 40404 30212
rect 40348 30158 40350 30210
rect 40350 30158 40402 30210
rect 40402 30158 40404 30210
rect 40348 30156 40404 30158
rect 44044 36428 44100 36484
rect 40908 33740 40964 33796
rect 41580 33740 41636 33796
rect 44044 33740 44100 33796
rect 41132 31836 41188 31892
rect 40796 29708 40852 29764
rect 41468 29932 41524 29988
rect 40348 29650 40404 29652
rect 40348 29598 40350 29650
rect 40350 29598 40402 29650
rect 40402 29598 40404 29650
rect 40348 29596 40404 29598
rect 41132 29596 41188 29652
rect 40460 29260 40516 29316
rect 40012 28754 40068 28756
rect 40012 28702 40014 28754
rect 40014 28702 40066 28754
rect 40066 28702 40068 28754
rect 40012 28700 40068 28702
rect 40460 28588 40516 28644
rect 41132 28642 41188 28644
rect 41132 28590 41134 28642
rect 41134 28590 41186 28642
rect 41186 28590 41188 28642
rect 41132 28588 41188 28590
rect 42700 30098 42756 30100
rect 42700 30046 42702 30098
rect 42702 30046 42754 30098
rect 42754 30046 42756 30098
rect 42700 30044 42756 30046
rect 44044 30044 44100 30100
rect 42588 29986 42644 29988
rect 42588 29934 42590 29986
rect 42590 29934 42642 29986
rect 42642 29934 42644 29986
rect 42588 29932 42644 29934
rect 41580 28700 41636 28756
rect 39900 27244 39956 27300
rect 40236 27020 40292 27076
rect 40124 26908 40180 26964
rect 39900 25618 39956 25620
rect 39900 25566 39902 25618
rect 39902 25566 39954 25618
rect 39954 25566 39956 25618
rect 39900 25564 39956 25566
rect 39676 25228 39732 25284
rect 39116 23996 39172 24052
rect 40796 27074 40852 27076
rect 40796 27022 40798 27074
rect 40798 27022 40850 27074
rect 40850 27022 40852 27074
rect 40796 27020 40852 27022
rect 40460 25506 40516 25508
rect 40460 25454 40462 25506
rect 40462 25454 40514 25506
rect 40514 25454 40516 25506
rect 40460 25452 40516 25454
rect 41132 25564 41188 25620
rect 40684 25394 40740 25396
rect 40684 25342 40686 25394
rect 40686 25342 40738 25394
rect 40738 25342 40740 25394
rect 40684 25340 40740 25342
rect 40124 23996 40180 24052
rect 40348 23548 40404 23604
rect 40684 23714 40740 23716
rect 40684 23662 40686 23714
rect 40686 23662 40738 23714
rect 40738 23662 40740 23714
rect 40684 23660 40740 23662
rect 38444 23100 38500 23156
rect 39452 23154 39508 23156
rect 39452 23102 39454 23154
rect 39454 23102 39506 23154
rect 39506 23102 39508 23154
rect 39452 23100 39508 23102
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35980 21532 36036 21588
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 31724 19234 31780 19236
rect 31724 19182 31726 19234
rect 31726 19182 31778 19234
rect 31778 19182 31780 19234
rect 31724 19180 31780 19182
rect 31612 18732 31668 18788
rect 31052 17388 31108 17444
rect 30940 17106 30996 17108
rect 30940 17054 30942 17106
rect 30942 17054 30994 17106
rect 30994 17054 30996 17106
rect 30940 17052 30996 17054
rect 31612 16882 31668 16884
rect 31612 16830 31614 16882
rect 31614 16830 31666 16882
rect 31666 16830 31668 16882
rect 31612 16828 31668 16830
rect 33180 19906 33236 19908
rect 33180 19854 33182 19906
rect 33182 19854 33234 19906
rect 33234 19854 33236 19906
rect 33180 19852 33236 19854
rect 32396 19180 32452 19236
rect 32172 18450 32228 18452
rect 32172 18398 32174 18450
rect 32174 18398 32226 18450
rect 32226 18398 32228 18450
rect 32172 18396 32228 18398
rect 32844 18396 32900 18452
rect 32956 17666 33012 17668
rect 32956 17614 32958 17666
rect 32958 17614 33010 17666
rect 33010 17614 33012 17666
rect 32956 17612 33012 17614
rect 32284 17442 32340 17444
rect 32284 17390 32286 17442
rect 32286 17390 32338 17442
rect 32338 17390 32340 17442
rect 32284 17388 32340 17390
rect 32956 17052 33012 17108
rect 33516 18396 33572 18452
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 34636 19068 34692 19124
rect 34524 18396 34580 18452
rect 35644 19122 35700 19124
rect 35644 19070 35646 19122
rect 35646 19070 35698 19122
rect 35698 19070 35700 19122
rect 35644 19068 35700 19070
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 34188 17612 34244 17668
rect 32508 15820 32564 15876
rect 32732 15820 32788 15876
rect 31948 14642 32004 14644
rect 31948 14590 31950 14642
rect 31950 14590 32002 14642
rect 32002 14590 32004 14642
rect 31948 14588 32004 14590
rect 33852 15986 33908 15988
rect 33852 15934 33854 15986
rect 33854 15934 33906 15986
rect 33906 15934 33908 15986
rect 33852 15932 33908 15934
rect 33180 15820 33236 15876
rect 34972 17388 35028 17444
rect 35532 16940 35588 16996
rect 34412 16098 34468 16100
rect 34412 16046 34414 16098
rect 34414 16046 34466 16098
rect 34466 16046 34468 16098
rect 34412 16044 34468 16046
rect 34300 15986 34356 15988
rect 34300 15934 34302 15986
rect 34302 15934 34354 15986
rect 34354 15934 34356 15986
rect 34300 15932 34356 15934
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35644 16268 35700 16324
rect 35868 16604 35924 16660
rect 40012 23324 40068 23380
rect 44044 25618 44100 25620
rect 44044 25566 44046 25618
rect 44046 25566 44098 25618
rect 44098 25566 44100 25618
rect 44044 25564 44100 25566
rect 40012 22482 40068 22484
rect 40012 22430 40014 22482
rect 40014 22430 40066 22482
rect 40066 22430 40068 22482
rect 40012 22428 40068 22430
rect 41020 22428 41076 22484
rect 37100 20188 37156 20244
rect 41692 23436 41748 23492
rect 41804 23660 41860 23716
rect 41580 21756 41636 21812
rect 42588 21810 42644 21812
rect 42588 21758 42590 21810
rect 42590 21758 42642 21810
rect 42642 21758 42644 21810
rect 42588 21756 42644 21758
rect 39788 20188 39844 20244
rect 40348 20188 40404 20244
rect 36428 17500 36484 17556
rect 36988 17554 37044 17556
rect 36988 17502 36990 17554
rect 36990 17502 37042 17554
rect 37042 17502 37044 17554
rect 36988 17500 37044 17502
rect 36092 16098 36148 16100
rect 36092 16046 36094 16098
rect 36094 16046 36146 16098
rect 36146 16046 36148 16098
rect 36092 16044 36148 16046
rect 37324 16156 37380 16212
rect 37436 16268 37492 16324
rect 39564 16210 39620 16212
rect 39564 16158 39566 16210
rect 39566 16158 39618 16210
rect 39618 16158 39620 16210
rect 39564 16156 39620 16158
rect 37100 15874 37156 15876
rect 37100 15822 37102 15874
rect 37102 15822 37154 15874
rect 37154 15822 37156 15874
rect 37100 15820 37156 15822
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 32956 14588 33012 14644
rect 35420 13970 35476 13972
rect 35420 13918 35422 13970
rect 35422 13918 35474 13970
rect 35474 13918 35476 13970
rect 35420 13916 35476 13918
rect 36540 13916 36596 13972
rect 35644 13692 35700 13748
rect 36316 13746 36372 13748
rect 36316 13694 36318 13746
rect 36318 13694 36370 13746
rect 36370 13694 36372 13746
rect 36316 13692 36372 13694
rect 34748 13634 34804 13636
rect 34748 13582 34750 13634
rect 34750 13582 34802 13634
rect 34802 13582 34804 13634
rect 34748 13580 34804 13582
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 36092 13074 36148 13076
rect 36092 13022 36094 13074
rect 36094 13022 36146 13074
rect 36146 13022 36148 13074
rect 36092 13020 36148 13022
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 40348 15820 40404 15876
rect 36988 11900 37044 11956
rect 31724 10834 31780 10836
rect 31724 10782 31726 10834
rect 31726 10782 31778 10834
rect 31778 10782 31780 10834
rect 31724 10780 31780 10782
rect 35196 11170 35252 11172
rect 35196 11118 35198 11170
rect 35198 11118 35250 11170
rect 35250 11118 35252 11170
rect 35196 11116 35252 11118
rect 31388 10050 31444 10052
rect 31388 9998 31390 10050
rect 31390 9998 31442 10050
rect 31442 9998 31444 10050
rect 31388 9996 31444 9998
rect 31052 9884 31108 9940
rect 32060 9884 32116 9940
rect 31836 9826 31892 9828
rect 31836 9774 31838 9826
rect 31838 9774 31890 9826
rect 31890 9774 31892 9826
rect 31836 9772 31892 9774
rect 30828 9714 30884 9716
rect 30828 9662 30830 9714
rect 30830 9662 30882 9714
rect 30882 9662 30884 9714
rect 30828 9660 30884 9662
rect 31948 9714 32004 9716
rect 31948 9662 31950 9714
rect 31950 9662 32002 9714
rect 32002 9662 32004 9714
rect 31948 9660 32004 9662
rect 31388 9548 31444 9604
rect 33964 9826 34020 9828
rect 33964 9774 33966 9826
rect 33966 9774 34018 9826
rect 34018 9774 34020 9826
rect 33964 9772 34020 9774
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 34524 9772 34580 9828
rect 33740 9714 33796 9716
rect 33740 9662 33742 9714
rect 33742 9662 33794 9714
rect 33794 9662 33796 9714
rect 33740 9660 33796 9662
rect 32060 9154 32116 9156
rect 32060 9102 32062 9154
rect 32062 9102 32114 9154
rect 32114 9102 32116 9154
rect 32060 9100 32116 9102
rect 32284 9042 32340 9044
rect 32284 8990 32286 9042
rect 32286 8990 32338 9042
rect 32338 8990 32340 9042
rect 32284 8988 32340 8990
rect 32172 8930 32228 8932
rect 32172 8878 32174 8930
rect 32174 8878 32226 8930
rect 32226 8878 32228 8930
rect 32172 8876 32228 8878
rect 33292 9154 33348 9156
rect 33292 9102 33294 9154
rect 33294 9102 33346 9154
rect 33346 9102 33348 9154
rect 33292 9100 33348 9102
rect 35644 9660 35700 9716
rect 33740 9042 33796 9044
rect 33740 8990 33742 9042
rect 33742 8990 33794 9042
rect 33794 8990 33796 9042
rect 33740 8988 33796 8990
rect 32844 8876 32900 8932
rect 32620 6636 32676 6692
rect 30268 5964 30324 6020
rect 29372 5906 29428 5908
rect 29372 5854 29374 5906
rect 29374 5854 29426 5906
rect 29426 5854 29428 5906
rect 29372 5852 29428 5854
rect 28476 5740 28532 5796
rect 29260 5794 29316 5796
rect 29260 5742 29262 5794
rect 29262 5742 29314 5794
rect 29314 5742 29316 5794
rect 29260 5740 29316 5742
rect 29596 5906 29652 5908
rect 29596 5854 29598 5906
rect 29598 5854 29650 5906
rect 29650 5854 29652 5906
rect 29596 5852 29652 5854
rect 30156 5906 30212 5908
rect 30156 5854 30158 5906
rect 30158 5854 30210 5906
rect 30210 5854 30212 5906
rect 30156 5852 30212 5854
rect 31276 5740 31332 5796
rect 33516 6860 33572 6916
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 34860 8428 34916 8484
rect 36428 8428 36484 8484
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 34860 6636 34916 6692
rect 35196 6860 35252 6916
rect 37660 11116 37716 11172
rect 39116 13074 39172 13076
rect 39116 13022 39118 13074
rect 39118 13022 39170 13074
rect 39170 13022 39172 13074
rect 39116 13020 39172 13022
rect 39788 11900 39844 11956
rect 37996 11116 38052 11172
rect 36988 8428 37044 8484
rect 38108 8428 38164 8484
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 31948 5122 32004 5124
rect 31948 5070 31950 5122
rect 31950 5070 32002 5122
rect 32002 5070 32004 5122
rect 31948 5068 32004 5070
rect 32620 5068 32676 5124
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
<< metal3 >>
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 28466 42140 28476 42196
rect 28532 42140 28542 42196
rect 28476 41972 28532 42140
rect 23202 41916 23212 41972
rect 23268 41916 24892 41972
rect 24948 41916 24958 41972
rect 28476 41916 30380 41972
rect 30436 41916 30446 41972
rect 31378 41916 31388 41972
rect 31444 41916 32508 41972
rect 32564 41916 32574 41972
rect 33730 41916 33740 41972
rect 33796 41916 36316 41972
rect 36372 41916 36382 41972
rect 13234 41804 13244 41860
rect 13300 41804 14476 41860
rect 14532 41804 14542 41860
rect 24658 41804 24668 41860
rect 24724 41804 25900 41860
rect 25956 41804 25966 41860
rect 36082 41804 36092 41860
rect 36148 41804 37324 41860
rect 37380 41804 37390 41860
rect 39890 41804 39900 41860
rect 39956 41804 41132 41860
rect 41188 41804 41198 41860
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 11554 40460 11564 40516
rect 11620 40460 12012 40516
rect 12068 40460 12348 40516
rect 12404 40460 12414 40516
rect 16930 40460 16940 40516
rect 16996 40460 31612 40516
rect 31668 40460 31678 40516
rect 2930 40348 2940 40404
rect 2996 40348 11340 40404
rect 11396 40348 11406 40404
rect 11666 40348 11676 40404
rect 11732 40348 12124 40404
rect 12180 40348 13916 40404
rect 13972 40348 13982 40404
rect 17826 40348 17836 40404
rect 17892 40348 20076 40404
rect 20132 40348 21420 40404
rect 21476 40348 21486 40404
rect 25330 40348 25340 40404
rect 25396 40348 28588 40404
rect 28644 40348 28654 40404
rect 38098 40348 38108 40404
rect 38164 40348 40460 40404
rect 40516 40348 41020 40404
rect 41076 40348 41086 40404
rect 5058 40236 5068 40292
rect 5124 40236 8428 40292
rect 12450 40236 12460 40292
rect 12516 40236 21084 40292
rect 21140 40236 21150 40292
rect 40338 40236 40348 40292
rect 40404 40236 41804 40292
rect 41860 40236 41870 40292
rect 42690 40236 42700 40292
rect 42756 40236 43932 40292
rect 43988 40236 43998 40292
rect 8372 40180 8428 40236
rect 8372 40124 13468 40180
rect 13524 40124 13534 40180
rect 14690 40124 14700 40180
rect 14756 40124 15484 40180
rect 15540 40124 15550 40180
rect 8978 40012 8988 40068
rect 9044 40012 17276 40068
rect 17332 40012 17342 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 16034 39676 16044 39732
rect 16100 39676 29260 39732
rect 29316 39676 29326 39732
rect 10994 39564 11004 39620
rect 11060 39564 12572 39620
rect 12628 39564 14252 39620
rect 14308 39564 14318 39620
rect 15586 39564 15596 39620
rect 15652 39564 18620 39620
rect 18676 39564 18686 39620
rect 28354 39564 28364 39620
rect 28420 39564 30268 39620
rect 30324 39564 30940 39620
rect 30996 39564 31948 39620
rect 32004 39564 34188 39620
rect 34244 39564 34254 39620
rect 8306 39452 8316 39508
rect 8372 39396 8428 39508
rect 12674 39452 12684 39508
rect 12740 39452 14028 39508
rect 14084 39452 14364 39508
rect 14420 39452 14812 39508
rect 14868 39452 14878 39508
rect 15810 39452 15820 39508
rect 15876 39452 16828 39508
rect 16884 39452 16894 39508
rect 8372 39340 10668 39396
rect 10724 39340 10734 39396
rect 14578 39340 14588 39396
rect 14644 39340 16380 39396
rect 16436 39340 16446 39396
rect 16930 39340 16940 39396
rect 16996 39340 26012 39396
rect 26068 39340 26078 39396
rect 39666 39340 39676 39396
rect 39732 39340 41132 39396
rect 41188 39340 41198 39396
rect 7186 39228 7196 39284
rect 7252 39228 11900 39284
rect 11956 39228 15148 39284
rect 15204 39228 16156 39284
rect 16212 39228 17052 39284
rect 17108 39228 17118 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 12002 39004 12012 39060
rect 12068 39004 15708 39060
rect 15764 39004 15932 39060
rect 15988 39004 15998 39060
rect 2706 38892 2716 38948
rect 2772 38892 11676 38948
rect 11732 38892 12572 38948
rect 12628 38892 12638 38948
rect 13804 38892 14924 38948
rect 14980 38892 14990 38948
rect 13804 38836 13860 38892
rect 10322 38780 10332 38836
rect 10388 38780 13804 38836
rect 13860 38780 13870 38836
rect 14018 38780 14028 38836
rect 14084 38780 15036 38836
rect 15092 38780 15596 38836
rect 15652 38780 15662 38836
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 22754 38108 22764 38164
rect 22820 38108 26012 38164
rect 26068 38108 28364 38164
rect 28420 38108 28430 38164
rect 39414 37996 39452 38052
rect 39508 37996 39518 38052
rect 36978 37884 36988 37940
rect 37044 37884 39900 37940
rect 39956 37884 39966 37940
rect 2258 37772 2268 37828
rect 2324 37772 3052 37828
rect 3108 37772 5740 37828
rect 5796 37772 6300 37828
rect 6356 37772 9772 37828
rect 9828 37772 9838 37828
rect 35298 37772 35308 37828
rect 35364 37772 37436 37828
rect 37492 37772 37502 37828
rect 39778 37772 39788 37828
rect 39844 37772 41916 37828
rect 41972 37772 41982 37828
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 37314 37436 37324 37492
rect 37380 37436 39788 37492
rect 39844 37436 42588 37492
rect 42644 37436 42654 37492
rect 3714 37324 3724 37380
rect 3780 37324 10332 37380
rect 10388 37324 10398 37380
rect 11218 37212 11228 37268
rect 11284 37212 11788 37268
rect 11844 37212 12236 37268
rect 12292 37212 12302 37268
rect 31602 37212 31612 37268
rect 31668 37212 32060 37268
rect 32116 37212 35308 37268
rect 35364 37212 35374 37268
rect 39218 37212 39228 37268
rect 39284 37212 39564 37268
rect 39620 37212 39630 37268
rect 11554 37100 11564 37156
rect 11620 37100 12460 37156
rect 12516 37100 14476 37156
rect 14532 37100 16716 37156
rect 16772 37100 20300 37156
rect 20356 37100 20366 37156
rect 10994 36988 11004 37044
rect 11060 36988 11676 37044
rect 11732 36988 12348 37044
rect 12404 36988 14588 37044
rect 14644 36988 14654 37044
rect 34412 36988 36988 37044
rect 37044 36988 37054 37044
rect 34412 36932 34468 36988
rect 34402 36876 34412 36932
rect 34468 36876 34478 36932
rect 38546 36876 38556 36932
rect 38612 36876 39900 36932
rect 39956 36876 40236 36932
rect 40292 36876 40302 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 6514 36764 6524 36820
rect 6580 36764 12012 36820
rect 12068 36764 13468 36820
rect 13524 36764 13534 36820
rect 38556 36708 38612 36876
rect 24546 36652 24556 36708
rect 24612 36652 25564 36708
rect 25620 36652 26460 36708
rect 26516 36652 28700 36708
rect 28756 36652 32284 36708
rect 32340 36652 32350 36708
rect 33506 36652 33516 36708
rect 33572 36652 35420 36708
rect 35476 36652 38612 36708
rect 5842 36540 5852 36596
rect 5908 36540 6972 36596
rect 7028 36540 7038 36596
rect 9986 36540 9996 36596
rect 10052 36540 12348 36596
rect 12404 36540 12414 36596
rect 12898 36540 12908 36596
rect 12964 36540 13804 36596
rect 13860 36540 15596 36596
rect 15652 36540 15662 36596
rect 30818 36540 30828 36596
rect 30884 36540 33852 36596
rect 33908 36540 33918 36596
rect 39414 36540 39452 36596
rect 39508 36540 39518 36596
rect 12562 36428 12572 36484
rect 12628 36428 13244 36484
rect 13300 36428 13310 36484
rect 13458 36428 13468 36484
rect 13524 36428 15036 36484
rect 15092 36428 15484 36484
rect 15540 36428 18004 36484
rect 18386 36428 18396 36484
rect 18452 36428 19068 36484
rect 19124 36428 20972 36484
rect 21028 36428 21038 36484
rect 39330 36428 39340 36484
rect 39396 36428 40348 36484
rect 40404 36428 44044 36484
rect 44100 36428 44110 36484
rect 17948 36372 18004 36428
rect 13682 36316 13692 36372
rect 13748 36316 16268 36372
rect 16324 36316 17724 36372
rect 17780 36316 17790 36372
rect 17948 36316 19628 36372
rect 19684 36316 19964 36372
rect 20020 36316 20748 36372
rect 20804 36316 20814 36372
rect 21746 36316 21756 36372
rect 21812 36316 24108 36372
rect 24164 36316 24174 36372
rect 34962 36316 34972 36372
rect 35028 36316 36652 36372
rect 36708 36316 36718 36372
rect 7074 36204 7084 36260
rect 7140 36204 10220 36260
rect 10276 36204 10286 36260
rect 32386 36204 32396 36260
rect 32452 36204 33852 36260
rect 33908 36204 34636 36260
rect 34692 36204 34702 36260
rect 37090 36204 37100 36260
rect 37156 36204 39116 36260
rect 39172 36204 39182 36260
rect 40002 36204 40012 36260
rect 40068 36204 40572 36260
rect 40628 36204 40638 36260
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 37426 35980 37436 36036
rect 37492 35980 38780 36036
rect 38836 35980 38846 36036
rect 40114 35980 40124 36036
rect 40180 35980 40908 36036
rect 40964 35980 40974 36036
rect 4834 35756 4844 35812
rect 4900 35756 13020 35812
rect 13076 35756 13086 35812
rect 20290 35756 20300 35812
rect 20356 35756 21756 35812
rect 21812 35756 21822 35812
rect 13234 35644 13244 35700
rect 13300 35644 13916 35700
rect 13972 35644 17276 35700
rect 17332 35644 17342 35700
rect 18386 35644 18396 35700
rect 18452 35644 20076 35700
rect 20132 35644 25228 35700
rect 25284 35644 25294 35700
rect 36530 35644 36540 35700
rect 36596 35644 37548 35700
rect 37604 35644 39564 35700
rect 39620 35644 39630 35700
rect 15026 35532 15036 35588
rect 15092 35532 18060 35588
rect 18116 35532 18126 35588
rect 27346 35532 27356 35588
rect 27412 35532 34636 35588
rect 34692 35532 37324 35588
rect 37380 35532 37390 35588
rect 16706 35420 16716 35476
rect 16772 35420 18844 35476
rect 18900 35420 18910 35476
rect 23426 35420 23436 35476
rect 23492 35420 24220 35476
rect 24276 35420 24286 35476
rect 10322 35308 10332 35364
rect 10388 35308 14252 35364
rect 14308 35308 14700 35364
rect 14756 35308 14766 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 18610 35084 18620 35140
rect 18676 35084 19180 35140
rect 19236 35084 19852 35140
rect 19908 35084 19918 35140
rect 26012 34972 29036 35028
rect 29092 34972 29102 35028
rect 26012 34916 26068 34972
rect 21634 34860 21644 34916
rect 21700 34860 26012 34916
rect 26068 34860 26078 34916
rect 28354 34860 28364 34916
rect 28420 34860 29372 34916
rect 29428 34860 31948 34916
rect 32004 34860 35084 34916
rect 35140 34860 35150 34916
rect 14802 34748 14812 34804
rect 14868 34748 15148 34804
rect 18386 34748 18396 34804
rect 18452 34748 19516 34804
rect 19572 34748 19582 34804
rect 15092 34692 15148 34748
rect 15092 34636 18956 34692
rect 19012 34636 19022 34692
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 19170 34300 19180 34356
rect 19236 34300 20076 34356
rect 20132 34020 20188 34356
rect 20132 33964 27468 34020
rect 27524 33964 27534 34020
rect 40898 33740 40908 33796
rect 40964 33740 41580 33796
rect 41636 33740 44044 33796
rect 44100 33740 44110 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 37426 33516 37436 33572
rect 37492 33516 39116 33572
rect 39172 33516 39182 33572
rect 6626 33404 6636 33460
rect 6692 33404 8988 33460
rect 9044 33404 9054 33460
rect 32274 33292 32284 33348
rect 32340 33292 33180 33348
rect 33236 33292 34076 33348
rect 34132 33292 34142 33348
rect 27346 33068 27356 33124
rect 27412 33068 29372 33124
rect 29428 33068 29438 33124
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 8978 32732 8988 32788
rect 9044 32732 9772 32788
rect 9828 32732 9838 32788
rect 8418 32620 8428 32676
rect 8484 32620 10444 32676
rect 10500 32620 10510 32676
rect 24658 32620 24668 32676
rect 24724 32620 25228 32676
rect 25284 32620 32284 32676
rect 32340 32620 32350 32676
rect 32498 32620 32508 32676
rect 32564 32620 34300 32676
rect 34356 32620 39228 32676
rect 39284 32620 40236 32676
rect 40292 32620 40302 32676
rect 24210 32508 24220 32564
rect 24276 32508 25340 32564
rect 25396 32508 25406 32564
rect 33506 32508 33516 32564
rect 33572 32508 35532 32564
rect 35588 32508 36428 32564
rect 36484 32508 36876 32564
rect 36932 32508 36942 32564
rect 34738 32396 34748 32452
rect 34804 32396 35980 32452
rect 36036 32396 37660 32452
rect 37716 32396 37726 32452
rect 25442 32284 25452 32340
rect 25508 32284 28140 32340
rect 28196 32284 29148 32340
rect 29204 32284 29214 32340
rect 33394 32172 33404 32228
rect 33460 32172 33852 32228
rect 33908 32172 33918 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 9986 31836 9996 31892
rect 10052 31836 16380 31892
rect 16436 31836 16828 31892
rect 16884 31836 16894 31892
rect 33282 31836 33292 31892
rect 33348 31836 40460 31892
rect 40516 31836 41132 31892
rect 41188 31836 41198 31892
rect 2258 31724 2268 31780
rect 2324 31724 2716 31780
rect 2772 31724 5964 31780
rect 6020 31724 6030 31780
rect 34402 31724 34412 31780
rect 34468 31724 39340 31780
rect 39396 31724 39406 31780
rect 24098 31612 24108 31668
rect 24164 31612 24780 31668
rect 24836 31612 24846 31668
rect 33506 31500 33516 31556
rect 33572 31500 34972 31556
rect 35028 31500 35038 31556
rect 36530 31500 36540 31556
rect 36596 31500 36988 31556
rect 37044 31500 37054 31556
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 5730 31052 5740 31108
rect 5796 31052 5964 31108
rect 6020 31052 10444 31108
rect 10500 31052 10510 31108
rect 15474 30940 15484 30996
rect 15540 30940 16492 30996
rect 16548 30940 16558 30996
rect 18284 30940 21420 30996
rect 21476 30940 21486 30996
rect 18284 30884 18340 30940
rect 3378 30828 3388 30884
rect 3444 30828 4956 30884
rect 5012 30828 5022 30884
rect 16818 30828 16828 30884
rect 16884 30828 18284 30884
rect 18340 30828 18350 30884
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 6626 30380 6636 30436
rect 6692 30380 8092 30436
rect 8148 30380 8764 30436
rect 8820 30380 8830 30436
rect 33058 30380 33068 30436
rect 33124 30380 34636 30436
rect 34692 30380 34702 30436
rect 9090 30268 9100 30324
rect 9156 30268 12012 30324
rect 12068 30268 12078 30324
rect 33170 30268 33180 30324
rect 33236 30268 34188 30324
rect 34244 30268 34254 30324
rect 5842 30156 5852 30212
rect 5908 30156 10108 30212
rect 10164 30156 11900 30212
rect 11956 30156 11966 30212
rect 24882 30156 24892 30212
rect 24948 30156 25676 30212
rect 25732 30156 26908 30212
rect 26964 30156 26974 30212
rect 37090 30156 37100 30212
rect 37156 30156 40348 30212
rect 40404 30156 40414 30212
rect 15922 30044 15932 30100
rect 15988 30044 17500 30100
rect 17556 30044 17566 30100
rect 42690 30044 42700 30100
rect 42756 30044 44044 30100
rect 44100 30044 44110 30100
rect 16034 29932 16044 29988
rect 16100 29932 16492 29988
rect 16548 29932 20300 29988
rect 20356 29932 26236 29988
rect 26292 29932 29372 29988
rect 29428 29932 29932 29988
rect 29988 29932 32620 29988
rect 32676 29932 32686 29988
rect 38994 29932 39004 29988
rect 39060 29932 41468 29988
rect 41524 29932 42588 29988
rect 42644 29932 42654 29988
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 34514 29708 34524 29764
rect 34580 29708 35756 29764
rect 35812 29708 37660 29764
rect 37716 29708 40796 29764
rect 40852 29708 40862 29764
rect 6962 29596 6972 29652
rect 7028 29596 28588 29652
rect 28644 29596 28654 29652
rect 37538 29596 37548 29652
rect 37604 29596 38892 29652
rect 38948 29596 38958 29652
rect 40338 29596 40348 29652
rect 40404 29596 41132 29652
rect 41188 29596 41198 29652
rect 9996 29484 12124 29540
rect 12180 29484 12190 29540
rect 14466 29484 14476 29540
rect 14532 29484 16156 29540
rect 16212 29484 18620 29540
rect 18676 29484 18686 29540
rect 36642 29484 36652 29540
rect 36708 29484 37212 29540
rect 37268 29484 38668 29540
rect 38724 29484 38734 29540
rect 9996 29428 10052 29484
rect 3378 29372 3388 29428
rect 3444 29372 4620 29428
rect 4676 29372 4686 29428
rect 5618 29372 5628 29428
rect 5684 29372 9996 29428
rect 10052 29372 10062 29428
rect 11442 29372 11452 29428
rect 11508 29372 13916 29428
rect 13972 29372 14364 29428
rect 14420 29372 14430 29428
rect 15474 29372 15484 29428
rect 15540 29372 17500 29428
rect 17556 29372 17566 29428
rect 18162 29372 18172 29428
rect 18228 29372 19292 29428
rect 19348 29372 19358 29428
rect 4620 29316 4676 29372
rect 4620 29260 6076 29316
rect 6132 29260 6142 29316
rect 11554 29260 11564 29316
rect 11620 29260 15596 29316
rect 15652 29260 19068 29316
rect 19124 29260 19134 29316
rect 23538 29260 23548 29316
rect 23604 29260 25340 29316
rect 25396 29260 25406 29316
rect 25554 29260 25564 29316
rect 25620 29260 26012 29316
rect 26068 29260 26684 29316
rect 26740 29260 28812 29316
rect 28868 29260 29372 29316
rect 29428 29260 40460 29316
rect 40516 29260 40526 29316
rect 4284 29148 4396 29204
rect 4452 29148 4462 29204
rect 9874 29148 9884 29204
rect 9940 29148 11676 29204
rect 11732 29148 11742 29204
rect 12124 29148 15484 29204
rect 15540 29148 15550 29204
rect 33170 29148 33180 29204
rect 33236 29148 33740 29204
rect 33796 29148 33806 29204
rect 34178 29148 34188 29204
rect 34244 29148 37548 29204
rect 37604 29148 37614 29204
rect 3266 28924 3276 28980
rect 3332 28924 3836 28980
rect 3892 28924 3902 28980
rect 4284 28868 4340 29148
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 12124 28980 12180 29148
rect 15922 29036 15932 29092
rect 15988 29036 16268 29092
rect 16324 29036 16334 29092
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 5058 28924 5068 28980
rect 5124 28924 6300 28980
rect 6356 28924 10780 28980
rect 10836 28924 12180 28980
rect 14924 28924 15708 28980
rect 15764 28924 16380 28980
rect 16436 28924 17388 28980
rect 17444 28924 17454 28980
rect 20132 28924 23996 28980
rect 24052 28924 24062 28980
rect 14924 28868 14980 28924
rect 4284 28812 4396 28868
rect 4452 28812 6412 28868
rect 6468 28812 6478 28868
rect 9650 28812 9660 28868
rect 9716 28812 14980 28868
rect 20132 28756 20188 28924
rect 28578 28812 28588 28868
rect 28644 28812 29372 28868
rect 29428 28812 35084 28868
rect 35140 28812 35980 28868
rect 36036 28812 36046 28868
rect 4050 28700 4060 28756
rect 4116 28700 8876 28756
rect 8932 28700 9548 28756
rect 9604 28700 9614 28756
rect 10882 28700 10892 28756
rect 10948 28700 15932 28756
rect 15988 28700 17276 28756
rect 17332 28700 17892 28756
rect 18050 28700 18060 28756
rect 18116 28700 18396 28756
rect 18452 28700 20188 28756
rect 31042 28700 31052 28756
rect 31108 28700 33852 28756
rect 33908 28700 33918 28756
rect 40002 28700 40012 28756
rect 40068 28700 41580 28756
rect 41636 28700 41646 28756
rect 17836 28644 17892 28700
rect 3154 28588 3164 28644
rect 3220 28588 3612 28644
rect 3668 28588 3678 28644
rect 4498 28588 4508 28644
rect 4564 28588 4574 28644
rect 4722 28588 4732 28644
rect 4788 28588 5964 28644
rect 6020 28588 7980 28644
rect 8036 28588 8046 28644
rect 8726 28588 8764 28644
rect 8820 28588 9884 28644
rect 9940 28588 9950 28644
rect 11218 28588 11228 28644
rect 11284 28588 12572 28644
rect 12628 28588 12638 28644
rect 14018 28588 14028 28644
rect 14084 28588 15148 28644
rect 15204 28588 16044 28644
rect 16100 28588 17612 28644
rect 17668 28588 17678 28644
rect 17836 28588 18508 28644
rect 18564 28588 18574 28644
rect 22866 28588 22876 28644
rect 22932 28588 26124 28644
rect 26180 28588 30268 28644
rect 30324 28588 31388 28644
rect 31444 28588 31454 28644
rect 40450 28588 40460 28644
rect 40516 28588 41132 28644
rect 41188 28588 41198 28644
rect 4508 28532 4564 28588
rect 3490 28476 3500 28532
rect 3556 28476 4284 28532
rect 4340 28476 4350 28532
rect 4508 28476 5068 28532
rect 5124 28476 5134 28532
rect 6514 28476 6524 28532
rect 6580 28476 6972 28532
rect 7028 28476 7038 28532
rect 8306 28476 8316 28532
rect 8372 28476 9212 28532
rect 9268 28476 10108 28532
rect 10164 28476 10174 28532
rect 12002 28476 12012 28532
rect 12068 28476 12078 28532
rect 12786 28476 12796 28532
rect 12852 28476 13580 28532
rect 13636 28476 13646 28532
rect 15092 28476 18844 28532
rect 18900 28476 18910 28532
rect 28242 28476 28252 28532
rect 28308 28476 32508 28532
rect 32564 28476 32574 28532
rect 4284 28420 4340 28476
rect 12012 28420 12068 28476
rect 15092 28420 15148 28476
rect 4284 28364 4508 28420
rect 4564 28364 4956 28420
rect 5012 28364 5022 28420
rect 5618 28364 5628 28420
rect 5684 28364 5964 28420
rect 6020 28364 6030 28420
rect 12012 28364 15148 28420
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 8194 28028 8204 28084
rect 8260 28028 9996 28084
rect 10052 28028 10892 28084
rect 10948 28028 10958 28084
rect 15092 27916 18060 27972
rect 18116 27916 18126 27972
rect 15092 27860 15148 27916
rect 3714 27804 3724 27860
rect 3780 27804 4732 27860
rect 4788 27804 5964 27860
rect 6020 27804 6030 27860
rect 12114 27804 12124 27860
rect 12180 27804 13468 27860
rect 13524 27804 15148 27860
rect 4274 27692 4284 27748
rect 4340 27692 5292 27748
rect 5348 27692 5358 27748
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 12562 27356 12572 27412
rect 12628 27356 26348 27412
rect 26404 27356 26414 27412
rect 20626 27244 20636 27300
rect 20692 27244 39900 27300
rect 39956 27244 39966 27300
rect 10658 27132 10668 27188
rect 10724 27132 14140 27188
rect 14196 27132 15260 27188
rect 15316 27132 15326 27188
rect 16146 27132 16156 27188
rect 16212 27132 17836 27188
rect 17892 27132 17902 27188
rect 21970 27132 21980 27188
rect 22036 27132 22540 27188
rect 22596 27132 25452 27188
rect 25508 27132 25900 27188
rect 25956 27132 36428 27188
rect 36484 27132 36764 27188
rect 36820 27132 37100 27188
rect 37156 27132 37166 27188
rect 20178 27020 20188 27076
rect 20244 27020 21756 27076
rect 21812 27020 27132 27076
rect 27188 27020 28252 27076
rect 28308 27020 28318 27076
rect 40226 27020 40236 27076
rect 40292 27020 40796 27076
rect 40852 27020 40862 27076
rect 17714 26908 17724 26964
rect 17780 26908 18060 26964
rect 18116 26908 18126 26964
rect 18834 26908 18844 26964
rect 18900 26908 20524 26964
rect 20580 26908 20590 26964
rect 21298 26908 21308 26964
rect 21364 26908 22204 26964
rect 22260 26908 22270 26964
rect 28354 26908 28364 26964
rect 28420 26908 29484 26964
rect 29540 26908 29550 26964
rect 29810 26908 29820 26964
rect 29876 26908 30268 26964
rect 30324 26908 30334 26964
rect 37650 26908 37660 26964
rect 37716 26908 38780 26964
rect 38836 26908 39452 26964
rect 39508 26908 40124 26964
rect 40180 26908 40190 26964
rect 12674 26796 12684 26852
rect 12740 26796 15596 26852
rect 15652 26796 15662 26852
rect 17266 26796 17276 26852
rect 17332 26796 17948 26852
rect 18004 26796 18508 26852
rect 18564 26796 18574 26852
rect 35298 26796 35308 26852
rect 35364 26796 36876 26852
rect 36932 26796 36942 26852
rect 3826 26684 3836 26740
rect 3892 26684 10780 26740
rect 10836 26684 10846 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 8978 26572 8988 26628
rect 9044 26572 14476 26628
rect 14532 26572 14542 26628
rect 14354 26460 14364 26516
rect 14420 26460 15260 26516
rect 15316 26460 15326 26516
rect 18274 26460 18284 26516
rect 18340 26460 19852 26516
rect 19908 26460 20188 26516
rect 37202 26460 37212 26516
rect 37268 26460 38220 26516
rect 38276 26460 38286 26516
rect 6402 26348 6412 26404
rect 6468 26348 10108 26404
rect 10164 26348 12236 26404
rect 12292 26348 12302 26404
rect 18050 26348 18060 26404
rect 18116 26348 19180 26404
rect 19236 26348 19246 26404
rect 9762 26236 9772 26292
rect 9828 26236 11116 26292
rect 11172 26236 12684 26292
rect 12740 26236 12750 26292
rect 14914 26236 14924 26292
rect 14980 26236 16044 26292
rect 16100 26236 16110 26292
rect 16258 26236 16268 26292
rect 16324 26236 17388 26292
rect 17444 26236 17454 26292
rect 18162 26236 18172 26292
rect 18228 26236 18956 26292
rect 19012 26236 19022 26292
rect 20132 26236 20188 26460
rect 20244 26236 20254 26292
rect 36866 26236 36876 26292
rect 36932 26236 37436 26292
rect 37492 26236 37502 26292
rect 16146 26124 16156 26180
rect 16212 26124 22876 26180
rect 22932 26124 22942 26180
rect 26786 26124 26796 26180
rect 26852 26124 30044 26180
rect 30100 26124 30110 26180
rect 35858 26124 35868 26180
rect 35924 26124 37324 26180
rect 37380 26124 37390 26180
rect 18722 26012 18732 26068
rect 18788 26012 23100 26068
rect 23156 26012 23166 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 10770 25676 10780 25732
rect 10836 25676 12236 25732
rect 12292 25676 12302 25732
rect 34738 25676 34748 25732
rect 34804 25676 35420 25732
rect 35476 25676 35486 25732
rect 8306 25564 8316 25620
rect 8372 25564 8876 25620
rect 8932 25564 8942 25620
rect 33954 25564 33964 25620
rect 34020 25564 37212 25620
rect 37268 25564 39900 25620
rect 39956 25564 41132 25620
rect 41188 25564 41198 25620
rect 43652 25564 44044 25620
rect 44100 25564 44110 25620
rect 43652 25508 43708 25564
rect 11778 25452 11788 25508
rect 11844 25452 14364 25508
rect 14420 25452 14430 25508
rect 21522 25452 21532 25508
rect 21588 25452 24220 25508
rect 24276 25452 24892 25508
rect 24948 25452 29820 25508
rect 29876 25452 29886 25508
rect 33842 25452 33852 25508
rect 33908 25452 35084 25508
rect 35140 25452 35150 25508
rect 40450 25452 40460 25508
rect 40516 25452 43708 25508
rect 17154 25340 17164 25396
rect 17220 25340 18172 25396
rect 18228 25340 20188 25396
rect 20132 25284 20188 25340
rect 21532 25284 21588 25452
rect 22754 25340 22764 25396
rect 22820 25340 24444 25396
rect 24500 25340 24510 25396
rect 27794 25340 27804 25396
rect 27860 25340 29260 25396
rect 29316 25340 29326 25396
rect 35186 25340 35196 25396
rect 35252 25340 36764 25396
rect 36820 25340 36830 25396
rect 38210 25340 38220 25396
rect 38276 25340 40684 25396
rect 40740 25340 40750 25396
rect 2930 25228 2940 25284
rect 2996 25228 5740 25284
rect 5796 25228 5806 25284
rect 6178 25228 6188 25284
rect 6244 25228 6748 25284
rect 6804 25228 6814 25284
rect 16370 25228 16380 25284
rect 16436 25228 18732 25284
rect 18788 25228 18798 25284
rect 20132 25228 21588 25284
rect 22866 25228 22876 25284
rect 22932 25228 27468 25284
rect 27524 25228 27534 25284
rect 29698 25228 29708 25284
rect 29764 25228 30156 25284
rect 30212 25228 39676 25284
rect 39732 25228 39742 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 8194 24780 8204 24836
rect 8260 24780 8764 24836
rect 8820 24780 12460 24836
rect 12516 24780 12526 24836
rect 14466 24668 14476 24724
rect 14532 24668 15148 24724
rect 15204 24668 15214 24724
rect 32722 24668 32732 24724
rect 32788 24668 33180 24724
rect 33236 24668 33246 24724
rect 27682 24556 27692 24612
rect 27748 24556 28476 24612
rect 28532 24556 28542 24612
rect 31714 24556 31724 24612
rect 31780 24556 33516 24612
rect 33572 24556 33582 24612
rect 3154 24444 3164 24500
rect 3220 24444 3724 24500
rect 3780 24444 3790 24500
rect 8978 24332 8988 24388
rect 9044 24332 10556 24388
rect 10612 24332 10622 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 5058 23996 5068 24052
rect 5124 23996 6860 24052
rect 6916 23996 7308 24052
rect 7364 23996 7374 24052
rect 21074 23996 21084 24052
rect 21140 23996 23436 24052
rect 23492 23996 23884 24052
rect 23940 23996 24332 24052
rect 24388 23996 24892 24052
rect 24948 23996 24958 24052
rect 31892 23996 34300 24052
rect 34356 23996 34366 24052
rect 35522 23996 35532 24052
rect 35588 23996 35868 24052
rect 35924 23996 39116 24052
rect 39172 23996 40124 24052
rect 40180 23996 40190 24052
rect 31892 23940 31948 23996
rect 2258 23884 2268 23940
rect 2324 23884 5852 23940
rect 5908 23884 5918 23940
rect 18946 23884 18956 23940
rect 19012 23884 19292 23940
rect 19348 23884 19358 23940
rect 30258 23884 30268 23940
rect 30324 23884 31052 23940
rect 31108 23884 31948 23940
rect 7410 23660 7420 23716
rect 7476 23660 8428 23716
rect 8484 23660 8494 23716
rect 28466 23660 28476 23716
rect 28532 23660 29484 23716
rect 29540 23660 40684 23716
rect 40740 23660 41804 23716
rect 41860 23660 41870 23716
rect 40338 23548 40348 23604
rect 40404 23548 40414 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 40348 23492 40404 23548
rect 20178 23436 20188 23492
rect 20244 23436 22876 23492
rect 22932 23436 22942 23492
rect 26002 23436 26012 23492
rect 26068 23436 33292 23492
rect 33348 23436 33358 23492
rect 36754 23436 36764 23492
rect 36820 23436 41692 23492
rect 41748 23436 41758 23492
rect 15026 23324 15036 23380
rect 15092 23324 15372 23380
rect 15428 23324 15438 23380
rect 20402 23324 20412 23380
rect 20468 23324 21532 23380
rect 21588 23324 21598 23380
rect 22642 23324 22652 23380
rect 22708 23324 23548 23380
rect 23604 23324 28924 23380
rect 28980 23324 28990 23380
rect 29922 23324 29932 23380
rect 29988 23324 40012 23380
rect 40068 23324 40078 23380
rect 2482 23100 2492 23156
rect 2548 23100 3388 23156
rect 5282 23100 5292 23156
rect 5348 23100 6860 23156
rect 6916 23100 7644 23156
rect 7700 23100 7710 23156
rect 11330 23100 11340 23156
rect 11396 23100 12684 23156
rect 12740 23100 12750 23156
rect 19842 23100 19852 23156
rect 19908 23100 20748 23156
rect 20804 23100 20814 23156
rect 3332 23044 3388 23100
rect 22652 23044 22708 23324
rect 29138 23212 29148 23268
rect 29204 23212 33068 23268
rect 33124 23212 33134 23268
rect 24434 23100 24444 23156
rect 24500 23100 25676 23156
rect 25732 23100 26348 23156
rect 26404 23100 26414 23156
rect 33170 23100 33180 23156
rect 33236 23100 33852 23156
rect 33908 23100 34972 23156
rect 35028 23100 35038 23156
rect 38434 23100 38444 23156
rect 38500 23100 39452 23156
rect 39508 23100 39518 23156
rect 3332 22988 5852 23044
rect 5908 22988 5918 23044
rect 17266 22988 17276 23044
rect 17332 22988 22708 23044
rect 23874 22988 23884 23044
rect 23940 22988 23950 23044
rect 23884 22932 23940 22988
rect 6402 22876 6412 22932
rect 6468 22876 23940 22932
rect 19170 22764 19180 22820
rect 19236 22764 19740 22820
rect 19796 22764 21084 22820
rect 21140 22764 21150 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 14476 22652 15932 22708
rect 15988 22652 15998 22708
rect 5394 22316 5404 22372
rect 5460 22316 13468 22372
rect 13524 22316 13534 22372
rect 14476 22260 14532 22652
rect 15698 22540 15708 22596
rect 15764 22540 17164 22596
rect 17220 22540 17230 22596
rect 18834 22540 18844 22596
rect 18900 22540 19404 22596
rect 19460 22540 19470 22596
rect 15138 22428 15148 22484
rect 15204 22428 15932 22484
rect 15988 22428 15998 22484
rect 25554 22428 25564 22484
rect 25620 22428 26236 22484
rect 26292 22428 26302 22484
rect 40002 22428 40012 22484
rect 40068 22428 41020 22484
rect 41076 22428 41086 22484
rect 15362 22316 15372 22372
rect 15428 22316 17164 22372
rect 17220 22316 17230 22372
rect 13010 22204 13020 22260
rect 13076 22204 14476 22260
rect 14532 22204 14542 22260
rect 17042 22204 17052 22260
rect 17108 22204 18844 22260
rect 18900 22204 18910 22260
rect 1810 22092 1820 22148
rect 1876 22092 21532 22148
rect 21588 22092 21598 22148
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 3602 21868 3612 21924
rect 3668 21868 6412 21924
rect 6468 21868 6478 21924
rect 13570 21756 13580 21812
rect 13636 21756 17052 21812
rect 17108 21756 17118 21812
rect 25218 21756 25228 21812
rect 25284 21756 25788 21812
rect 25844 21756 26236 21812
rect 26292 21756 26572 21812
rect 26628 21756 26638 21812
rect 41570 21756 41580 21812
rect 41636 21756 42588 21812
rect 42644 21756 42654 21812
rect 19058 21644 19068 21700
rect 19124 21644 28924 21700
rect 28980 21644 28990 21700
rect 29586 21644 29596 21700
rect 29652 21644 30604 21700
rect 30660 21644 30670 21700
rect 7410 21532 7420 21588
rect 7476 21532 11340 21588
rect 11396 21532 11406 21588
rect 30146 21532 30156 21588
rect 30212 21532 35980 21588
rect 36036 21532 36046 21588
rect 6738 21308 6748 21364
rect 6804 21308 25228 21364
rect 25284 21308 25900 21364
rect 25956 21308 25966 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 9986 20748 9996 20804
rect 10052 20748 10892 20804
rect 10948 20748 10958 20804
rect 11330 20636 11340 20692
rect 11396 20636 15036 20692
rect 15092 20636 15102 20692
rect 9314 20524 9324 20580
rect 9380 20524 14028 20580
rect 14084 20524 14094 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 11218 20188 11228 20244
rect 11284 20188 13692 20244
rect 13748 20188 13758 20244
rect 30482 20188 30492 20244
rect 30548 20188 31276 20244
rect 31332 20188 31342 20244
rect 37090 20188 37100 20244
rect 37156 20188 39788 20244
rect 39844 20188 40348 20244
rect 40404 20188 40414 20244
rect 8530 20076 8540 20132
rect 8596 20076 10220 20132
rect 10276 20076 10286 20132
rect 8866 19964 8876 20020
rect 8932 19964 14588 20020
rect 14644 19964 14654 20020
rect 19058 19964 19068 20020
rect 19124 19964 19740 20020
rect 19796 19964 19806 20020
rect 28018 19964 28028 20020
rect 28084 19964 29484 20020
rect 29540 19964 31948 20020
rect 31892 19908 31948 19964
rect 5058 19852 5068 19908
rect 5124 19852 5852 19908
rect 5908 19852 5918 19908
rect 10210 19852 10220 19908
rect 10276 19852 10892 19908
rect 10948 19852 11452 19908
rect 11508 19852 11518 19908
rect 31892 19852 33180 19908
rect 33236 19852 33246 19908
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 4722 19292 4732 19348
rect 4788 19292 6076 19348
rect 6132 19292 8428 19348
rect 8484 19292 8494 19348
rect 11442 19292 11452 19348
rect 11508 19292 17836 19348
rect 17892 19292 20188 19348
rect 20244 19292 20254 19348
rect 24770 19292 24780 19348
rect 24836 19292 28028 19348
rect 28084 19292 28094 19348
rect 31714 19180 31724 19236
rect 31780 19180 32396 19236
rect 32452 19180 32462 19236
rect 24322 19068 24332 19124
rect 24388 19068 25452 19124
rect 25508 19068 25518 19124
rect 34626 19068 34636 19124
rect 34692 19068 35644 19124
rect 35700 19068 35710 19124
rect 25218 18956 25228 19012
rect 25284 18956 29820 19012
rect 29876 18956 30268 19012
rect 30324 18956 30334 19012
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 30594 18732 30604 18788
rect 30660 18732 31612 18788
rect 31668 18732 31678 18788
rect 10210 18620 10220 18676
rect 10276 18620 10668 18676
rect 10724 18620 11228 18676
rect 11284 18620 11294 18676
rect 14242 18620 14252 18676
rect 14308 18620 14812 18676
rect 14868 18620 14878 18676
rect 1810 18508 1820 18564
rect 1876 18508 5068 18564
rect 5124 18508 5134 18564
rect 5282 18508 5292 18564
rect 5348 18508 5740 18564
rect 5796 18508 6076 18564
rect 6132 18508 10108 18564
rect 10164 18508 10174 18564
rect 10546 18508 10556 18564
rect 10612 18508 14476 18564
rect 14532 18508 15036 18564
rect 15092 18508 15102 18564
rect 19058 18508 19068 18564
rect 19124 18508 23212 18564
rect 23268 18508 23278 18564
rect 23426 18508 23436 18564
rect 23492 18508 24444 18564
rect 24500 18508 27580 18564
rect 27636 18508 27646 18564
rect 2594 18396 2604 18452
rect 2660 18396 3388 18452
rect 9426 18396 9436 18452
rect 9492 18396 10444 18452
rect 10500 18396 10510 18452
rect 14354 18396 14364 18452
rect 14420 18396 15708 18452
rect 15764 18396 15774 18452
rect 19282 18396 19292 18452
rect 19348 18396 20188 18452
rect 20244 18396 20748 18452
rect 20804 18396 20814 18452
rect 23538 18396 23548 18452
rect 23604 18396 24108 18452
rect 24164 18396 24174 18452
rect 32162 18396 32172 18452
rect 32228 18396 32844 18452
rect 32900 18396 33516 18452
rect 33572 18396 34524 18452
rect 34580 18396 34590 18452
rect 3332 18340 3388 18396
rect 19292 18340 19348 18396
rect 3332 18284 3948 18340
rect 4004 18284 4014 18340
rect 4834 18284 4844 18340
rect 4900 18284 11004 18340
rect 11060 18284 19348 18340
rect 20132 18284 25228 18340
rect 25284 18284 25294 18340
rect 20132 18228 20188 18284
rect 4274 18172 4284 18228
rect 4340 18172 5964 18228
rect 6020 18172 6030 18228
rect 15250 18172 15260 18228
rect 15316 18172 16156 18228
rect 16212 18172 20188 18228
rect 20290 18172 20300 18228
rect 20356 18172 22652 18228
rect 22708 18172 23884 18228
rect 23940 18172 30492 18228
rect 30548 18172 30558 18228
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 4844 17948 14476 18004
rect 14532 17948 14542 18004
rect 17938 17948 17948 18004
rect 18004 17948 22876 18004
rect 22932 17948 22942 18004
rect 4844 17892 4900 17948
rect 4498 17836 4508 17892
rect 4564 17836 4900 17892
rect 10434 17836 10444 17892
rect 10500 17836 15036 17892
rect 15092 17836 16828 17892
rect 16884 17836 17500 17892
rect 17556 17836 17566 17892
rect 11442 17724 11452 17780
rect 11508 17724 12012 17780
rect 12068 17724 14308 17780
rect 14466 17724 14476 17780
rect 14532 17724 26124 17780
rect 26180 17724 26190 17780
rect 14018 17612 14028 17668
rect 14084 17612 14094 17668
rect 14028 17444 14084 17612
rect 14252 17556 14308 17724
rect 15474 17612 15484 17668
rect 15540 17612 17276 17668
rect 17332 17612 17342 17668
rect 22866 17612 22876 17668
rect 22932 17612 23436 17668
rect 23492 17612 23502 17668
rect 32946 17612 32956 17668
rect 33012 17612 34188 17668
rect 34244 17612 34254 17668
rect 14252 17500 26012 17556
rect 26068 17500 26078 17556
rect 36418 17500 36428 17556
rect 36484 17500 36988 17556
rect 37044 17500 37054 17556
rect 6738 17388 6748 17444
rect 6804 17388 11116 17444
rect 11172 17388 11182 17444
rect 14028 17388 17276 17444
rect 17332 17388 17342 17444
rect 31042 17388 31052 17444
rect 31108 17388 32284 17444
rect 32340 17388 34972 17444
rect 35028 17388 35038 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 30482 17052 30492 17108
rect 30548 17052 30940 17108
rect 30996 17052 31006 17108
rect 31892 17052 32956 17108
rect 33012 17052 33022 17108
rect 5058 16940 5068 16996
rect 5124 16940 6076 16996
rect 6132 16940 9660 16996
rect 9716 16940 9726 16996
rect 31892 16884 31948 17052
rect 35522 16940 35532 16996
rect 35588 16940 35924 16996
rect 6178 16828 6188 16884
rect 6244 16828 11564 16884
rect 11620 16828 11630 16884
rect 17266 16828 17276 16884
rect 17332 16828 18396 16884
rect 18452 16828 20636 16884
rect 20692 16828 20702 16884
rect 29586 16828 29596 16884
rect 29652 16828 31612 16884
rect 31668 16828 31948 16884
rect 35868 16660 35924 16940
rect 35858 16604 35868 16660
rect 35924 16604 35934 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 23090 16268 23100 16324
rect 23156 16268 23436 16324
rect 23492 16268 23996 16324
rect 24052 16268 24062 16324
rect 35634 16268 35644 16324
rect 35700 16268 37436 16324
rect 37492 16268 37502 16324
rect 37314 16156 37324 16212
rect 37380 16156 39564 16212
rect 39620 16156 39630 16212
rect 12898 16044 12908 16100
rect 12964 16044 13804 16100
rect 13860 16044 18956 16100
rect 19012 16044 19022 16100
rect 34402 16044 34412 16100
rect 34468 16044 36092 16100
rect 36148 16044 36158 16100
rect 5842 15932 5852 15988
rect 5908 15932 11004 15988
rect 11060 15932 11900 15988
rect 11956 15932 12572 15988
rect 12628 15932 12638 15988
rect 24994 15932 25004 15988
rect 25060 15932 33852 15988
rect 33908 15932 34300 15988
rect 34356 15932 34366 15988
rect 15698 15820 15708 15876
rect 15764 15820 19964 15876
rect 20020 15820 25340 15876
rect 25396 15820 28700 15876
rect 28756 15820 32508 15876
rect 32564 15820 32574 15876
rect 32722 15820 32732 15876
rect 32788 15820 33180 15876
rect 33236 15820 37100 15876
rect 37156 15820 40348 15876
rect 40404 15820 40414 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 24210 15596 24220 15652
rect 24276 15596 25788 15652
rect 25844 15596 25854 15652
rect 17602 15484 17612 15540
rect 17668 15484 19516 15540
rect 19572 15484 19852 15540
rect 19908 15484 20188 15540
rect 25330 15484 25340 15540
rect 25396 15484 25406 15540
rect 20132 15428 20188 15484
rect 20132 15372 23212 15428
rect 23268 15372 23278 15428
rect 24210 15260 24220 15316
rect 24276 15260 25004 15316
rect 25060 15260 25070 15316
rect 25340 15204 25396 15484
rect 18050 15148 18060 15204
rect 18116 15148 25396 15204
rect 12450 15036 12460 15092
rect 12516 15036 19628 15092
rect 19684 15036 20076 15092
rect 20132 15036 21868 15092
rect 21924 15036 22540 15092
rect 22596 15036 22606 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 24658 14700 24668 14756
rect 24724 14700 25452 14756
rect 25508 14700 25518 14756
rect 23202 14588 23212 14644
rect 23268 14588 24444 14644
rect 24500 14588 25564 14644
rect 25620 14588 29260 14644
rect 29316 14588 29326 14644
rect 30034 14588 30044 14644
rect 30100 14588 31948 14644
rect 32004 14588 32956 14644
rect 33012 14588 33022 14644
rect 20514 14476 20524 14532
rect 20580 14476 22988 14532
rect 23044 14476 23054 14532
rect 15474 14364 15484 14420
rect 15540 14364 15820 14420
rect 15876 14364 15886 14420
rect 4834 14252 4844 14308
rect 4900 14252 6188 14308
rect 6244 14252 10668 14308
rect 10724 14252 10734 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 8530 13916 8540 13972
rect 8596 13916 9996 13972
rect 10052 13916 13692 13972
rect 13748 13916 13758 13972
rect 35410 13916 35420 13972
rect 35476 13916 36540 13972
rect 36596 13916 36606 13972
rect 24546 13804 24556 13860
rect 24612 13804 27244 13860
rect 27300 13804 27310 13860
rect 10210 13692 10220 13748
rect 10276 13692 14364 13748
rect 14420 13692 15036 13748
rect 15092 13692 15102 13748
rect 26562 13692 26572 13748
rect 26628 13692 30044 13748
rect 30100 13692 30110 13748
rect 35634 13692 35644 13748
rect 35700 13692 36316 13748
rect 36372 13692 36382 13748
rect 14130 13580 14140 13636
rect 14196 13580 14924 13636
rect 14980 13580 15596 13636
rect 15652 13580 15662 13636
rect 20402 13580 20412 13636
rect 20468 13580 34748 13636
rect 34804 13580 34814 13636
rect 1922 13468 1932 13524
rect 1988 13468 5180 13524
rect 5236 13468 5964 13524
rect 6020 13468 6030 13524
rect 15362 13468 15372 13524
rect 15428 13468 16044 13524
rect 16100 13468 16110 13524
rect 7298 13356 7308 13412
rect 7364 13356 8428 13412
rect 8484 13356 8494 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 2594 13020 2604 13076
rect 2660 13020 5740 13076
rect 5796 13020 5806 13076
rect 6962 13020 6972 13076
rect 7028 13020 8764 13076
rect 8820 13020 8830 13076
rect 15474 13020 15484 13076
rect 15540 13020 17836 13076
rect 17892 13020 17902 13076
rect 21074 13020 21084 13076
rect 21140 13020 21868 13076
rect 21924 13020 21934 13076
rect 36082 13020 36092 13076
rect 36148 13020 39116 13076
rect 39172 13020 39182 13076
rect 6066 12908 6076 12964
rect 6132 12908 8652 12964
rect 8708 12908 8718 12964
rect 8978 12908 8988 12964
rect 9044 12908 9548 12964
rect 9604 12908 12516 12964
rect 12460 12852 12516 12908
rect 5058 12796 5068 12852
rect 5124 12796 5852 12852
rect 5908 12796 5918 12852
rect 7410 12796 7420 12852
rect 7476 12796 8876 12852
rect 8932 12796 9884 12852
rect 9940 12796 9950 12852
rect 12450 12796 12460 12852
rect 12516 12796 14028 12852
rect 14084 12796 14094 12852
rect 7420 12740 7476 12796
rect 4946 12684 4956 12740
rect 5012 12684 5964 12740
rect 6020 12684 7476 12740
rect 22978 12684 22988 12740
rect 23044 12684 23212 12740
rect 23268 12684 24444 12740
rect 24500 12684 24510 12740
rect 22642 12572 22652 12628
rect 22708 12572 23436 12628
rect 23492 12572 23772 12628
rect 23828 12572 23838 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 6626 12460 6636 12516
rect 6692 12460 10108 12516
rect 10164 12460 11452 12516
rect 11508 12460 13244 12516
rect 13300 12460 13310 12516
rect 9426 12348 9436 12404
rect 9492 12348 9772 12404
rect 9828 12348 9838 12404
rect 10994 12348 11004 12404
rect 11060 12348 13356 12404
rect 13412 12348 13422 12404
rect 20738 12348 20748 12404
rect 20804 12348 22204 12404
rect 22260 12348 23100 12404
rect 23156 12348 23166 12404
rect 23874 12348 23884 12404
rect 23940 12348 24556 12404
rect 24612 12348 24622 12404
rect 7522 12236 7532 12292
rect 7588 12236 8316 12292
rect 8372 12236 9548 12292
rect 9604 12236 9614 12292
rect 24098 12236 24108 12292
rect 24164 12236 24668 12292
rect 24724 12236 25452 12292
rect 25508 12236 25518 12292
rect 5618 12124 5628 12180
rect 5684 12124 6748 12180
rect 6804 12124 6814 12180
rect 9650 12124 9660 12180
rect 9716 12124 10668 12180
rect 10724 12124 10734 12180
rect 21634 12124 21644 12180
rect 21700 12124 22428 12180
rect 22484 12124 23996 12180
rect 24052 12124 24062 12180
rect 9762 12012 9772 12068
rect 9828 12012 11004 12068
rect 11060 12012 11070 12068
rect 21298 11900 21308 11956
rect 21364 11900 22092 11956
rect 22148 11900 22158 11956
rect 36978 11900 36988 11956
rect 37044 11900 39788 11956
rect 39844 11900 39854 11956
rect 5058 11788 5068 11844
rect 5124 11788 5516 11844
rect 5572 11788 6076 11844
rect 6132 11788 6860 11844
rect 6916 11788 6926 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 4834 11676 4844 11732
rect 4900 11676 7308 11732
rect 7364 11676 7374 11732
rect 14354 11452 14364 11508
rect 14420 11452 14924 11508
rect 14980 11452 23212 11508
rect 23268 11452 23278 11508
rect 4386 11340 4396 11396
rect 4452 11340 6748 11396
rect 6804 11340 6814 11396
rect 19618 11340 19628 11396
rect 19684 11340 21756 11396
rect 21812 11340 22652 11396
rect 22708 11340 22718 11396
rect 24658 11340 24668 11396
rect 24724 11340 25340 11396
rect 25396 11340 25406 11396
rect 4162 11228 4172 11284
rect 4228 11228 5964 11284
rect 6020 11228 6030 11284
rect 13906 11228 13916 11284
rect 13972 11228 14140 11284
rect 14196 11228 14206 11284
rect 24210 11228 24220 11284
rect 24276 11228 27356 11284
rect 27412 11228 27422 11284
rect 2594 11116 2604 11172
rect 2660 11116 4284 11172
rect 4340 11116 4350 11172
rect 5842 11116 5852 11172
rect 5908 11116 12012 11172
rect 12068 11116 12078 11172
rect 12898 11116 12908 11172
rect 12964 11116 20412 11172
rect 20468 11116 20478 11172
rect 35186 11116 35196 11172
rect 35252 11116 37660 11172
rect 37716 11116 37996 11172
rect 38052 11116 38062 11172
rect 12908 11060 12964 11116
rect 7074 11004 7084 11060
rect 7140 11004 7644 11060
rect 7700 11004 12964 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 6178 10780 6188 10836
rect 6244 10780 11676 10836
rect 11732 10780 11742 10836
rect 13234 10780 13244 10836
rect 13300 10780 15260 10836
rect 15316 10780 15326 10836
rect 28578 10780 28588 10836
rect 28644 10780 30044 10836
rect 30100 10780 31724 10836
rect 31780 10780 31790 10836
rect 17266 10668 17276 10724
rect 17332 10668 20524 10724
rect 20580 10668 20590 10724
rect 11778 10556 11788 10612
rect 11844 10556 12236 10612
rect 12292 10556 13468 10612
rect 13524 10556 14588 10612
rect 14644 10556 14654 10612
rect 18274 10444 18284 10500
rect 18340 10444 19628 10500
rect 19684 10444 19694 10500
rect 14914 10332 14924 10388
rect 14980 10332 14990 10388
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 12002 10108 12012 10164
rect 12068 10108 12908 10164
rect 12964 10108 12974 10164
rect 14924 10052 14980 10332
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 14924 9996 17836 10052
rect 17892 9996 17902 10052
rect 19618 9996 19628 10052
rect 19684 9996 20412 10052
rect 20468 9996 20478 10052
rect 30146 9996 30156 10052
rect 30212 9996 31388 10052
rect 31444 9996 31454 10052
rect 7746 9884 7756 9940
rect 7812 9884 9436 9940
rect 9492 9884 9502 9940
rect 12114 9884 12124 9940
rect 12180 9884 13804 9940
rect 13860 9884 14028 9940
rect 14084 9884 14094 9940
rect 14924 9716 14980 9996
rect 31042 9884 31052 9940
rect 31108 9884 32060 9940
rect 32116 9884 32126 9940
rect 15810 9772 15820 9828
rect 15876 9772 17500 9828
rect 17556 9772 17566 9828
rect 29922 9772 29932 9828
rect 29988 9772 30604 9828
rect 30660 9772 30670 9828
rect 31826 9772 31836 9828
rect 31892 9772 33964 9828
rect 34020 9772 34524 9828
rect 34580 9772 34590 9828
rect 11554 9660 11564 9716
rect 11620 9660 12348 9716
rect 12404 9660 12414 9716
rect 12562 9660 12572 9716
rect 12628 9660 12796 9716
rect 12852 9660 14980 9716
rect 30818 9660 30828 9716
rect 30884 9660 31948 9716
rect 32004 9660 32116 9716
rect 33730 9660 33740 9716
rect 33796 9660 35644 9716
rect 35700 9660 35710 9716
rect 19282 9548 19292 9604
rect 19348 9548 20300 9604
rect 20356 9548 20366 9604
rect 26450 9548 26460 9604
rect 26516 9548 30604 9604
rect 30660 9548 31388 9604
rect 31444 9548 31454 9604
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 18722 9324 18732 9380
rect 18788 9324 19628 9380
rect 19684 9324 19694 9380
rect 18274 9212 18284 9268
rect 18340 9212 19516 9268
rect 19572 9212 20076 9268
rect 20132 9212 20142 9268
rect 32060 9156 32116 9660
rect 32050 9100 32060 9156
rect 32116 9100 33292 9156
rect 33348 9100 33358 9156
rect 17826 8988 17836 9044
rect 17892 8988 18508 9044
rect 18564 8988 18574 9044
rect 30482 8988 30492 9044
rect 30548 8988 32284 9044
rect 32340 8988 33740 9044
rect 33796 8988 33806 9044
rect 18386 8876 18396 8932
rect 18452 8876 19628 8932
rect 19684 8876 19694 8932
rect 32162 8876 32172 8932
rect 32228 8876 32844 8932
rect 32900 8876 32910 8932
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 34850 8428 34860 8484
rect 34916 8428 36428 8484
rect 36484 8428 36988 8484
rect 37044 8428 38108 8484
rect 38164 8428 38174 8484
rect 20402 8316 20412 8372
rect 20468 8316 21420 8372
rect 21476 8316 25116 8372
rect 25172 8316 25182 8372
rect 18946 8204 18956 8260
rect 19012 8204 19852 8260
rect 19908 8204 19918 8260
rect 20412 8148 20468 8316
rect 14578 8092 14588 8148
rect 14644 8092 18284 8148
rect 18340 8092 18844 8148
rect 18900 8092 19180 8148
rect 19236 8092 19246 8148
rect 20132 8092 20468 8148
rect 20132 8036 20188 8092
rect 5170 7980 5180 8036
rect 5236 7980 7084 8036
rect 7140 7980 10556 8036
rect 10612 7980 10622 8036
rect 17826 7980 17836 8036
rect 17892 7980 20188 8036
rect 23426 7980 23436 8036
rect 23492 7980 23884 8036
rect 23940 7980 25676 8036
rect 25732 7980 25742 8036
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 24546 7644 24556 7700
rect 24612 7644 25340 7700
rect 25396 7644 27804 7700
rect 27860 7644 28364 7700
rect 28420 7644 28430 7700
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 33506 6860 33516 6916
rect 33572 6860 35196 6916
rect 35252 6860 35262 6916
rect 13010 6748 13020 6804
rect 13076 6748 13804 6804
rect 13860 6748 15484 6804
rect 15540 6748 16044 6804
rect 16100 6748 16110 6804
rect 21858 6748 21868 6804
rect 21924 6748 22988 6804
rect 23044 6748 24556 6804
rect 24612 6748 24622 6804
rect 27458 6636 27468 6692
rect 27524 6636 29820 6692
rect 29876 6636 29886 6692
rect 32610 6636 32620 6692
rect 32676 6636 34860 6692
rect 34916 6636 34926 6692
rect 20066 6412 20076 6468
rect 20132 6412 21756 6468
rect 21812 6412 21822 6468
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 17378 6076 17388 6132
rect 17444 6076 19068 6132
rect 19124 6076 20748 6132
rect 20804 6076 20814 6132
rect 28690 5964 28700 6020
rect 28756 5964 30268 6020
rect 30324 5964 30334 6020
rect 29372 5908 29428 5964
rect 10210 5852 10220 5908
rect 10276 5852 10556 5908
rect 10612 5852 13468 5908
rect 13524 5852 13534 5908
rect 29362 5852 29372 5908
rect 29428 5852 29438 5908
rect 29586 5852 29596 5908
rect 29652 5852 30156 5908
rect 30212 5852 30222 5908
rect 18610 5740 18620 5796
rect 18676 5740 20300 5796
rect 20356 5740 20366 5796
rect 25666 5740 25676 5796
rect 25732 5740 26796 5796
rect 26852 5740 26862 5796
rect 27682 5740 27692 5796
rect 27748 5740 28476 5796
rect 28532 5740 28542 5796
rect 29250 5740 29260 5796
rect 29316 5740 31276 5796
rect 31332 5740 31342 5796
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 15250 5068 15260 5124
rect 15316 5068 15932 5124
rect 15988 5068 15998 5124
rect 31938 5068 31948 5124
rect 32004 5068 32620 5124
rect 32676 5068 32686 5124
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 12450 4284 12460 4340
rect 12516 4284 15708 4340
rect 15764 4284 17388 4340
rect 17444 4284 17454 4340
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 39452 37996 39508 38052
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 39452 36540 39508 36596
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 8764 28588 8820 28644
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 8764 24780 8820 24836
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 41580 4768 42396
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 19808 42364 20128 42396
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 8764 28644 8820 28654
rect 8764 24836 8820 28588
rect 8764 24770 8820 24780
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 41580 35488 42396
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 39452 38052 39508 38062
rect 39452 36596 39508 37996
rect 39452 36530 39508 36540
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _337_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 25312 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _338_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 29568 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _339_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _340_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25424 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _341_
timestamp 1698431365
transform -1 0 26656 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _342_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25648 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _343_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27664 0 -1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _344_
timestamp 1698431365
transform -1 0 29680 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _345_
timestamp 1698431365
transform -1 0 28672 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _346_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20496 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _347_
timestamp 1698431365
transform -1 0 18816 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _348_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19376 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _349_
timestamp 1698431365
transform -1 0 22176 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _350_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19488 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _351_
timestamp 1698431365
transform -1 0 14672 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _352_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7504 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _353_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11312 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _354_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16240 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _355_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7168 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _356_
timestamp 1698431365
transform 1 0 9632 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _357_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13104 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _358_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29680 0 1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _359_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32144 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _360_
timestamp 1698431365
transform -1 0 38192 0 -1 15680
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _361_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30800 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _362_
timestamp 1698431365
transform 1 0 15680 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _363_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14224 0 1 25088
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _364_
timestamp 1698431365
transform 1 0 15792 0 1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _365_
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _366_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10528 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _367_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8288 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _368_
timestamp 1698431365
transform 1 0 6272 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _369_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9520 0 -1 21952
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _370_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16912 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _371_
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _372_
timestamp 1698431365
transform -1 0 14224 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _373_
timestamp 1698431365
transform -1 0 11088 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _374_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10080 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _375_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10640 0 -1 23520
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _376_
timestamp 1698431365
transform -1 0 10304 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _377_
timestamp 1698431365
transform 1 0 9632 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _378_
timestamp 1698431365
transform -1 0 9184 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _379_
timestamp 1698431365
transform 1 0 9856 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _380_
timestamp 1698431365
transform 1 0 15008 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _381_
timestamp 1698431365
transform 1 0 14896 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _382_
timestamp 1698431365
transform -1 0 10416 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _383_
timestamp 1698431365
transform 1 0 14448 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _384_
timestamp 1698431365
transform 1 0 9520 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _385_
timestamp 1698431365
transform -1 0 5824 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _386_
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _387_
timestamp 1698431365
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _388_
timestamp 1698431365
transform 1 0 7168 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _389_
timestamp 1698431365
transform 1 0 8064 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _390_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _391_
timestamp 1698431365
transform 1 0 15008 0 1 23520
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _392_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _393_
timestamp 1698431365
transform 1 0 9744 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _394_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12208 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _395_
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _396_
timestamp 1698431365
transform 1 0 14896 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _397_
timestamp 1698431365
transform 1 0 6832 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _398_
timestamp 1698431365
transform 1 0 13776 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _399_
timestamp 1698431365
transform 1 0 10080 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _400_
timestamp 1698431365
transform -1 0 16912 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _401_
timestamp 1698431365
transform -1 0 20272 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _402_
timestamp 1698431365
transform -1 0 19712 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _403_
timestamp 1698431365
transform 1 0 14336 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _404_
timestamp 1698431365
transform 1 0 11536 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _405_
timestamp 1698431365
transform -1 0 18592 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _406_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15232 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _407_
timestamp 1698431365
transform 1 0 12880 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _408_
timestamp 1698431365
transform 1 0 14448 0 1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _409_
timestamp 1698431365
transform -1 0 12880 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _410_
timestamp 1698431365
transform -1 0 12320 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _411_
timestamp 1698431365
transform 1 0 19824 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _412_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10864 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _413_
timestamp 1698431365
transform -1 0 10864 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _414_
timestamp 1698431365
transform 1 0 14224 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _415_
timestamp 1698431365
transform 1 0 13664 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _416_
timestamp 1698431365
transform -1 0 11872 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _417_
timestamp 1698431365
transform 1 0 11984 0 -1 37632
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _418_
timestamp 1698431365
transform -1 0 12768 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _419_
timestamp 1698431365
transform 1 0 15344 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _420_
timestamp 1698431365
transform 1 0 16688 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _421_
timestamp 1698431365
transform 1 0 13888 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _422_
timestamp 1698431365
transform 1 0 15792 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _423_
timestamp 1698431365
transform 1 0 15232 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _424_
timestamp 1698431365
transform 1 0 16464 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _425_
timestamp 1698431365
transform 1 0 14896 0 1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _426_
timestamp 1698431365
transform -1 0 11424 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _427_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8512 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _428_
timestamp 1698431365
transform 1 0 24080 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _429_
timestamp 1698431365
transform 1 0 25312 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _430_
timestamp 1698431365
transform 1 0 34160 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _431_
timestamp 1698431365
transform -1 0 25984 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _432_
timestamp 1698431365
transform -1 0 32592 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _433_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30912 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _434_
timestamp 1698431365
transform -1 0 32144 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _435_
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _436_
timestamp 1698431365
transform -1 0 22736 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _437_
timestamp 1698431365
transform -1 0 20944 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _438_
timestamp 1698431365
transform 1 0 31696 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _439_
timestamp 1698431365
transform -1 0 31248 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _440_
timestamp 1698431365
transform 1 0 30912 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _441_
timestamp 1698431365
transform -1 0 36064 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _442_
timestamp 1698431365
transform 1 0 35056 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _443_
timestamp 1698431365
transform 1 0 24752 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _444_
timestamp 1698431365
transform 1 0 34720 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _445_
timestamp 1698431365
transform -1 0 34720 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _446_
timestamp 1698431365
transform 1 0 35728 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _447_
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _448_
timestamp 1698431365
transform -1 0 36736 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _449_
timestamp 1698431365
transform -1 0 21056 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _450_
timestamp 1698431365
transform -1 0 35840 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _451_
timestamp 1698431365
transform 1 0 35728 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _452_
timestamp 1698431365
transform -1 0 35280 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _453_
timestamp 1698431365
transform -1 0 34272 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _454_
timestamp 1698431365
transform -1 0 35616 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _455_
timestamp 1698431365
transform 1 0 35280 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _456_
timestamp 1698431365
transform -1 0 32592 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _457_
timestamp 1698431365
transform 1 0 25648 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _458_
timestamp 1698431365
transform -1 0 32480 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _459_
timestamp 1698431365
transform -1 0 33824 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _460_
timestamp 1698431365
transform 1 0 30352 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _461_
timestamp 1698431365
transform -1 0 32368 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _462_
timestamp 1698431365
transform -1 0 30352 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _463_
timestamp 1698431365
transform 1 0 29904 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _464_
timestamp 1698431365
transform 1 0 29008 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _465_
timestamp 1698431365
transform -1 0 26880 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _466_
timestamp 1698431365
transform -1 0 29008 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _467_
timestamp 1698431365
transform -1 0 28000 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _468_
timestamp 1698431365
transform -1 0 25872 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _469_
timestamp 1698431365
transform 1 0 32144 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _470_
timestamp 1698431365
transform 1 0 23968 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _471_
timestamp 1698431365
transform 1 0 23968 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _472_
timestamp 1698431365
transform 1 0 33936 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _473_
timestamp 1698431365
transform 1 0 34944 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _474_
timestamp 1698431365
transform -1 0 29904 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _475_
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _476_
timestamp 1698431365
transform 1 0 36960 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _477_
timestamp 1698431365
transform 1 0 36400 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _478_
timestamp 1698431365
transform 1 0 34272 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _479_
timestamp 1698431365
transform 1 0 33040 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _480_
timestamp 1698431365
transform 1 0 35280 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _481_
timestamp 1698431365
transform -1 0 34944 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _482_
timestamp 1698431365
transform 1 0 36960 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _483_
timestamp 1698431365
transform 1 0 39312 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _484_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 34272 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _485_
timestamp 1698431365
transform -1 0 42896 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _486_
timestamp 1698431365
transform -1 0 37744 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _487_
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _488_
timestamp 1698431365
transform 1 0 32032 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _489_
timestamp 1698431365
transform 1 0 40656 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _490_
timestamp 1698431365
transform 1 0 39424 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _491_
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _492_
timestamp 1698431365
transform 1 0 28896 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _493_
timestamp 1698431365
transform 1 0 29344 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _494_
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _495_
timestamp 1698431365
transform -1 0 41888 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _496_
timestamp 1698431365
transform 1 0 40096 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _497_
timestamp 1698431365
transform 1 0 40544 0 1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _498_
timestamp 1698431365
transform -1 0 41440 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _499_
timestamp 1698431365
transform -1 0 39760 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _500_
timestamp 1698431365
transform -1 0 40096 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _501_
timestamp 1698431365
transform 1 0 37184 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _502_
timestamp 1698431365
transform -1 0 39424 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _503_
timestamp 1698431365
transform 1 0 28672 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _504_
timestamp 1698431365
transform 1 0 34496 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _505_
timestamp 1698431365
transform -1 0 34496 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _506_
timestamp 1698431365
transform -1 0 33936 0 1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _507_
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _508_
timestamp 1698431365
transform -1 0 37856 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _509_
timestamp 1698431365
transform -1 0 34272 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _510_
timestamp 1698431365
transform -1 0 42896 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _511_
timestamp 1698431365
transform 1 0 36176 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _512_
timestamp 1698431365
transform 1 0 38528 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _513_
timestamp 1698431365
transform -1 0 39536 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _514_
timestamp 1698431365
transform 1 0 40320 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _515_
timestamp 1698431365
transform -1 0 41664 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _516_
timestamp 1698431365
transform 1 0 26208 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _517_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42000 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _518_
timestamp 1698431365
transform -1 0 42896 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _519_
timestamp 1698431365
transform -1 0 40880 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _520_
timestamp 1698431365
transform -1 0 41664 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _521_
timestamp 1698431365
transform 1 0 39200 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _522_
timestamp 1698431365
transform 1 0 40656 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _523_
timestamp 1698431365
transform -1 0 42000 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _524_
timestamp 1698431365
transform -1 0 36064 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _525_
timestamp 1698431365
transform 1 0 34720 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _526_
timestamp 1698431365
transform 1 0 38080 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _527_
timestamp 1698431365
transform 1 0 36624 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _528_
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _529_
timestamp 1698431365
transform -1 0 35616 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _530_
timestamp 1698431365
transform -1 0 33824 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _531_
timestamp 1698431365
transform 1 0 37072 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _532_
timestamp 1698431365
transform 1 0 35168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _533_
timestamp 1698431365
transform 1 0 20048 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _534_
timestamp 1698431365
transform 1 0 10528 0 -1 26656
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _535_
timestamp 1698431365
transform 1 0 12208 0 -1 25088
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _536_
timestamp 1698431365
transform -1 0 16240 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _537_
timestamp 1698431365
transform -1 0 20608 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _538_
timestamp 1698431365
transform 1 0 20608 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _539_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15680 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _540_
timestamp 1698431365
transform -1 0 17584 0 1 21952
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _541_
timestamp 1698431365
transform -1 0 19824 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _542_
timestamp 1698431365
transform 1 0 19152 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _543_
timestamp 1698431365
transform 1 0 19600 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _544_
timestamp 1698431365
transform 1 0 18928 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _545_
timestamp 1698431365
transform -1 0 6384 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _546_
timestamp 1698431365
transform -1 0 23072 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _547_
timestamp 1698431365
transform -1 0 12208 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _548_
timestamp 1698431365
transform 1 0 18704 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _549_
timestamp 1698431365
transform -1 0 13104 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _550_
timestamp 1698431365
transform 1 0 4480 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _551_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _552_
timestamp 1698431365
transform -1 0 4480 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _553_
timestamp 1698431365
transform -1 0 11760 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _554_
timestamp 1698431365
transform -1 0 10640 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _555_
timestamp 1698431365
transform -1 0 11200 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _556_
timestamp 1698431365
transform 1 0 10416 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _557_
timestamp 1698431365
transform 1 0 10864 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _558_
timestamp 1698431365
transform 1 0 19376 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _559_
timestamp 1698431365
transform -1 0 17808 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _560_
timestamp 1698431365
transform -1 0 14000 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _561_
timestamp 1698431365
transform -1 0 14672 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _562_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15904 0 -1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _563_
timestamp 1698431365
transform 1 0 4592 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _564_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10640 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _565_
timestamp 1698431365
transform -1 0 5824 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _566_
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _567_
timestamp 1698431365
transform 1 0 6496 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _568_
timestamp 1698431365
transform -1 0 4592 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _569_
timestamp 1698431365
transform -1 0 6384 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _570_
timestamp 1698431365
transform 1 0 4816 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _571_
timestamp 1698431365
transform 1 0 11984 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _572_
timestamp 1698431365
transform 1 0 6832 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _573_
timestamp 1698431365
transform 1 0 8176 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _574_
timestamp 1698431365
transform -1 0 24640 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _575_
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _576_
timestamp 1698431365
transform 1 0 8064 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _577_
timestamp 1698431365
transform -1 0 10416 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _578_
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _579_
timestamp 1698431365
transform 1 0 14112 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _580_
timestamp 1698431365
transform -1 0 14560 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _581_
timestamp 1698431365
transform 1 0 14560 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _582_
timestamp 1698431365
transform -1 0 14000 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _583_
timestamp 1698431365
transform -1 0 15568 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _584_
timestamp 1698431365
transform -1 0 12992 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _585_
timestamp 1698431365
transform -1 0 12432 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _586_
timestamp 1698431365
transform -1 0 12656 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _587_
timestamp 1698431365
transform -1 0 11760 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _588_
timestamp 1698431365
transform -1 0 15344 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _589_
timestamp 1698431365
transform -1 0 15232 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _590_
timestamp 1698431365
transform -1 0 15008 0 -1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _591_
timestamp 1698431365
transform -1 0 23744 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _592_
timestamp 1698431365
transform -1 0 14672 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _593_
timestamp 1698431365
transform -1 0 14224 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _594_
timestamp 1698431365
transform -1 0 18816 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _595_
timestamp 1698431365
transform 1 0 13664 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _596_
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _597_
timestamp 1698431365
transform -1 0 19936 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _598_
timestamp 1698431365
transform 1 0 18256 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _599_
timestamp 1698431365
transform -1 0 18592 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _600_
timestamp 1698431365
transform -1 0 25984 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _601_
timestamp 1698431365
transform -1 0 18256 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _602_
timestamp 1698431365
transform 1 0 19488 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _603_
timestamp 1698431365
transform -1 0 20608 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _604_
timestamp 1698431365
transform -1 0 19376 0 1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _605_
timestamp 1698431365
transform 1 0 19712 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _606_
timestamp 1698431365
transform 1 0 15120 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _607_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18480 0 1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _608_
timestamp 1698431365
transform 1 0 20272 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _609_
timestamp 1698431365
transform -1 0 23968 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _610_
timestamp 1698431365
transform 1 0 21952 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _611_
timestamp 1698431365
transform 1 0 20944 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _612_
timestamp 1698431365
transform -1 0 22848 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _613_
timestamp 1698431365
transform 1 0 22960 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _614_
timestamp 1698431365
transform -1 0 25984 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _615_
timestamp 1698431365
transform 1 0 23856 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _616_
timestamp 1698431365
transform -1 0 24864 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _617_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22848 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _618_
timestamp 1698431365
transform 1 0 23968 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _619_
timestamp 1698431365
transform -1 0 25760 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _620_
timestamp 1698431365
transform 1 0 23408 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _621_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24640 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _622_
timestamp 1698431365
transform 1 0 23184 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _623_
timestamp 1698431365
transform 1 0 23072 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _624_
timestamp 1698431365
transform 1 0 23632 0 -1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _625_
timestamp 1698431365
transform -1 0 24640 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _626_
timestamp 1698431365
transform 1 0 23072 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _627_
timestamp 1698431365
transform 1 0 22848 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _628_
timestamp 1698431365
transform 1 0 23632 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _629_
timestamp 1698431365
transform 1 0 23856 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _630_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19712 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _631_
timestamp 1698431365
transform -1 0 9296 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _632_
timestamp 1698431365
transform 1 0 10192 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _633_
timestamp 1698431365
transform -1 0 8624 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _634_
timestamp 1698431365
transform -1 0 9184 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _635_
timestamp 1698431365
transform -1 0 8512 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _636_
timestamp 1698431365
transform -1 0 6160 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _637_
timestamp 1698431365
transform -1 0 6832 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _638_
timestamp 1698431365
transform 1 0 10304 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _639_
timestamp 1698431365
transform -1 0 6720 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _640_
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _641_
timestamp 1698431365
transform -1 0 5600 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _642_
timestamp 1698431365
transform 1 0 3584 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _643_
timestamp 1698431365
transform -1 0 3920 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _644_
timestamp 1698431365
transform -1 0 9184 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _645_
timestamp 1698431365
transform -1 0 4928 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _646_
timestamp 1698431365
transform 1 0 3920 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _647_
timestamp 1698431365
transform -1 0 5376 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _648_
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _649_
timestamp 1698431365
transform 1 0 8512 0 1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _650_
timestamp 1698431365
transform -1 0 15904 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _651_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12320 0 1 28224
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _652_
timestamp 1698431365
transform -1 0 4032 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _653_
timestamp 1698431365
transform -1 0 19264 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _654_
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _655_
timestamp 1698431365
transform 1 0 19264 0 -1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _656_
timestamp 1698431365
transform 1 0 15904 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _657_
timestamp 1698431365
transform 1 0 15904 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _658_
timestamp 1698431365
transform 1 0 17024 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _659_
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _660_
timestamp 1698431365
transform -1 0 16128 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _661_
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _662_
timestamp 1698431365
transform -1 0 19376 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _663_
timestamp 1698431365
transform 1 0 20384 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _664_
timestamp 1698431365
transform 1 0 27440 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _665_
timestamp 1698431365
transform 1 0 29008 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _666_
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _667_
timestamp 1698431365
transform 1 0 24640 0 1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _668_
timestamp 1698431365
transform -1 0 24752 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _669_
timestamp 1698431365
transform -1 0 24640 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _670_
timestamp 1698431365
transform 1 0 24192 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _671_
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _672_
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _673_
timestamp 1698431365
transform 1 0 27328 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _674_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17696 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _675_
timestamp 1698431365
transform 1 0 2016 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _676_
timestamp 1698431365
transform 1 0 20160 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _677_
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _678_
timestamp 1698431365
transform 1 0 28336 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _679_
timestamp 1698431365
transform 1 0 30688 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _680_
timestamp 1698431365
transform 1 0 5936 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _681_
timestamp 1698431365
transform -1 0 36624 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _682_
timestamp 1698431365
transform 1 0 29232 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _683_
timestamp 1698431365
transform -1 0 32704 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _684_
timestamp 1698431365
transform -1 0 40544 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _685_
timestamp 1698431365
transform -1 0 40096 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _686_
timestamp 1698431365
transform 1 0 34608 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _687_
timestamp 1698431365
transform -1 0 36176 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _688_
timestamp 1698431365
transform 1 0 28224 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _689_
timestamp 1698431365
transform -1 0 32256 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _690_
timestamp 1698431365
transform 1 0 24304 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _691_
timestamp 1698431365
transform 1 0 6272 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _692_
timestamp 1698431365
transform 1 0 2800 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _693_
timestamp 1698431365
transform 1 0 1792 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _694_
timestamp 1698431365
transform -1 0 35056 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _695_
timestamp 1698431365
transform -1 0 31808 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _696_
timestamp 1698431365
transform -1 0 37744 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _697_
timestamp 1698431365
transform 1 0 40880 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _698_
timestamp 1698431365
transform 1 0 40992 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _699_
timestamp 1698431365
transform 1 0 40992 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _700_
timestamp 1698431365
transform 1 0 37744 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _701_
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _702_
timestamp 1698431365
transform 1 0 30128 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _703_
timestamp 1698431365
transform -1 0 40544 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _704_
timestamp 1698431365
transform 1 0 40992 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _705_
timestamp 1698431365
transform 1 0 40992 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _706_
timestamp 1698431365
transform 1 0 40544 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _707_
timestamp 1698431365
transform 1 0 36176 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _708_
timestamp 1698431365
transform 1 0 30800 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _709_
timestamp 1698431365
transform 1 0 33824 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _710_
timestamp 1698431365
transform -1 0 20944 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _711_
timestamp 1698431365
transform 1 0 1680 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _712_
timestamp 1698431365
transform 1 0 5824 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _713_
timestamp 1698431365
transform 1 0 13776 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _714_
timestamp 1698431365
transform 1 0 1680 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _715_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1680 0 1 14112
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _716_
timestamp 1698431365
transform 1 0 6832 0 1 7840
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _717_
timestamp 1698431365
transform -1 0 18816 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _718_
timestamp 1698431365
transform 1 0 9968 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _719_
timestamp 1698431365
transform 1 0 12208 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _720_
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _721_
timestamp 1698431365
transform -1 0 22736 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _722_
timestamp 1698431365
transform 1 0 21616 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _723_
timestamp 1698431365
transform -1 0 28336 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _724_
timestamp 1698431365
transform 1 0 26320 0 -1 14112
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _725_
timestamp 1698431365
transform 1 0 24528 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _726_
timestamp 1698431365
transform -1 0 9744 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _727_
timestamp 1698431365
transform 1 0 2016 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _728_
timestamp 1698431365
transform 1 0 2016 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _729_
timestamp 1698431365
transform 1 0 2464 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _730_
timestamp 1698431365
transform 1 0 2240 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _731_
timestamp 1698431365
transform -1 0 21728 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _732_
timestamp 1698431365
transform -1 0 16576 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _733_
timestamp 1698431365
transform 1 0 20048 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _734_
timestamp 1698431365
transform -1 0 30464 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _735_
timestamp 1698431365
transform 1 0 22512 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _736_
timestamp 1698431365
transform 1 0 22624 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _737_
timestamp 1698431365
transform 1 0 26544 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__362__I $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15456 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__363__B
timestamp 1698431365
transform 1 0 18144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__395__A1
timestamp 1698431365
transform 1 0 11984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__408__A1
timestamp 1698431365
transform 1 0 15456 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__411__I
timestamp 1698431365
transform 1 0 19600 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__412__B
timestamp 1698431365
transform -1 0 12544 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__417__C
timestamp 1698431365
transform 1 0 16688 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__428__I
timestamp 1698431365
transform 1 0 23408 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__430__A2
timestamp 1698431365
transform 1 0 33936 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__433__A1
timestamp 1698431365
transform 1 0 29792 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__435__I
timestamp 1698431365
transform 1 0 20720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__436__I
timestamp 1698431365
transform 1 0 21840 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__439__A1
timestamp 1698431365
transform 1 0 30464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__443__I
timestamp 1698431365
transform 1 0 23856 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__445__A1
timestamp 1698431365
transform 1 0 33824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__450__B
timestamp 1698431365
transform 1 0 34720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__454__B
timestamp 1698431365
transform 1 0 34496 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__I
timestamp 1698431365
transform 1 0 25424 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__B
timestamp 1698431365
transform 1 0 31360 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__462__A1
timestamp 1698431365
transform -1 0 29456 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__463__B
timestamp 1698431365
transform -1 0 31248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__465__I
timestamp 1698431365
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__468__A1
timestamp 1698431365
transform -1 0 26320 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__470__I
timestamp 1698431365
transform 1 0 24864 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__474__I
timestamp 1698431365
transform -1 0 30352 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__475__I
timestamp 1698431365
transform -1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__476__I
timestamp 1698431365
transform 1 0 36736 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__477__A1
timestamp 1698431365
transform 1 0 36176 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__480__I
timestamp 1698431365
transform 1 0 35056 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__482__I
timestamp 1698431365
transform 1 0 36400 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__484__A2
timestamp 1698431365
transform -1 0 34496 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__484__C
timestamp 1698431365
transform 1 0 35392 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__490__C
timestamp 1698431365
transform 1 0 40544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__494__I
timestamp 1698431365
transform 1 0 29904 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__495__A2
timestamp 1698431365
transform 1 0 42112 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__497__A1
timestamp 1698431365
transform -1 0 40544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__502__C
timestamp 1698431365
transform 1 0 39984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__506__A1
timestamp 1698431365
transform 1 0 32928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__509__B
timestamp 1698431365
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__511__I
timestamp 1698431365
transform 1 0 35952 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__514__A1
timestamp 1698431365
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__515__A1
timestamp 1698431365
transform 1 0 40320 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__517__A2
timestamp 1698431365
transform 1 0 39984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__517__C
timestamp 1698431365
transform 1 0 40432 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__520__A2
timestamp 1698431365
transform 1 0 40320 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__521__A1
timestamp 1698431365
transform -1 0 39200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__522__A1
timestamp 1698431365
transform 1 0 39984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__523__A2
timestamp 1698431365
transform 1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__523__C
timestamp 1698431365
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__524__I
timestamp 1698431365
transform -1 0 35616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__527__A1
timestamp 1698431365
transform -1 0 36624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__530__B
timestamp 1698431365
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__532__A2
timestamp 1698431365
transform 1 0 34944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__537__A1
timestamp 1698431365
transform 1 0 21504 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__539__B
timestamp 1698431365
transform -1 0 14224 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__540__B
timestamp 1698431365
transform -1 0 15456 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__542__I
timestamp 1698431365
transform 1 0 18928 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__547__I
timestamp 1698431365
transform 1 0 12432 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__552__A1
timestamp 1698431365
transform 1 0 4480 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__557__B
timestamp 1698431365
transform 1 0 11984 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__558__I
timestamp 1698431365
transform 1 0 20048 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__562__C
timestamp 1698431365
transform 1 0 16128 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__567__B
timestamp 1698431365
transform 1 0 7616 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__571__I
timestamp 1698431365
transform 1 0 12880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__575__C
timestamp 1698431365
transform 1 0 6608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__578__C
timestamp 1698431365
transform 1 0 11424 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__581__C
timestamp 1698431365
transform 1 0 16016 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__586__B
timestamp 1698431365
transform 1 0 12880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__591__A1
timestamp 1698431365
transform 1 0 22624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__592__B2
timestamp 1698431365
transform 1 0 14896 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__593__C
timestamp 1698431365
transform 1 0 15232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__597__B
timestamp 1698431365
transform 1 0 18256 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__600__I
timestamp 1698431365
transform 1 0 26208 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__601__B
timestamp 1698431365
transform 1 0 17808 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__603__A2
timestamp 1698431365
transform 1 0 19712 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__605__B
timestamp 1698431365
transform 1 0 21392 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__610__B
timestamp 1698431365
transform 1 0 21728 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__611__A1
timestamp 1698431365
transform 1 0 21840 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__613__A1
timestamp 1698431365
transform 1 0 23856 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__617__A3
timestamp 1698431365
transform 1 0 24416 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__618__B
timestamp 1698431365
transform 1 0 25312 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__622__A1
timestamp 1698431365
transform 1 0 22960 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__624__C
timestamp 1698431365
transform -1 0 25088 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__626__A1
timestamp 1698431365
transform 1 0 22848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__628__A1
timestamp 1698431365
transform 1 0 22624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__632__B
timestamp 1698431365
transform -1 0 11536 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__635__A1
timestamp 1698431365
transform -1 0 7952 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__638__I
timestamp 1698431365
transform 1 0 10640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__639__A2
timestamp 1698431365
transform 1 0 6944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__640__B
timestamp 1698431365
transform -1 0 6832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__643__C
timestamp 1698431365
transform 1 0 3584 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__647__B
timestamp 1698431365
transform 1 0 6048 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__648__A3
timestamp 1698431365
transform 1 0 10864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__651__C
timestamp 1698431365
transform 1 0 12544 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__655__A1
timestamp 1698431365
transform 1 0 20272 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__656__A2
timestamp 1698431365
transform 1 0 17248 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__659__C
timestamp 1698431365
transform 1 0 18368 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__663__A1
timestamp 1698431365
transform -1 0 20384 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__664__A2
timestamp 1698431365
transform 1 0 28336 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__665__A1
timestamp 1698431365
transform 1 0 28784 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__668__A1
timestamp 1698431365
transform 1 0 23968 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__671__A1
timestamp 1698431365
transform 1 0 25984 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__672__A1
timestamp 1698431365
transform 1 0 28896 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__672__B
timestamp 1698431365
transform 1 0 30128 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__673__A1
timestamp 1698431365
transform 1 0 28448 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__673__C
timestamp 1698431365
transform 1 0 27104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__674__CLK
timestamp 1698431365
transform 1 0 21392 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__675__CLK
timestamp 1698431365
transform -1 0 5712 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__676__CLK
timestamp 1698431365
transform -1 0 20160 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__677__CLK
timestamp 1698431365
transform 1 0 28336 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__678__CLK
timestamp 1698431365
transform -1 0 32032 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__679__CLK
timestamp 1698431365
transform 1 0 34160 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__680__CLK
timestamp 1698431365
transform -1 0 9856 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__681__CLK
timestamp 1698431365
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__682__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__683__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__684__CLK
timestamp 1698431365
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__685__CLK
timestamp 1698431365
transform 1 0 36624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__686__CLK
timestamp 1698431365
transform 1 0 38080 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__687__CLK
timestamp 1698431365
transform 1 0 36400 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__688__CLK
timestamp 1698431365
transform 1 0 31696 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__689__CLK
timestamp 1698431365
transform -1 0 32704 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__690__CLK
timestamp 1698431365
transform 1 0 27776 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__691__CLK
timestamp 1698431365
transform 1 0 9744 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__692__CLK
timestamp 1698431365
transform 1 0 6272 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__693__CLK
timestamp 1698431365
transform 1 0 5712 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__694__CLK
timestamp 1698431365
transform 1 0 35280 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__695__CLK
timestamp 1698431365
transform 1 0 32032 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__696__CLK
timestamp 1698431365
transform -1 0 38192 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__697__CLK
timestamp 1698431365
transform -1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__698__CLK
timestamp 1698431365
transform 1 0 40320 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__699__CLK
timestamp 1698431365
transform 1 0 40768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__700__CLK
timestamp 1698431365
transform 1 0 37520 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__701__CLK
timestamp 1698431365
transform 1 0 36400 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__702__CLK
timestamp 1698431365
transform 1 0 33600 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__703__CLK
timestamp 1698431365
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__704__CLK
timestamp 1698431365
transform 1 0 40320 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__705__CLK
timestamp 1698431365
transform -1 0 39984 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__706__CLK
timestamp 1698431365
transform 1 0 40320 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__707__CLK
timestamp 1698431365
transform -1 0 39872 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__708__CLK
timestamp 1698431365
transform 1 0 34272 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__709__CLK
timestamp 1698431365
transform -1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__710__CLK
timestamp 1698431365
transform 1 0 21392 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__711__CLK
timestamp 1698431365
transform 1 0 4928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__712__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__713__CLK
timestamp 1698431365
transform 1 0 17248 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__714__CLK
timestamp 1698431365
transform 1 0 5152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__715__CLK
timestamp 1698431365
transform 1 0 5152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__716__CLK
timestamp 1698431365
transform 1 0 10528 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__717__CLK
timestamp 1698431365
transform 1 0 19040 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__718__CLK
timestamp 1698431365
transform 1 0 13440 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__719__CLK
timestamp 1698431365
transform 1 0 15680 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__720__CLK
timestamp 1698431365
transform 1 0 20720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__721__CLK
timestamp 1698431365
transform 1 0 22960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__722__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__723__CLK
timestamp 1698431365
transform 1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__724__CLK
timestamp 1698431365
transform 1 0 30016 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__725__CLK
timestamp 1698431365
transform 1 0 28000 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__726__CLK
timestamp 1698431365
transform 1 0 9968 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__727__CLK
timestamp 1698431365
transform -1 0 5936 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__728__CLK
timestamp 1698431365
transform 1 0 5712 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__729__CLK
timestamp 1698431365
transform 1 0 5936 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__730__CLK
timestamp 1698431365
transform -1 0 5936 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__731__CLK
timestamp 1698431365
transform 1 0 18256 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__732__CLK
timestamp 1698431365
transform 1 0 16800 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__733__CLK
timestamp 1698431365
transform 1 0 19824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__734__CLK
timestamp 1698431365
transform 1 0 30688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__735__CLK
timestamp 1698431365
transform 1 0 25984 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__736__CLK
timestamp 1698431365
transform 1 0 26096 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__737__CLK
timestamp 1698431365
transform 1 0 30016 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 21616 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_0__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 15680 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_1__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 19936 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_2__f_wb_clk_i_I
timestamp 1698431365
transform -1 0 16576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_3__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 20272 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_4__f_wb_clk_i_I
timestamp 1698431365
transform -1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_5__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 32480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_6__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 29904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_7__f_wb_clk_i_I
timestamp 1698431365
transform -1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 5152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output10_I
timestamp 1698431365
transform 1 0 39760 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21616 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1698431365
transform -1 0 15456 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1698431365
transform 1 0 14112 0 1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1698431365
transform -1 0 15680 0 -1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1698431365
transform 1 0 14448 0 1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1698431365
transform 1 0 29232 0 1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1698431365
transform 1 0 33040 0 -1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_376 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_72 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_88
timestamp 1698431365
transform 1 0 11200 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_96 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12096 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_126 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15456 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_130
timestamp 1698431365
transform 1 0 15904 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_138
timestamp 1698431365
transform 1 0 16800 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_158
timestamp 1698431365
transform 1 0 19040 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_191
timestamp 1698431365
transform 1 0 22736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_195
timestamp 1698431365
transform 1 0 23184 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_203
timestamp 1698431365
transform 1 0 24080 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698431365
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698431365
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698431365
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_346
timestamp 1698431365
transform 1 0 40096 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_123
timestamp 1698431365
transform 1 0 15120 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_127
timestamp 1698431365
transform 1 0 15568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_166
timestamp 1698431365
transform 1 0 19936 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_174
timestamp 1698431365
transform 1 0 20832 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_193
timestamp 1698431365
transform 1 0 22960 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_201
timestamp 1698431365
transform 1 0 23856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_234
timestamp 1698431365
transform 1 0 27552 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_238
timestamp 1698431365
transform 1 0 28000 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_242
timestamp 1698431365
transform 1 0 28448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_244
timestamp 1698431365
transform 1 0 28672 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_276
timestamp 1698431365
transform 1 0 32256 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_280
timestamp 1698431365
transform 1 0 32704 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_312
timestamp 1698431365
transform 1 0 36288 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_314
timestamp 1698431365
transform 1 0 36512 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_381
timestamp 1698431365
transform 1 0 44016 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_383
timestamp 1698431365
transform 1 0 44240 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_76
timestamp 1698431365
transform 1 0 9856 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_106
timestamp 1698431365
transform 1 0 13216 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_110
timestamp 1698431365
transform 1 0 13664 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_126
timestamp 1698431365
transform 1 0 15456 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_134
timestamp 1698431365
transform 1 0 16352 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_138
timestamp 1698431365
transform 1 0 16800 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_171
timestamp 1698431365
transform 1 0 20496 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_175
timestamp 1698431365
transform 1 0 20944 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_207
timestamp 1698431365
transform 1 0 24528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_209
timestamp 1698431365
transform 1 0 24752 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_219
timestamp 1698431365
transform 1 0 25872 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_223
timestamp 1698431365
transform 1 0 26320 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_225
timestamp 1698431365
transform 1 0 26544 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_238
timestamp 1698431365
transform 1 0 28000 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_263
timestamp 1698431365
transform 1 0 30800 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_267
timestamp 1698431365
transform 1 0 31248 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_275
timestamp 1698431365
transform 1 0 32144 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_279
timestamp 1698431365
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_311
timestamp 1698431365
transform 1 0 36176 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_315
timestamp 1698431365
transform 1 0 36624 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_347
timestamp 1698431365
transform 1 0 40208 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_349
timestamp 1698431365
transform 1 0 40432 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_115
timestamp 1698431365
transform 1 0 14224 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_125
timestamp 1698431365
transform 1 0 15344 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_141
timestamp 1698431365
transform 1 0 17136 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_149
timestamp 1698431365
transform 1 0 18032 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_156
timestamp 1698431365
transform 1 0 18816 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_172
timestamp 1698431365
transform 1 0 20608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698431365
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_251
timestamp 1698431365
transform 1 0 29456 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_290
timestamp 1698431365
transform 1 0 33824 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_306
timestamp 1698431365
transform 1 0 35616 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_314
timestamp 1698431365
transform 1 0 36512 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_381
timestamp 1698431365
transform 1 0 44016 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_383
timestamp 1698431365
transform 1 0 44240 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_174
timestamp 1698431365
transform 1 0 20832 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_178
timestamp 1698431365
transform 1 0 21280 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_180
timestamp 1698431365
transform 1 0 21504 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_216
timestamp 1698431365
transform 1 0 25536 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_248
timestamp 1698431365
transform 1 0 29120 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_264
timestamp 1698431365
transform 1 0 30912 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_272
timestamp 1698431365
transform 1 0 31808 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_279
timestamp 1698431365
transform 1 0 32592 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_45
timestamp 1698431365
transform 1 0 6384 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_80
timestamp 1698431365
transform 1 0 10304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_84
timestamp 1698431365
transform 1 0 10752 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_100
timestamp 1698431365
transform 1 0 12544 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_104
timestamp 1698431365
transform 1 0 12992 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_113
timestamp 1698431365
transform 1 0 14000 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_121
timestamp 1698431365
transform 1 0 14896 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_131
timestamp 1698431365
transform 1 0 16016 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_161
timestamp 1698431365
transform 1 0 19376 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_163
timestamp 1698431365
transform 1 0 19600 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_172
timestamp 1698431365
transform 1 0 20608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1698431365
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_181
timestamp 1698431365
transform 1 0 21616 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_189
timestamp 1698431365
transform 1 0 22512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_199
timestamp 1698431365
transform 1 0 23632 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_203
timestamp 1698431365
transform 1 0 24080 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_235
timestamp 1698431365
transform 1 0 27664 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_243
timestamp 1698431365
transform 1 0 28560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_381
timestamp 1698431365
transform 1 0 44016 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_383
timestamp 1698431365
transform 1 0 44240 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_88
timestamp 1698431365
transform 1 0 11200 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_96
timestamp 1698431365
transform 1 0 12096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_98
timestamp 1698431365
transform 1 0 12320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_104
timestamp 1698431365
transform 1 0 12992 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_159
timestamp 1698431365
transform 1 0 19152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_161
timestamp 1698431365
transform 1 0 19376 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_170
timestamp 1698431365
transform 1 0 20384 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_202
timestamp 1698431365
transform 1 0 23968 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_244
timestamp 1698431365
transform 1 0 28672 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_260
timestamp 1698431365
transform 1 0 30464 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_278
timestamp 1698431365
transform 1 0 32480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_290
timestamp 1698431365
transform 1 0 33824 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_294
timestamp 1698431365
transform 1 0 34272 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_296
timestamp 1698431365
transform 1 0 34496 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_326
timestamp 1698431365
transform 1 0 37856 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_330
timestamp 1698431365
transform 1 0 38304 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_346
timestamp 1698431365
transform 1 0 40096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_69
timestamp 1698431365
transform 1 0 9072 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_85
timestamp 1698431365
transform 1 0 10864 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_109
timestamp 1698431365
transform 1 0 13552 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_124
timestamp 1698431365
transform 1 0 15232 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_140
timestamp 1698431365
transform 1 0 17024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_172
timestamp 1698431365
transform 1 0 20608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_174
timestamp 1698431365
transform 1 0 20832 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698431365
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_277
timestamp 1698431365
transform 1 0 32368 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_285
timestamp 1698431365
transform 1 0 33264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_287
timestamp 1698431365
transform 1 0 33488 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_294
timestamp 1698431365
transform 1 0 34272 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_310
timestamp 1698431365
transform 1 0 36064 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_314
timestamp 1698431365
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_381
timestamp 1698431365
transform 1 0 44016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_383
timestamp 1698431365
transform 1 0 44240 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_32
timestamp 1698431365
transform 1 0 4928 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_36
timestamp 1698431365
transform 1 0 5376 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_68
timestamp 1698431365
transform 1 0 8960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_88
timestamp 1698431365
transform 1 0 11200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_99
timestamp 1698431365
transform 1 0 12432 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_103
timestamp 1698431365
transform 1 0 12880 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_122
timestamp 1698431365
transform 1 0 15008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_126
timestamp 1698431365
transform 1 0 15456 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_134
timestamp 1698431365
transform 1 0 16352 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_138
timestamp 1698431365
transform 1 0 16800 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_150
timestamp 1698431365
transform 1 0 18144 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_153
timestamp 1698431365
transform 1 0 18480 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_161
timestamp 1698431365
transform 1 0 19376 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_163
timestamp 1698431365
transform 1 0 19600 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_166
timestamp 1698431365
transform 1 0 19936 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_198
timestamp 1698431365
transform 1 0 23520 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698431365
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_216
timestamp 1698431365
transform 1 0 25536 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_232
timestamp 1698431365
transform 1 0 27328 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_269
timestamp 1698431365
transform 1 0 31472 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_273
timestamp 1698431365
transform 1 0 31920 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_277
timestamp 1698431365
transform 1 0 32368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_279
timestamp 1698431365
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_290
timestamp 1698431365
transform 1 0 33824 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_294
timestamp 1698431365
transform 1 0 34272 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_309
timestamp 1698431365
transform 1 0 35952 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_341
timestamp 1698431365
transform 1 0 39536 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_349
timestamp 1698431365
transform 1 0 40432 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_18
timestamp 1698431365
transform 1 0 3360 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_22
timestamp 1698431365
transform 1 0 3808 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_54
timestamp 1698431365
transform 1 0 7392 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_58
timestamp 1698431365
transform 1 0 7840 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_90
timestamp 1698431365
transform 1 0 11424 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_98
timestamp 1698431365
transform 1 0 12320 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_102
timestamp 1698431365
transform 1 0 12768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_104
timestamp 1698431365
transform 1 0 12992 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_109
timestamp 1698431365
transform 1 0 13552 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_119
timestamp 1698431365
transform 1 0 14672 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_123
timestamp 1698431365
transform 1 0 15120 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_155
timestamp 1698431365
transform 1 0 18704 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698431365
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_181
timestamp 1698431365
transform 1 0 21616 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_192
timestamp 1698431365
transform 1 0 22848 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_210
timestamp 1698431365
transform 1 0 24864 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_241
timestamp 1698431365
transform 1 0 28336 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_279
timestamp 1698431365
transform 1 0 32592 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_295
timestamp 1698431365
transform 1 0 34384 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_306
timestamp 1698431365
transform 1 0 35616 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_314
timestamp 1698431365
transform 1 0 36512 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_381
timestamp 1698431365
transform 1 0 44016 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_383
timestamp 1698431365
transform 1 0 44240 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_34
timestamp 1698431365
transform 1 0 5152 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_40
timestamp 1698431365
transform 1 0 5824 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_44
timestamp 1698431365
transform 1 0 6272 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_46
timestamp 1698431365
transform 1 0 6496 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_49
timestamp 1698431365
transform 1 0 6832 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_57
timestamp 1698431365
transform 1 0 7728 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_88
timestamp 1698431365
transform 1 0 11200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_92
timestamp 1698431365
transform 1 0 11648 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_124
timestamp 1698431365
transform 1 0 15232 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_158
timestamp 1698431365
transform 1 0 19040 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_166
timestamp 1698431365
transform 1 0 19936 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_168
timestamp 1698431365
transform 1 0 20160 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698431365
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_314
timestamp 1698431365
transform 1 0 36512 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_317
timestamp 1698431365
transform 1 0 36848 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_349
timestamp 1698431365
transform 1 0 40432 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_18
timestamp 1698431365
transform 1 0 3360 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_26
timestamp 1698431365
transform 1 0 4256 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_30
timestamp 1698431365
transform 1 0 4704 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_47
timestamp 1698431365
transform 1 0 6608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_56
timestamp 1698431365
transform 1 0 7616 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_92
timestamp 1698431365
transform 1 0 11648 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_94
timestamp 1698431365
transform 1 0 11872 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_115
timestamp 1698431365
transform 1 0 14224 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_156
timestamp 1698431365
transform 1 0 18816 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_160
timestamp 1698431365
transform 1 0 19264 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_168
timestamp 1698431365
transform 1 0 20160 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_172
timestamp 1698431365
transform 1 0 20608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698431365
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_181
timestamp 1698431365
transform 1 0 21616 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_185
timestamp 1698431365
transform 1 0 22064 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_193
timestamp 1698431365
transform 1 0 22960 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_204
timestamp 1698431365
transform 1 0 24192 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_208
timestamp 1698431365
transform 1 0 24640 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_212
timestamp 1698431365
transform 1 0 25088 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_220
timestamp 1698431365
transform 1 0 25984 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_236
timestamp 1698431365
transform 1 0 27776 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698431365
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_279
timestamp 1698431365
transform 1 0 32592 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_295
timestamp 1698431365
transform 1 0 34384 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_303
timestamp 1698431365
transform 1 0 35280 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_313
timestamp 1698431365
transform 1 0 36400 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_346
timestamp 1698431365
transform 1 0 40096 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_378
timestamp 1698431365
transform 1 0 43680 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_382
timestamp 1698431365
transform 1 0 44128 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_36
timestamp 1698431365
transform 1 0 5376 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_68
timestamp 1698431365
transform 1 0 8960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_81
timestamp 1698431365
transform 1 0 10416 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_89
timestamp 1698431365
transform 1 0 11312 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_97
timestamp 1698431365
transform 1 0 12208 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_101
timestamp 1698431365
transform 1 0 12656 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_109
timestamp 1698431365
transform 1 0 13552 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_129
timestamp 1698431365
transform 1 0 15792 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_133
timestamp 1698431365
transform 1 0 16240 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_137
timestamp 1698431365
transform 1 0 16688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698431365
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698431365
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_220
timestamp 1698431365
transform 1 0 25984 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_222
timestamp 1698431365
transform 1 0 26208 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_254
timestamp 1698431365
transform 1 0 29792 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_258
timestamp 1698431365
transform 1 0 30240 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_274
timestamp 1698431365
transform 1 0 32032 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_278
timestamp 1698431365
transform 1 0 32480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_316
timestamp 1698431365
transform 1 0 36736 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_348
timestamp 1698431365
transform 1 0 40320 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_45
timestamp 1698431365
transform 1 0 6384 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_77
timestamp 1698431365
transform 1 0 9968 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_93
timestamp 1698431365
transform 1 0 11760 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698431365
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_111
timestamp 1698431365
transform 1 0 13776 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_113
timestamp 1698431365
transform 1 0 14000 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_119
timestamp 1698431365
transform 1 0 14672 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_121
timestamp 1698431365
transform 1 0 14896 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_128
timestamp 1698431365
transform 1 0 15680 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_160
timestamp 1698431365
transform 1 0 19264 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_164
timestamp 1698431365
transform 1 0 19712 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_166
timestamp 1698431365
transform 1 0 19936 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_169
timestamp 1698431365
transform 1 0 20272 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698431365
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_185
timestamp 1698431365
transform 1 0 22064 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_189
timestamp 1698431365
transform 1 0 22512 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_191
timestamp 1698431365
transform 1 0 22736 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_208
timestamp 1698431365
transform 1 0 24640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_212
timestamp 1698431365
transform 1 0 25088 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_218
timestamp 1698431365
transform 1 0 25760 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_234
timestamp 1698431365
transform 1 0 27552 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_242
timestamp 1698431365
transform 1 0 28448 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_297
timestamp 1698431365
transform 1 0 34608 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_313
timestamp 1698431365
transform 1 0 36400 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_381
timestamp 1698431365
transform 1 0 44016 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_383
timestamp 1698431365
transform 1 0 44240 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698431365
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698431365
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_158
timestamp 1698431365
transform 1 0 19040 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_160
timestamp 1698431365
transform 1 0 19264 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_167
timestamp 1698431365
transform 1 0 20048 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_176
timestamp 1698431365
transform 1 0 21056 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_192
timestamp 1698431365
transform 1 0 22848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_249
timestamp 1698431365
transform 1 0 29232 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_286
timestamp 1698431365
transform 1 0 33376 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_290
timestamp 1698431365
transform 1 0 33824 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_329
timestamp 1698431365
transform 1 0 38192 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_345
timestamp 1698431365
transform 1 0 39984 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_349
timestamp 1698431365
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_69
timestamp 1698431365
transform 1 0 9072 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_93
timestamp 1698431365
transform 1 0 11760 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_97
timestamp 1698431365
transform 1 0 12208 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_113
timestamp 1698431365
transform 1 0 14000 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_164
timestamp 1698431365
transform 1 0 19712 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_168
timestamp 1698431365
transform 1 0 20160 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698431365
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_200
timestamp 1698431365
transform 1 0 23744 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_232
timestamp 1698431365
transform 1 0 27328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_240
timestamp 1698431365
transform 1 0 28224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698431365
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_263
timestamp 1698431365
transform 1 0 30800 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_270
timestamp 1698431365
transform 1 0 31584 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_286
timestamp 1698431365
transform 1 0 33376 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_304
timestamp 1698431365
transform 1 0 35392 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_306
timestamp 1698431365
transform 1 0 35616 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_350
timestamp 1698431365
transform 1 0 40544 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_382
timestamp 1698431365
transform 1 0 44128 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_34
timestamp 1698431365
transform 1 0 5152 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_38
timestamp 1698431365
transform 1 0 5600 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_69
timestamp 1698431365
transform 1 0 9072 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_126
timestamp 1698431365
transform 1 0 15456 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_130
timestamp 1698431365
transform 1 0 15904 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698431365
transform 1 0 16800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_147
timestamp 1698431365
transform 1 0 17808 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_163
timestamp 1698431365
transform 1 0 19600 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_175
timestamp 1698431365
transform 1 0 20944 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698431365
transform 1 0 24528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698431365
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_244
timestamp 1698431365
transform 1 0 28672 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_267
timestamp 1698431365
transform 1 0 31248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_275
timestamp 1698431365
transform 1 0 32144 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_277
timestamp 1698431365
transform 1 0 32368 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_332
timestamp 1698431365
transform 1 0 38528 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_348
timestamp 1698431365
transform 1 0 40320 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_18
timestamp 1698431365
transform 1 0 3360 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_26
timestamp 1698431365
transform 1 0 4256 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_30
timestamp 1698431365
transform 1 0 4704 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_46
timestamp 1698431365
transform 1 0 6496 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_62
timestamp 1698431365
transform 1 0 8288 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_83
timestamp 1698431365
transform 1 0 10640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_93
timestamp 1698431365
transform 1 0 11760 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_97
timestamp 1698431365
transform 1 0 12208 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_140
timestamp 1698431365
transform 1 0 17024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_144
timestamp 1698431365
transform 1 0 17472 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_160
timestamp 1698431365
transform 1 0 19264 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_168
timestamp 1698431365
transform 1 0 20160 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_172
timestamp 1698431365
transform 1 0 20608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698431365
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_185
timestamp 1698431365
transform 1 0 22064 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_189
timestamp 1698431365
transform 1 0 22512 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_191
timestamp 1698431365
transform 1 0 22736 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_202
timestamp 1698431365
transform 1 0 23968 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_208
timestamp 1698431365
transform 1 0 24640 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_240
timestamp 1698431365
transform 1 0 28224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698431365
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_263
timestamp 1698431365
transform 1 0 30800 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_284
timestamp 1698431365
transform 1 0 33152 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_300
timestamp 1698431365
transform 1 0 34944 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_310
timestamp 1698431365
transform 1 0 36064 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_314
timestamp 1698431365
transform 1 0 36512 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_323
timestamp 1698431365
transform 1 0 37520 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_355
timestamp 1698431365
transform 1 0 41104 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_371
timestamp 1698431365
transform 1 0 42896 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_379
timestamp 1698431365
transform 1 0 43792 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_383
timestamp 1698431365
transform 1 0 44240 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_18
timestamp 1698431365
transform 1 0 3360 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_40
timestamp 1698431365
transform 1 0 5824 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_56
timestamp 1698431365
transform 1 0 7616 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_64
timestamp 1698431365
transform 1 0 8512 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698431365
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_74
timestamp 1698431365
transform 1 0 9632 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_88
timestamp 1698431365
transform 1 0 11200 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_104
timestamp 1698431365
transform 1 0 12992 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_108
timestamp 1698431365
transform 1 0 13440 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_110
timestamp 1698431365
transform 1 0 13664 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_130
timestamp 1698431365
transform 1 0 15904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_134
timestamp 1698431365
transform 1 0 16352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1698431365
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_150
timestamp 1698431365
transform 1 0 18144 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_154
timestamp 1698431365
transform 1 0 18592 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_156
timestamp 1698431365
transform 1 0 18816 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_175
timestamp 1698431365
transform 1 0 20944 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_183
timestamp 1698431365
transform 1 0 21840 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_187
timestamp 1698431365
transform 1 0 22288 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_189
timestamp 1698431365
transform 1 0 22512 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_244
timestamp 1698431365
transform 1 0 28672 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_260
timestamp 1698431365
transform 1 0 30464 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_268
timestamp 1698431365
transform 1 0 31360 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_270
timestamp 1698431365
transform 1 0 31584 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_290
timestamp 1698431365
transform 1 0 33824 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_299
timestamp 1698431365
transform 1 0 34832 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_331
timestamp 1698431365
transform 1 0 38416 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_347
timestamp 1698431365
transform 1 0 40208 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_349
timestamp 1698431365
transform 1 0 40432 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698431365
transform 1 0 4928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_45
timestamp 1698431365
transform 1 0 6384 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_61
timestamp 1698431365
transform 1 0 8176 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_69
timestamp 1698431365
transform 1 0 9072 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_73
timestamp 1698431365
transform 1 0 9520 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_78
timestamp 1698431365
transform 1 0 10080 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_94
timestamp 1698431365
transform 1 0 11872 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_102
timestamp 1698431365
transform 1 0 12768 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698431365
transform 1 0 12992 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_115
timestamp 1698431365
transform 1 0 14224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_119
timestamp 1698431365
transform 1 0 14672 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_125
timestamp 1698431365
transform 1 0 15344 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_141
timestamp 1698431365
transform 1 0 17136 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_145
timestamp 1698431365
transform 1 0 17584 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_181
timestamp 1698431365
transform 1 0 21616 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_197
timestamp 1698431365
transform 1 0 23408 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_236
timestamp 1698431365
transform 1 0 27776 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_240
timestamp 1698431365
transform 1 0 28224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698431365
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_251
timestamp 1698431365
transform 1 0 29456 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_253
timestamp 1698431365
transform 1 0 29680 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_264
timestamp 1698431365
transform 1 0 30912 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_275
timestamp 1698431365
transform 1 0 32144 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_283
timestamp 1698431365
transform 1 0 33040 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_285
timestamp 1698431365
transform 1 0 33264 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_321
timestamp 1698431365
transform 1 0 37296 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_353
timestamp 1698431365
transform 1 0 40880 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_369
timestamp 1698431365
transform 1 0 42672 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_377
timestamp 1698431365
transform 1 0 43568 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_381
timestamp 1698431365
transform 1 0 44016 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_383
timestamp 1698431365
transform 1 0 44240 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_18
timestamp 1698431365
transform 1 0 3360 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_26
timestamp 1698431365
transform 1 0 4256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_30
timestamp 1698431365
transform 1 0 4704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_34
timestamp 1698431365
transform 1 0 5152 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_50
timestamp 1698431365
transform 1 0 6944 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_58
timestamp 1698431365
transform 1 0 7840 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_74
timestamp 1698431365
transform 1 0 9632 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_87
timestamp 1698431365
transform 1 0 11088 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_103
timestamp 1698431365
transform 1 0 12880 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_111
timestamp 1698431365
transform 1 0 13776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_115
timestamp 1698431365
transform 1 0 14224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_133
timestamp 1698431365
transform 1 0 16240 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_137
timestamp 1698431365
transform 1 0 16688 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698431365
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_158
timestamp 1698431365
transform 1 0 19040 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_162
timestamp 1698431365
transform 1 0 19488 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_171
timestamp 1698431365
transform 1 0 20496 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_203
timestamp 1698431365
transform 1 0 24080 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_207
timestamp 1698431365
transform 1 0 24528 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_244
timestamp 1698431365
transform 1 0 28672 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_248
timestamp 1698431365
transform 1 0 29120 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698431365
transform 1 0 32480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_286
timestamp 1698431365
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_53
timestamp 1698431365
transform 1 0 7280 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_57
timestamp 1698431365
transform 1 0 7728 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_59
timestamp 1698431365
transform 1 0 7952 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_92
timestamp 1698431365
transform 1 0 11648 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_100
timestamp 1698431365
transform 1 0 12544 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698431365
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_152
timestamp 1698431365
transform 1 0 18368 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_168
timestamp 1698431365
transform 1 0 20160 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_172
timestamp 1698431365
transform 1 0 20608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_209
timestamp 1698431365
transform 1 0 24752 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_211
timestamp 1698431365
transform 1 0 24976 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_220
timestamp 1698431365
transform 1 0 25984 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_224
timestamp 1698431365
transform 1 0 26432 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_240
timestamp 1698431365
transform 1 0 28224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_251
timestamp 1698431365
transform 1 0 29456 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_263
timestamp 1698431365
transform 1 0 30800 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_295
timestamp 1698431365
transform 1 0 34384 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_333
timestamp 1698431365
transform 1 0 38640 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_341
timestamp 1698431365
transform 1 0 39536 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_345
timestamp 1698431365
transform 1 0 39984 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_347
timestamp 1698431365
transform 1 0 40208 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_379
timestamp 1698431365
transform 1 0 43792 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_383
timestamp 1698431365
transform 1 0 44240 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_34
timestamp 1698431365
transform 1 0 5152 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_42
timestamp 1698431365
transform 1 0 6048 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_56
timestamp 1698431365
transform 1 0 7616 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_64
timestamp 1698431365
transform 1 0 8512 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698431365
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_113
timestamp 1698431365
transform 1 0 14000 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_121
timestamp 1698431365
transform 1 0 14896 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_123
timestamp 1698431365
transform 1 0 15120 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_126
timestamp 1698431365
transform 1 0 15456 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_134
timestamp 1698431365
transform 1 0 16352 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_138
timestamp 1698431365
transform 1 0 16800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_150
timestamp 1698431365
transform 1 0 18144 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_154
timestamp 1698431365
transform 1 0 18592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_161
timestamp 1698431365
transform 1 0 19376 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_193
timestamp 1698431365
transform 1 0 22960 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_201
timestamp 1698431365
transform 1 0 23856 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_205
timestamp 1698431365
transform 1 0 24304 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_207
timestamp 1698431365
transform 1 0 24528 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_228
timestamp 1698431365
transform 1 0 26880 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_244
timestamp 1698431365
transform 1 0 28672 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_259
timestamp 1698431365
transform 1 0 30352 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_275
timestamp 1698431365
transform 1 0 32144 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698431365
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_298
timestamp 1698431365
transform 1 0 34720 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_306
timestamp 1698431365
transform 1 0 35616 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_310
timestamp 1698431365
transform 1 0 36064 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_340
timestamp 1698431365
transform 1 0 39424 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_344
timestamp 1698431365
transform 1 0 39872 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_348
timestamp 1698431365
transform 1 0 40320 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_360
timestamp 1698431365
transform 1 0 41664 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_364
timestamp 1698431365
transform 1 0 42112 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_366
timestamp 1698431365
transform 1 0 42336 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_371
timestamp 1698431365
transform 1 0 42896 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_379
timestamp 1698431365
transform 1 0 43792 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_383
timestamp 1698431365
transform 1 0 44240 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698431365
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_123
timestamp 1698431365
transform 1 0 15120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_125
timestamp 1698431365
transform 1 0 15344 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_145
timestamp 1698431365
transform 1 0 17584 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_153
timestamp 1698431365
transform 1 0 18480 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_165
timestamp 1698431365
transform 1 0 19824 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_173
timestamp 1698431365
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_231
timestamp 1698431365
transform 1 0 27216 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_239
timestamp 1698431365
transform 1 0 28112 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_243
timestamp 1698431365
transform 1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698431365
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_333
timestamp 1698431365
transform 1 0 38640 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_341
timestamp 1698431365
transform 1 0 39536 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_347
timestamp 1698431365
transform 1 0 40208 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_357
timestamp 1698431365
transform 1 0 41328 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_373
timestamp 1698431365
transform 1 0 43120 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_381
timestamp 1698431365
transform 1 0 44016 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_383
timestamp 1698431365
transform 1 0 44240 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_6
timestamp 1698431365
transform 1 0 2016 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_37
timestamp 1698431365
transform 1 0 5488 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_41
timestamp 1698431365
transform 1 0 5936 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_57
timestamp 1698431365
transform 1 0 7728 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_65
timestamp 1698431365
transform 1 0 8624 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_80
timestamp 1698431365
transform 1 0 10304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_82
timestamp 1698431365
transform 1 0 10528 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_126
timestamp 1698431365
transform 1 0 15456 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_133
timestamp 1698431365
transform 1 0 16240 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698431365
transform 1 0 16688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698431365
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_150
timestamp 1698431365
transform 1 0 18144 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_154
timestamp 1698431365
transform 1 0 18592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_178
timestamp 1698431365
transform 1 0 21280 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_182
timestamp 1698431365
transform 1 0 21728 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_208
timestamp 1698431365
transform 1 0 24640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_228
timestamp 1698431365
transform 1 0 26880 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_258
timestamp 1698431365
transform 1 0 30240 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_274
timestamp 1698431365
transform 1 0 32032 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698431365
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_287
timestamp 1698431365
transform 1 0 33488 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_295
timestamp 1698431365
transform 1 0 34384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_297
timestamp 1698431365
transform 1 0 34608 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_310
timestamp 1698431365
transform 1 0 36064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_312
timestamp 1698431365
transform 1 0 36288 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_323
timestamp 1698431365
transform 1 0 37520 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_331
timestamp 1698431365
transform 1 0 38416 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_335
timestamp 1698431365
transform 1 0 38864 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_363
timestamp 1698431365
transform 1 0 42000 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_379
timestamp 1698431365
transform 1 0 43792 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_383
timestamp 1698431365
transform 1 0 44240 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_41
timestamp 1698431365
transform 1 0 5936 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_43
timestamp 1698431365
transform 1 0 6160 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_56
timestamp 1698431365
transform 1 0 7616 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_72
timestamp 1698431365
transform 1 0 9408 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_76
timestamp 1698431365
transform 1 0 9856 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_94
timestamp 1698431365
transform 1 0 11872 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_102
timestamp 1698431365
transform 1 0 12768 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_104
timestamp 1698431365
transform 1 0 12992 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_115
timestamp 1698431365
transform 1 0 14224 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_119
timestamp 1698431365
transform 1 0 14672 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_121
timestamp 1698431365
transform 1 0 14896 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_165
timestamp 1698431365
transform 1 0 19824 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_173
timestamp 1698431365
transform 1 0 20720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_185
timestamp 1698431365
transform 1 0 22064 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_194
timestamp 1698431365
transform 1 0 23072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_196
timestamp 1698431365
transform 1 0 23296 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_199
timestamp 1698431365
transform 1 0 23632 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_215
timestamp 1698431365
transform 1 0 25424 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_231
timestamp 1698431365
transform 1 0 27216 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_239
timestamp 1698431365
transform 1 0 28112 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698431365
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_253
timestamp 1698431365
transform 1 0 29680 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_257
timestamp 1698431365
transform 1 0 30128 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_261
timestamp 1698431365
transform 1 0 30576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_292
timestamp 1698431365
transform 1 0 34048 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_296
timestamp 1698431365
transform 1 0 34496 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_310
timestamp 1698431365
transform 1 0 36064 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698431365
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_349
timestamp 1698431365
transform 1 0 40432 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_353
timestamp 1698431365
transform 1 0 40880 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_369
timestamp 1698431365
transform 1 0 42672 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_377
timestamp 1698431365
transform 1 0 43568 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_381
timestamp 1698431365
transform 1 0 44016 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_383
timestamp 1698431365
transform 1 0 44240 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_34
timestamp 1698431365
transform 1 0 5152 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_50
timestamp 1698431365
transform 1 0 6944 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_54
timestamp 1698431365
transform 1 0 7392 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_63
timestamp 1698431365
transform 1 0 8400 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_67
timestamp 1698431365
transform 1 0 8848 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_69
timestamp 1698431365
transform 1 0 9072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_88
timestamp 1698431365
transform 1 0 11200 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_96
timestamp 1698431365
transform 1 0 12096 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_134
timestamp 1698431365
transform 1 0 16352 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698431365
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_150
timestamp 1698431365
transform 1 0 18144 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_154
timestamp 1698431365
transform 1 0 18592 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_156
timestamp 1698431365
transform 1 0 18816 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_159
timestamp 1698431365
transform 1 0 19152 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_191
timestamp 1698431365
transform 1 0 22736 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_207
timestamp 1698431365
transform 1 0 24528 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698431365
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_228
timestamp 1698431365
transform 1 0 26880 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_236
timestamp 1698431365
transform 1 0 27776 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_240
timestamp 1698431365
transform 1 0 28224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_244
timestamp 1698431365
transform 1 0 28672 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_248
timestamp 1698431365
transform 1 0 29120 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_264
timestamp 1698431365
transform 1 0 30912 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_272
timestamp 1698431365
transform 1 0 31808 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_276
timestamp 1698431365
transform 1 0 32256 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_290
timestamp 1698431365
transform 1 0 33824 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_322
timestamp 1698431365
transform 1 0 37408 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_326
timestamp 1698431365
transform 1 0 37856 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_336
timestamp 1698431365
transform 1 0 38976 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_344
timestamp 1698431365
transform 1 0 39872 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_360
timestamp 1698431365
transform 1 0 41664 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_376
timestamp 1698431365
transform 1 0 43456 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_45
timestamp 1698431365
transform 1 0 6384 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_49
timestamp 1698431365
transform 1 0 6832 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_57
timestamp 1698431365
transform 1 0 7728 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_61
timestamp 1698431365
transform 1 0 8176 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_63
timestamp 1698431365
transform 1 0 8400 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_70
timestamp 1698431365
transform 1 0 9184 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_86
timestamp 1698431365
transform 1 0 10976 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_90
timestamp 1698431365
transform 1 0 11424 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_92
timestamp 1698431365
transform 1 0 11648 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_148
timestamp 1698431365
transform 1 0 17920 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_152
timestamp 1698431365
transform 1 0 18368 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_168
timestamp 1698431365
transform 1 0 20160 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698431365
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698431365
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_193
timestamp 1698431365
transform 1 0 22960 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_201
timestamp 1698431365
transform 1 0 23856 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_208
timestamp 1698431365
transform 1 0 24640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_212
timestamp 1698431365
transform 1 0 25088 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_228
timestamp 1698431365
transform 1 0 26880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698431365
transform 1 0 28448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698431365
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_255
timestamp 1698431365
transform 1 0 29904 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_259
timestamp 1698431365
transform 1 0 30352 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_291
timestamp 1698431365
transform 1 0 33936 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_299
timestamp 1698431365
transform 1 0 34832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_310
timestamp 1698431365
transform 1 0 36064 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698431365
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_321
timestamp 1698431365
transform 1 0 37296 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_337
timestamp 1698431365
transform 1 0 39088 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_341
timestamp 1698431365
transform 1 0 39536 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_353
timestamp 1698431365
transform 1 0 40880 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_383
timestamp 1698431365
transform 1 0 44240 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_18
timestamp 1698431365
transform 1 0 3360 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_24
timestamp 1698431365
transform 1 0 4032 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_40
timestamp 1698431365
transform 1 0 5824 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_49
timestamp 1698431365
transform 1 0 6832 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_65
timestamp 1698431365
transform 1 0 8624 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_69
timestamp 1698431365
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_80
timestamp 1698431365
transform 1 0 10304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_119
timestamp 1698431365
transform 1 0 14672 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_133
timestamp 1698431365
transform 1 0 16240 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_137
timestamp 1698431365
transform 1 0 16688 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698431365
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_161
timestamp 1698431365
transform 1 0 19376 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_196
timestamp 1698431365
transform 1 0 23296 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_204
timestamp 1698431365
transform 1 0 24192 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698431365
transform 1 0 24640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_220
timestamp 1698431365
transform 1 0 25984 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_224
timestamp 1698431365
transform 1 0 26432 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_254
timestamp 1698431365
transform 1 0 29792 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_258
timestamp 1698431365
transform 1 0 30240 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_274
timestamp 1698431365
transform 1 0 32032 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_278
timestamp 1698431365
transform 1 0 32480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_327
timestamp 1698431365
transform 1 0 37968 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_343
timestamp 1698431365
transform 1 0 39760 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_345
timestamp 1698431365
transform 1 0 39984 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_348
timestamp 1698431365
transform 1 0 40320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698431365
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_111
timestamp 1698431365
transform 1 0 13776 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_134
timestamp 1698431365
transform 1 0 16352 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_138
timestamp 1698431365
transform 1 0 16800 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_148
timestamp 1698431365
transform 1 0 17920 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_164
timestamp 1698431365
transform 1 0 19712 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_191
timestamp 1698431365
transform 1 0 22736 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_207
timestamp 1698431365
transform 1 0 24528 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_225
timestamp 1698431365
transform 1 0 26544 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698431365
transform 1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_255
timestamp 1698431365
transform 1 0 29904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_259
timestamp 1698431365
transform 1 0 30352 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_291
timestamp 1698431365
transform 1 0 33936 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_299
timestamp 1698431365
transform 1 0 34832 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_306
timestamp 1698431365
transform 1 0 35616 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_310
timestamp 1698431365
transform 1 0 36064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_312
timestamp 1698431365
transform 1 0 36288 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_324
timestamp 1698431365
transform 1 0 37632 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_332
timestamp 1698431365
transform 1 0 38528 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_336
timestamp 1698431365
transform 1 0 38976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_338
timestamp 1698431365
transform 1 0 39200 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_347
timestamp 1698431365
transform 1 0 40208 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_360
timestamp 1698431365
transform 1 0 41664 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_376
timestamp 1698431365
transform 1 0 43456 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_18
timestamp 1698431365
transform 1 0 3360 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_38
timestamp 1698431365
transform 1 0 5600 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_83
timestamp 1698431365
transform 1 0 10640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_87
timestamp 1698431365
transform 1 0 11088 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_119
timestamp 1698431365
transform 1 0 14672 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_123
timestamp 1698431365
transform 1 0 15120 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_125
timestamp 1698431365
transform 1 0 15344 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_128
timestamp 1698431365
transform 1 0 15680 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698431365
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_151
timestamp 1698431365
transform 1 0 18256 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_185
timestamp 1698431365
transform 1 0 22064 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_201
timestamp 1698431365
transform 1 0 23856 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698431365
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698431365
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_286
timestamp 1698431365
transform 1 0 33376 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_290
timestamp 1698431365
transform 1 0 33824 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_322
timestamp 1698431365
transform 1 0 37408 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_338
timestamp 1698431365
transform 1 0 39200 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698431365
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_360
timestamp 1698431365
transform 1 0 41664 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_376
timestamp 1698431365
transform 1 0 43456 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_10
timestamp 1698431365
transform 1 0 2464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_12
timestamp 1698431365
transform 1 0 2688 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_48
timestamp 1698431365
transform 1 0 6720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_52
timestamp 1698431365
transform 1 0 7168 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_56
timestamp 1698431365
transform 1 0 7616 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_98
timestamp 1698431365
transform 1 0 12320 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_102
timestamp 1698431365
transform 1 0 12768 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_104
timestamp 1698431365
transform 1 0 12992 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_115
timestamp 1698431365
transform 1 0 14224 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_123
timestamp 1698431365
transform 1 0 15120 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_127
timestamp 1698431365
transform 1 0 15568 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_129
timestamp 1698431365
transform 1 0 15792 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_140
timestamp 1698431365
transform 1 0 17024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_144
timestamp 1698431365
transform 1 0 17472 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_154
timestamp 1698431365
transform 1 0 18592 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_170
timestamp 1698431365
transform 1 0 20384 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_185
timestamp 1698431365
transform 1 0 22064 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_189
timestamp 1698431365
transform 1 0 22512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_219
timestamp 1698431365
transform 1 0 25872 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_223
timestamp 1698431365
transform 1 0 26320 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_239
timestamp 1698431365
transform 1 0 28112 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_243
timestamp 1698431365
transform 1 0 28560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_255
timestamp 1698431365
transform 1 0 29904 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_294
timestamp 1698431365
transform 1 0 34272 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_298
timestamp 1698431365
transform 1 0 34720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_300
timestamp 1698431365
transform 1 0 34944 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_309
timestamp 1698431365
transform 1 0 35952 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_313
timestamp 1698431365
transform 1 0 36400 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_333
timestamp 1698431365
transform 1 0 38640 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_341
timestamp 1698431365
transform 1 0 39536 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_347
timestamp 1698431365
transform 1 0 40208 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_351
timestamp 1698431365
transform 1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_363
timestamp 1698431365
transform 1 0 42000 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_379
timestamp 1698431365
transform 1 0 43792 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_383
timestamp 1698431365
transform 1 0 44240 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_18
timestamp 1698431365
transform 1 0 3360 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_40
timestamp 1698431365
transform 1 0 5824 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_44
timestamp 1698431365
transform 1 0 6272 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_60
timestamp 1698431365
transform 1 0 8064 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_86
timestamp 1698431365
transform 1 0 10976 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_88
timestamp 1698431365
transform 1 0 11200 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_103
timestamp 1698431365
transform 1 0 12880 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_111
timestamp 1698431365
transform 1 0 13776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_119
timestamp 1698431365
transform 1 0 14672 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_123
timestamp 1698431365
transform 1 0 15120 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_167
timestamp 1698431365
transform 1 0 20048 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_171
timestamp 1698431365
transform 1 0 20496 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_203
timestamp 1698431365
transform 1 0 24080 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_207
timestamp 1698431365
transform 1 0 24528 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_209
timestamp 1698431365
transform 1 0 24752 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_218
timestamp 1698431365
transform 1 0 25760 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_222
timestamp 1698431365
transform 1 0 26208 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_238
timestamp 1698431365
transform 1 0 28000 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_240
timestamp 1698431365
transform 1 0 28224 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_243
timestamp 1698431365
transform 1 0 28560 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_253
timestamp 1698431365
transform 1 0 29680 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_257
timestamp 1698431365
transform 1 0 30128 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_273
timestamp 1698431365
transform 1 0 31920 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_277
timestamp 1698431365
transform 1 0 32368 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_279
timestamp 1698431365
transform 1 0 32592 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_287
timestamp 1698431365
transform 1 0 33488 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_303
timestamp 1698431365
transform 1 0 35280 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_307
timestamp 1698431365
transform 1 0 35728 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_317
timestamp 1698431365
transform 1 0 36848 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_326
timestamp 1698431365
transform 1 0 37856 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_330
timestamp 1698431365
transform 1 0 38304 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_340
timestamp 1698431365
transform 1 0 39424 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_383
timestamp 1698431365
transform 1 0 44240 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_53
timestamp 1698431365
transform 1 0 7280 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_61
timestamp 1698431365
transform 1 0 8176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_71
timestamp 1698431365
transform 1 0 9296 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_81
timestamp 1698431365
transform 1 0 10416 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_85
timestamp 1698431365
transform 1 0 10864 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698431365
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_115
timestamp 1698431365
transform 1 0 14224 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_167
timestamp 1698431365
transform 1 0 20048 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698431365
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_193
timestamp 1698431365
transform 1 0 22960 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_201
timestamp 1698431365
transform 1 0 23856 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_203
timestamp 1698431365
transform 1 0 24080 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_216
timestamp 1698431365
transform 1 0 25536 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_232
timestamp 1698431365
transform 1 0 27328 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_299
timestamp 1698431365
transform 1 0 34832 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_350
timestamp 1698431365
transform 1 0 40544 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_366
timestamp 1698431365
transform 1 0 42336 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_371
timestamp 1698431365
transform 1 0 42896 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_379
timestamp 1698431365
transform 1 0 43792 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_383
timestamp 1698431365
transform 1 0 44240 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698431365
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_76
timestamp 1698431365
transform 1 0 9856 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_132
timestamp 1698431365
transform 1 0 16128 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698431365
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_150
timestamp 1698431365
transform 1 0 18144 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_182
timestamp 1698431365
transform 1 0 21728 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_198
timestamp 1698431365
transform 1 0 23520 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_209
timestamp 1698431365
transform 1 0 24752 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_228
timestamp 1698431365
transform 1 0 26880 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_230
timestamp 1698431365
transform 1 0 27104 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_260
timestamp 1698431365
transform 1 0 30464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_264
timestamp 1698431365
transform 1 0 30912 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_272
timestamp 1698431365
transform 1 0 31808 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_276
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_333
timestamp 1698431365
transform 1 0 38640 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698431365
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_41
timestamp 1698431365
transform 1 0 5936 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_136
timestamp 1698431365
transform 1 0 16576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_140
timestamp 1698431365
transform 1 0 17024 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_172
timestamp 1698431365
transform 1 0 20608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_174
timestamp 1698431365
transform 1 0 20832 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_193
timestamp 1698431365
transform 1 0 22960 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_201
timestamp 1698431365
transform 1 0 23856 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_215
timestamp 1698431365
transform 1 0 25424 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_231
timestamp 1698431365
transform 1 0 27216 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_239
timestamp 1698431365
transform 1 0 28112 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_243
timestamp 1698431365
transform 1 0 28560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_279
timestamp 1698431365
transform 1 0 32592 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_281
timestamp 1698431365
transform 1 0 32816 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_301
timestamp 1698431365
transform 1 0 35056 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_309
timestamp 1698431365
transform 1 0 35952 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_323
timestamp 1698431365
transform 1 0 37520 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_331
timestamp 1698431365
transform 1 0 38416 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_341
timestamp 1698431365
transform 1 0 39536 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_373
timestamp 1698431365
transform 1 0 43120 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_381
timestamp 1698431365
transform 1 0 44016 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_383
timestamp 1698431365
transform 1 0 44240 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_39
timestamp 1698431365
transform 1 0 5712 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_43
timestamp 1698431365
transform 1 0 6160 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_65
timestamp 1698431365
transform 1 0 8624 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_82
timestamp 1698431365
transform 1 0 10528 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_114
timestamp 1698431365
transform 1 0 14112 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_130
timestamp 1698431365
transform 1 0 15904 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_138
timestamp 1698431365
transform 1 0 16800 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_174
timestamp 1698431365
transform 1 0 20832 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_190
timestamp 1698431365
transform 1 0 22624 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_198
timestamp 1698431365
transform 1 0 23520 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_208
timestamp 1698431365
transform 1 0 24640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_220
timestamp 1698431365
transform 1 0 25984 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_252
timestamp 1698431365
transform 1 0 29568 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_268
timestamp 1698431365
transform 1 0 31360 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_272
timestamp 1698431365
transform 1 0 31808 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_311
timestamp 1698431365
transform 1 0 36176 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_315
timestamp 1698431365
transform 1 0 36624 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_347
timestamp 1698431365
transform 1 0 40208 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_349
timestamp 1698431365
transform 1 0 40432 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_45
timestamp 1698431365
transform 1 0 6384 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_75
timestamp 1698431365
transform 1 0 9744 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_87
timestamp 1698431365
transform 1 0 11088 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_91
timestamp 1698431365
transform 1 0 11536 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_99
timestamp 1698431365
transform 1 0 12432 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_103
timestamp 1698431365
transform 1 0 12880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698431365
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698431365
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_253
timestamp 1698431365
transform 1 0 29680 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_269
timestamp 1698431365
transform 1 0 31472 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_277
timestamp 1698431365
transform 1 0 32368 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_281
timestamp 1698431365
transform 1 0 32816 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_297
timestamp 1698431365
transform 1 0 34608 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_313
timestamp 1698431365
transform 1 0 36400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_333
timestamp 1698431365
transform 1 0 38640 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_341
timestamp 1698431365
transform 1 0 39536 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_345
timestamp 1698431365
transform 1 0 39984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_347
timestamp 1698431365
transform 1 0 40208 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_362
timestamp 1698431365
transform 1 0 41888 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_366
timestamp 1698431365
transform 1 0 42336 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_382
timestamp 1698431365
transform 1 0 44128 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698431365
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_104
timestamp 1698431365
transform 1 0 12992 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_108
timestamp 1698431365
transform 1 0 13440 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_110
timestamp 1698431365
transform 1 0 13664 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_117
timestamp 1698431365
transform 1 0 14448 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_133
timestamp 1698431365
transform 1 0 16240 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_137
timestamp 1698431365
transform 1 0 16688 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_139
timestamp 1698431365
transform 1 0 16912 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_150
timestamp 1698431365
transform 1 0 18144 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_154
timestamp 1698431365
transform 1 0 18592 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_156
timestamp 1698431365
transform 1 0 18816 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_161
timestamp 1698431365
transform 1 0 19376 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_193
timestamp 1698431365
transform 1 0 22960 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_209
timestamp 1698431365
transform 1 0 24752 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698431365
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_314
timestamp 1698431365
transform 1 0 36512 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_324
timestamp 1698431365
transform 1 0 37632 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_340
timestamp 1698431365
transform 1 0 39424 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_383
timestamp 1698431365
transform 1 0 44240 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_115
timestamp 1698431365
transform 1 0 14224 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_124
timestamp 1698431365
transform 1 0 15232 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_132
timestamp 1698431365
transform 1 0 16128 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_134
timestamp 1698431365
transform 1 0 16352 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_139
timestamp 1698431365
transform 1 0 16912 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_147
timestamp 1698431365
transform 1 0 17808 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_149
timestamp 1698431365
transform 1 0 18032 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_169
timestamp 1698431365
transform 1 0 20272 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_183
timestamp 1698431365
transform 1 0 21840 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_215
timestamp 1698431365
transform 1 0 25424 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_225
timestamp 1698431365
transform 1 0 26544 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_229
timestamp 1698431365
transform 1 0 26992 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_231
timestamp 1698431365
transform 1 0 27216 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_244
timestamp 1698431365
transform 1 0 28672 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_252
timestamp 1698431365
transform 1 0 29568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_284
timestamp 1698431365
transform 1 0 33152 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_308
timestamp 1698431365
transform 1 0 35840 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_312
timestamp 1698431365
transform 1 0 36288 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_314
timestamp 1698431365
transform 1 0 36512 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_319
timestamp 1698431365
transform 1 0 37072 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_325
timestamp 1698431365
transform 1 0 37744 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_341
timestamp 1698431365
transform 1 0 39536 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_345
timestamp 1698431365
transform 1 0 39984 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_356
timestamp 1698431365
transform 1 0 41216 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_372
timestamp 1698431365
transform 1 0 43008 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_380
timestamp 1698431365
transform 1 0 43904 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_76
timestamp 1698431365
transform 1 0 9856 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_86
timestamp 1698431365
transform 1 0 10976 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_102
timestamp 1698431365
transform 1 0 12768 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_111
timestamp 1698431365
transform 1 0 13776 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_115
timestamp 1698431365
transform 1 0 14224 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_129
timestamp 1698431365
transform 1 0 15792 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_137
timestamp 1698431365
transform 1 0 16688 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_139
timestamp 1698431365
transform 1 0 16912 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_171
timestamp 1698431365
transform 1 0 20496 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_173
timestamp 1698431365
transform 1 0 20720 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_186
timestamp 1698431365
transform 1 0 22176 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_202
timestamp 1698431365
transform 1 0 23968 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_235
timestamp 1698431365
transform 1 0 27664 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_267
timestamp 1698431365
transform 1 0 31248 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_275
timestamp 1698431365
transform 1 0 32144 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_279
timestamp 1698431365
transform 1 0 32592 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_290
timestamp 1698431365
transform 1 0 33824 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_294
timestamp 1698431365
transform 1 0 34272 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_300
timestamp 1698431365
transform 1 0 34944 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_308
timestamp 1698431365
transform 1 0 35840 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_310
timestamp 1698431365
transform 1 0 36064 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_321
timestamp 1698431365
transform 1 0 37296 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_337
timestamp 1698431365
transform 1 0 39088 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_345
timestamp 1698431365
transform 1 0 39984 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_349
timestamp 1698431365
transform 1 0 40432 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_45
timestamp 1698431365
transform 1 0 6384 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_53
timestamp 1698431365
transform 1 0 7280 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_85
timestamp 1698431365
transform 1 0 10864 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_93
timestamp 1698431365
transform 1 0 11760 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_124
timestamp 1698431365
transform 1 0 15232 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_128
timestamp 1698431365
transform 1 0 15680 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_144
timestamp 1698431365
transform 1 0 17472 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_148
timestamp 1698431365
transform 1 0 17920 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_162
timestamp 1698431365
transform 1 0 19488 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_164
timestamp 1698431365
transform 1 0 19712 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698431365
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_193
timestamp 1698431365
transform 1 0 22960 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_201
timestamp 1698431365
transform 1 0 23856 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_214
timestamp 1698431365
transform 1 0 25312 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_226
timestamp 1698431365
transform 1 0 26656 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_242
timestamp 1698431365
transform 1 0 28448 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_244
timestamp 1698431365
transform 1 0 28672 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_263
timestamp 1698431365
transform 1 0 30800 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_271
timestamp 1698431365
transform 1 0 31696 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_279
timestamp 1698431365
transform 1 0 32592 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_283
timestamp 1698431365
transform 1 0 33040 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_302
timestamp 1698431365
transform 1 0 35168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_306
timestamp 1698431365
transform 1 0 35616 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_314
timestamp 1698431365
transform 1 0 36512 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_325
timestamp 1698431365
transform 1 0 37744 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_333
timestamp 1698431365
transform 1 0 38640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_343
timestamp 1698431365
transform 1 0 39760 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_347
timestamp 1698431365
transform 1 0 40208 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_349
timestamp 1698431365
transform 1 0 40432 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_352
timestamp 1698431365
transform 1 0 40768 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_10
timestamp 1698431365
transform 1 0 2464 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_12
timestamp 1698431365
transform 1 0 2688 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_42
timestamp 1698431365
transform 1 0 6048 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_46
timestamp 1698431365
transform 1 0 6496 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_62
timestamp 1698431365
transform 1 0 8288 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_74
timestamp 1698431365
transform 1 0 9632 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_93
timestamp 1698431365
transform 1 0 11760 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_135
timestamp 1698431365
transform 1 0 16464 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_139
timestamp 1698431365
transform 1 0 16912 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_158
timestamp 1698431365
transform 1 0 19040 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_162
timestamp 1698431365
transform 1 0 19488 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_165
timestamp 1698431365
transform 1 0 19824 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_197
timestamp 1698431365
transform 1 0 23408 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_205
timestamp 1698431365
transform 1 0 24304 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698431365
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_218
timestamp 1698431365
transform 1 0 25760 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_234
timestamp 1698431365
transform 1 0 27552 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_242
timestamp 1698431365
transform 1 0 28448 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_272
timestamp 1698431365
transform 1 0 31808 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698431365
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_290
timestamp 1698431365
transform 1 0 33824 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_296
timestamp 1698431365
transform 1 0 34496 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_328
timestamp 1698431365
transform 1 0 38080 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_383
timestamp 1698431365
transform 1 0 44240 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_33
timestamp 1698431365
transform 1 0 5040 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_41
timestamp 1698431365
transform 1 0 5936 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_43
timestamp 1698431365
transform 1 0 6160 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_73
timestamp 1698431365
transform 1 0 9520 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_77
timestamp 1698431365
transform 1 0 9968 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_85
timestamp 1698431365
transform 1 0 10864 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_89
timestamp 1698431365
transform 1 0 11312 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_96
timestamp 1698431365
transform 1 0 12096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_100
timestamp 1698431365
transform 1 0 12544 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_104
timestamp 1698431365
transform 1 0 12992 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_171
timestamp 1698431365
transform 1 0 20496 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_185
timestamp 1698431365
transform 1 0 22064 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_218
timestamp 1698431365
transform 1 0 25760 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_222
timestamp 1698431365
transform 1 0 26208 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_238
timestamp 1698431365
transform 1 0 28000 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_242
timestamp 1698431365
transform 1 0 28448 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_244
timestamp 1698431365
transform 1 0 28672 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_263
timestamp 1698431365
transform 1 0 30800 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_271
timestamp 1698431365
transform 1 0 31696 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_301
timestamp 1698431365
transform 1 0 35056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_305
timestamp 1698431365
transform 1 0 35504 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_313
timestamp 1698431365
transform 1 0 36400 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_325
timestamp 1698431365
transform 1 0 37744 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_333
timestamp 1698431365
transform 1 0 38640 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_337
timestamp 1698431365
transform 1 0 39088 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_346
timestamp 1698431365
transform 1 0 40096 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_350
timestamp 1698431365
transform 1 0 40544 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_354
timestamp 1698431365
transform 1 0 40992 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_370
timestamp 1698431365
transform 1 0 42784 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_378
timestamp 1698431365
transform 1 0 43680 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_382
timestamp 1698431365
transform 1 0 44128 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_66
timestamp 1698431365
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_88
timestamp 1698431365
transform 1 0 11200 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_96
timestamp 1698431365
transform 1 0 12096 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_98
timestamp 1698431365
transform 1 0 12320 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_103
timestamp 1698431365
transform 1 0 12880 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_107
timestamp 1698431365
transform 1 0 13328 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_109
timestamp 1698431365
transform 1 0 13552 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_118
timestamp 1698431365
transform 1 0 14560 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_120
timestamp 1698431365
transform 1 0 14784 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_131
timestamp 1698431365
transform 1 0 16016 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_139
timestamp 1698431365
transform 1 0 16912 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_206
timestamp 1698431365
transform 1 0 24416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_276
timestamp 1698431365
transform 1 0 32256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_346
timestamp 1698431365
transform 1 0 40096 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_53
timestamp 1698431365
transform 1 0 7280 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_57
timestamp 1698431365
transform 1 0 7728 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_64
timestamp 1698431365
transform 1 0 8512 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_80
timestamp 1698431365
transform 1 0 10304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_98
timestamp 1698431365
transform 1 0 12320 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_102
timestamp 1698431365
transform 1 0 12768 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_104
timestamp 1698431365
transform 1 0 12992 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_111
timestamp 1698431365
transform 1 0 13776 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_120
timestamp 1698431365
transform 1 0 14784 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_128
timestamp 1698431365
transform 1 0 15680 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_143
timestamp 1698431365
transform 1 0 17360 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_145
timestamp 1698431365
transform 1 0 17584 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_181
timestamp 1698431365
transform 1 0 21616 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_213
timestamp 1698431365
transform 1 0 25200 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_229
timestamp 1698431365
transform 1 0 26992 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_237
timestamp 1698431365
transform 1 0 27888 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_243
timestamp 1698431365
transform 1 0 28560 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_255
timestamp 1698431365
transform 1 0 29904 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_259
timestamp 1698431365
transform 1 0 30352 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_261
timestamp 1698431365
transform 1 0 30576 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_291
timestamp 1698431365
transform 1 0 33936 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_295
timestamp 1698431365
transform 1 0 34384 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_311
timestamp 1698431365
transform 1 0 36176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_321
timestamp 1698431365
transform 1 0 37296 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_358
timestamp 1698431365
transform 1 0 41440 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_366
timestamp 1698431365
transform 1 0 42336 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_371
timestamp 1698431365
transform 1 0 42896 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_379
timestamp 1698431365
transform 1 0 43792 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_383
timestamp 1698431365
transform 1 0 44240 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_35
timestamp 1698431365
transform 1 0 5264 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_39
timestamp 1698431365
transform 1 0 5712 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_76
timestamp 1698431365
transform 1 0 9856 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_84
timestamp 1698431365
transform 1 0 10752 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_88
timestamp 1698431365
transform 1 0 11200 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_102
timestamp 1698431365
transform 1 0 12768 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_110
timestamp 1698431365
transform 1 0 13664 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_114
timestamp 1698431365
transform 1 0 14112 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_121
timestamp 1698431365
transform 1 0 14896 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_123
timestamp 1698431365
transform 1 0 15120 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_129
timestamp 1698431365
transform 1 0 15792 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_133
timestamp 1698431365
transform 1 0 16240 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_158
timestamp 1698431365
transform 1 0 19040 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_197
timestamp 1698431365
transform 1 0 23408 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_205
timestamp 1698431365
transform 1 0 24304 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_209
timestamp 1698431365
transform 1 0 24752 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_270
timestamp 1698431365
transform 1 0 31584 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_274
timestamp 1698431365
transform 1 0 32032 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_278
timestamp 1698431365
transform 1 0 32480 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_290
timestamp 1698431365
transform 1 0 33824 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_294
timestamp 1698431365
transform 1 0 34272 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_325
timestamp 1698431365
transform 1 0 37744 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_329
timestamp 1698431365
transform 1 0 38192 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_345
timestamp 1698431365
transform 1 0 39984 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_347
timestamp 1698431365
transform 1 0 40208 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_382
timestamp 1698431365
transform 1 0 44128 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_101
timestamp 1698431365
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_171
timestamp 1698431365
transform 1 0 20496 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_241
timestamp 1698431365
transform 1 0 28336 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_311
timestamp 1698431365
transform 1 0 36176 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_333
timestamp 1698431365
transform 1 0 38640 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_341
timestamp 1698431365
transform 1 0 39536 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_345
timestamp 1698431365
transform 1 0 39984 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_353
timestamp 1698431365
transform 1 0 40880 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_357
timestamp 1698431365
transform 1 0 41328 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_18
timestamp 1698431365
transform 1 0 3360 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_26
timestamp 1698431365
transform 1 0 4256 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_30
timestamp 1698431365
transform 1 0 4704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_36
timestamp 1698431365
transform 1 0 5376 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_38
timestamp 1698431365
transform 1 0 5600 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_45
timestamp 1698431365
transform 1 0 6384 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_61
timestamp 1698431365
transform 1 0 8176 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_65
timestamp 1698431365
transform 1 0 8624 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_70
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_79
timestamp 1698431365
transform 1 0 10192 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_95
timestamp 1698431365
transform 1 0 11984 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_99
timestamp 1698431365
transform 1 0 12432 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_101
timestamp 1698431365
transform 1 0 12656 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_104
timestamp 1698431365
transform 1 0 12992 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_106
timestamp 1698431365
transform 1 0 13216 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_133
timestamp 1698431365
transform 1 0 16240 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_135
timestamp 1698431365
transform 1 0 16464 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_138
timestamp 1698431365
transform 1 0 16800 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_140
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_167
timestamp 1698431365
transform 1 0 20048 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_169
timestamp 1698431365
transform 1 0 20272 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_172
timestamp 1698431365
transform 1 0 20608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_174
timestamp 1698431365
transform 1 0 20832 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_201
timestamp 1698431365
transform 1 0 23856 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_203
timestamp 1698431365
transform 1 0 24080 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_206
timestamp 1698431365
transform 1 0 24416 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_208
timestamp 1698431365
transform 1 0 24640 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_235
timestamp 1698431365
transform 1 0 27664 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_237
timestamp 1698431365
transform 1 0 27888 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_240
timestamp 1698431365
transform 1 0 28224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_242
timestamp 1698431365
transform 1 0 28448 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_269
timestamp 1698431365
transform 1 0 31472 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_271
timestamp 1698431365
transform 1 0 31696 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_274
timestamp 1698431365
transform 1 0 32032 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_276
timestamp 1698431365
transform 1 0 32256 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_303
timestamp 1698431365
transform 1 0 35280 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_305
timestamp 1698431365
transform 1 0 35504 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_308
timestamp 1698431365
transform 1 0 35840 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_310
timestamp 1698431365
transform 1 0 36064 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_337
timestamp 1698431365
transform 1 0 39088 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_339
timestamp 1698431365
transform 1 0 39312 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_342
timestamp 1698431365
transform 1 0 39648 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_344
timestamp 1698431365
transform 1 0 39872 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_371
timestamp 1698431365
transform 1 0 42896 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_373
timestamp 1698431365
transform 1 0 43120 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_376
timestamp 1698431365
transform 1 0 43456 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input1
timestamp 1698431365
transform 1 0 9520 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input2
timestamp 1698431365
transform 1 0 5712 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698431365
transform 1 0 17136 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698431365
transform 1 0 20944 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698431365
transform 1 0 24752 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698431365
transform 1 0 28560 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698431365
transform 1 0 32368 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698431365
transform 1 0 36176 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698431365
transform 1 0 39984 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698431365
transform -1 0 44352 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_50 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 44576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_51
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 44576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_52
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 44576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_53
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 44576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_54
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 44576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_55
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 44576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_56
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 44576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_57
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 44576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_58
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 44576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_59
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 44576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_60
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 44576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_61
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 44576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_62
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 44576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_63
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 44576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_64
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 44576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_65
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 44576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_66
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 44576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_67
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 44576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_68
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 44576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_69
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 44576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_70
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 44576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_71
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 44576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_72
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 44576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_73
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 44576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_74
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 44576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_75
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 44576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_76
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 44576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_77
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 44576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_78
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 44576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 44576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 44576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 44576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 44576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 44576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 44576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 44576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 44576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 44576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 44576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 44576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 44576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 44576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 44576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 44576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 44576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 44576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 44576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 44576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 44576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 44576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_100 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_101
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_102
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_103
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_104
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_105
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_106
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_107
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_108
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_109
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_110
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_111
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_112
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_113
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_114
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_115
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_116
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_117
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_118
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_119
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_120
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_121
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_122
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_123
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_124
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_125
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_126
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_127
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_128
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_129
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_130
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_131
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_132
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_133
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_134
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_135
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_136
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_137
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_138
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_139
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_140
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_141
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_142
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_143
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_144
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_145
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_146
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_147
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_148
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_149
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_150
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_151
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_152
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_153
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_154
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_155
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_156
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_157
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_158
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_159
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_160
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_161
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_162
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_163
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_164
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_165
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_166
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_167
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_168
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_169
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_170
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_171
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_172
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_173
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_174
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_175
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_176
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_177
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_178
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_179
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_180
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_181
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_182
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_183
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_184
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_185
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_186
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_187
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_188
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_189
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_190
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_191
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_192
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_193
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_194
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_195
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_196
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_197
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_198
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_199
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_200
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_201
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_202
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_203
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_204
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_205
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_206
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_207
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_208
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_209
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_210
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_211
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_212
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_213
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_214
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_215
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_216
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_217
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_218
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_219
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_220
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_221
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_222
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_223
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_224
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_225
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_226
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_227
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_228
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_229
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_230
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_231
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_232
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_233
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_234
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_235
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_236
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_237
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_238
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_239
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_240
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_241
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_242
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_243
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_244
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_245
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_246
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_247
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_248
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_249
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_250
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_251
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_252
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_253
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_254
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_255
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_256
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_257
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_258
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_259
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_260
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_261
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_262
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_263
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_264
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_265
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_266
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_267
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_268
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_269
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_270
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_271
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_272
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_273
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_274
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_275
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_276
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_277
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_278
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_279
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_280
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_281
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_282
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_283
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_284
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_285
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_286
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_287
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_288
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_289
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_290
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_291
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_292
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_293
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_294
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_295
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_296
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_297
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_298
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_299
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_300
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_301
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_302
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_303
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_304
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_305
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_306
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_307
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_308
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_309
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_310
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_311
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_312
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_313
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_314
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_315
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_316
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_317
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_318
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_319
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_320
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_321
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_322
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_323
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_324
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_325
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_326
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_327
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_328
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_329
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_330
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_331
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_332
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_333
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_334
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_335
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_336
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_337
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_338
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_339
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_340
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_341
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_342
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_343
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_344
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_345
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_346
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_347
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_348
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_349
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_350
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_351
timestamp 1698431365
transform 1 0 5152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_352
timestamp 1698431365
transform 1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_353
timestamp 1698431365
transform 1 0 12768 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_354
timestamp 1698431365
transform 1 0 16576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_355
timestamp 1698431365
transform 1 0 20384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_356
timestamp 1698431365
transform 1 0 24192 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_357
timestamp 1698431365
transform 1 0 28000 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_358
timestamp 1698431365
transform 1 0 31808 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_359
timestamp 1698431365
transform 1 0 35616 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_360
timestamp 1698431365
transform 1 0 39424 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_361
timestamp 1698431365
transform 1 0 43232 0 -1 42336
box -86 -86 310 870
<< labels >>
flabel metal2 s 9408 45200 9520 46000 0 FreeSans 448 90 0 0 io_in
port 0 nsew signal input
flabel metal2 s 13216 45200 13328 46000 0 FreeSans 448 90 0 0 io_out[0]
port 1 nsew signal tristate
flabel metal2 s 17024 45200 17136 46000 0 FreeSans 448 90 0 0 io_out[1]
port 2 nsew signal tristate
flabel metal2 s 20832 45200 20944 46000 0 FreeSans 448 90 0 0 io_out[2]
port 3 nsew signal tristate
flabel metal2 s 24640 45200 24752 46000 0 FreeSans 448 90 0 0 io_out[3]
port 4 nsew signal tristate
flabel metal2 s 28448 45200 28560 46000 0 FreeSans 448 90 0 0 io_out[4]
port 5 nsew signal tristate
flabel metal2 s 32256 45200 32368 46000 0 FreeSans 448 90 0 0 io_out[5]
port 6 nsew signal tristate
flabel metal2 s 36064 45200 36176 46000 0 FreeSans 448 90 0 0 io_out[6]
port 7 nsew signal tristate
flabel metal2 s 39872 45200 39984 46000 0 FreeSans 448 90 0 0 io_out[7]
port 8 nsew signal tristate
flabel metal2 s 43680 45200 43792 46000 0 FreeSans 448 90 0 0 io_out[8]
port 9 nsew signal tristate
flabel metal2 s 5600 45200 5712 46000 0 FreeSans 448 90 0 0 rst_n
port 10 nsew signal input
flabel metal4 s 4448 3076 4768 42396 0 FreeSans 1280 90 0 0 vdd
port 11 nsew power bidirectional
flabel metal4 s 35168 3076 35488 42396 0 FreeSans 1280 90 0 0 vdd
port 11 nsew power bidirectional
flabel metal4 s 19808 3076 20128 42396 0 FreeSans 1280 90 0 0 vss
port 12 nsew ground bidirectional
flabel metal2 s 1792 45200 1904 46000 0 FreeSans 448 90 0 0 wb_clk_i
port 13 nsew signal input
rlabel metal1 22960 41552 22960 41552 0 vdd
rlabel metal1 22960 42336 22960 42336 0 vss
rlabel metal3 7168 40376 7168 40376 0 _000_
rlabel metal3 16800 40264 16800 40264 0 _001_
rlabel metal2 26040 39816 26040 39816 0 _002_
rlabel metal2 29288 39984 29288 39984 0 _003_
rlabel metal2 31640 40096 31640 40096 0 _004_
rlabel metal3 17136 39592 17136 39592 0 _005_
rlabel metal2 8008 39872 8008 39872 0 _006_
rlabel metal2 34664 18704 34664 18704 0 _007_
rlabel metal2 30184 19656 30184 19656 0 _008_
rlabel metal2 31752 15456 31752 15456 0 _009_
rlabel metal3 38472 16184 38472 16184 0 _010_
rlabel metal3 37632 13048 37632 13048 0 _011_
rlabel metal2 35560 9800 35560 9800 0 _012_
rlabel metal2 35224 6440 35224 6440 0 _013_
rlabel metal2 29176 10248 29176 10248 0 _014_
rlabel metal2 31304 5488 31304 5488 0 _015_
rlabel metal2 25256 5432 25256 5432 0 _016_
rlabel metal2 11928 39312 11928 39312 0 _017_
rlabel metal3 12096 38808 12096 38808 0 _018_
rlabel metal2 2744 38528 2744 38528 0 _019_
rlabel metal2 34552 37240 34552 37240 0 _020_
rlabel metal2 30856 36848 30856 36848 0 _021_
rlabel metal2 37128 39200 37128 39200 0 _022_
rlabel metal2 40320 40264 40320 40264 0 _023_
rlabel metal2 41328 33544 41328 33544 0 _024_
rlabel metal2 41944 37576 41944 37576 0 _025_
rlabel metal2 38472 37296 38472 37296 0 _026_
rlabel metal3 33656 32200 33656 32200 0 _027_
rlabel metal2 33992 28672 33992 28672 0 _028_
rlabel metal2 39592 30576 39592 30576 0 _029_
rlabel metal2 41944 29008 41944 29008 0 _030_
rlabel metal2 41384 24976 41384 24976 0 _031_
rlabel metal2 41496 22120 41496 22120 0 _032_
rlabel metal2 37128 21728 37128 21728 0 _033_
rlabel metal2 31752 24304 31752 24304 0 _034_
rlabel metal2 35448 25648 35448 25648 0 _035_
rlabel metal2 19992 19040 19992 19040 0 _036_
rlabel metal2 2632 18760 2632 18760 0 _037_
rlabel metal2 6776 17192 6776 17192 0 _038_
rlabel metal2 14728 18200 14728 18200 0 _039_
rlabel metal2 2632 10920 2632 10920 0 _040_
rlabel metal2 2632 13720 2632 13720 0 _041_
rlabel metal2 7784 9128 7784 9128 0 _042_
rlabel metal3 16688 13048 16688 13048 0 _043_
rlabel metal2 11088 9912 11088 9912 0 _044_
rlabel metal2 13160 4704 13160 4704 0 _045_
rlabel metal2 18088 5992 18088 5992 0 _046_
rlabel metal2 21784 5432 21784 5432 0 _047_
rlabel metal2 22568 7784 22568 7784 0 _048_
rlabel metal3 25816 11256 25816 11256 0 _049_
rlabel metal3 25928 13832 25928 13832 0 _050_
rlabel metal3 24920 19096 24920 19096 0 _051_
rlabel metal2 8344 32984 8344 32984 0 _052_
rlabel metal2 2968 24640 2968 24640 0 _053_
rlabel metal2 2912 31640 2912 31640 0 _054_
rlabel metal2 5096 30240 5096 30240 0 _055_
rlabel metal2 3192 23856 3192 23856 0 _056_
rlabel metal2 20216 30240 20216 30240 0 _057_
rlabel metal2 15848 31416 15848 31416 0 _058_
rlabel metal2 21000 26600 21000 26600 0 _059_
rlabel metal2 29512 30072 29512 30072 0 _060_
rlabel metal2 24360 34104 24360 34104 0 _061_
rlabel metal2 23576 29008 23576 29008 0 _062_
rlabel metal2 27552 26152 27552 26152 0 _063_
rlabel metal2 21784 35952 21784 35952 0 _064_
rlabel metal3 23856 34888 23856 34888 0 _065_
rlabel metal2 25256 31780 25256 31780 0 _066_
rlabel metal2 25760 34888 25760 34888 0 _067_
rlabel metal2 26264 35504 26264 35504 0 _068_
rlabel metal2 25928 35336 25928 35336 0 _069_
rlabel metal2 18424 35504 18424 35504 0 _070_
rlabel metal2 25032 31836 25032 31836 0 _071_
rlabel metal2 27496 34384 27496 34384 0 _072_
rlabel metal2 19376 35672 19376 35672 0 _073_
rlabel metal2 18256 35112 18256 35112 0 _074_
rlabel metal2 19096 35112 19096 35112 0 _075_
rlabel metal2 21000 36120 21000 36120 0 _076_
rlabel metal3 17808 35448 17808 35448 0 _077_
rlabel metal3 12936 29400 12936 29400 0 _078_
rlabel metal2 8232 24752 8232 24752 0 _079_
rlabel metal2 15624 26152 15624 26152 0 _080_
rlabel metal2 16240 24808 16240 24808 0 _081_
rlabel metal2 12488 25984 12488 25984 0 _082_
rlabel metal2 10808 25144 10808 25144 0 _083_
rlabel metal3 13104 25480 13104 25480 0 _084_
rlabel metal2 30632 21224 30632 21224 0 _085_
rlabel metal2 30408 21280 30408 21280 0 _086_
rlabel metal2 30184 21168 30184 21168 0 _087_
rlabel metal2 29792 26936 29792 26936 0 _088_
rlabel metal2 17640 26208 17640 26208 0 _089_
rlabel metal2 17696 23800 17696 23800 0 _090_
rlabel metal2 17304 20412 17304 20412 0 _091_
rlabel metal3 25368 15344 25368 15344 0 _092_
rlabel metal2 11032 12320 11032 12320 0 _093_
rlabel metal2 10304 20216 10304 20216 0 _094_
rlabel metal3 9408 21560 9408 21560 0 _095_
rlabel metal2 17080 21280 17080 21280 0 _096_
rlabel metal2 15736 22400 15736 22400 0 _097_
rlabel metal3 15624 28616 15624 28616 0 _098_
rlabel metal2 12264 24696 12264 24696 0 _099_
rlabel metal2 10472 21896 10472 21896 0 _100_
rlabel metal2 11368 23408 11368 23408 0 _101_
rlabel metal2 15176 23408 15176 23408 0 _102_
rlabel metal3 11256 26264 11256 26264 0 _103_
rlabel metal2 10024 20440 10024 20440 0 _104_
rlabel metal2 9016 24864 9016 24864 0 _105_
rlabel metal2 11368 20776 11368 20776 0 _106_
rlabel metal3 15680 14392 15680 14392 0 _107_
rlabel metal2 15176 19768 15176 19768 0 _108_
rlabel metal3 11760 19992 11760 19992 0 _109_
rlabel metal2 15512 20496 15512 20496 0 _110_
rlabel metal2 10696 18592 10696 18592 0 _111_
rlabel metal3 9464 22344 9464 22344 0 _112_
rlabel metal2 13832 21448 13832 21448 0 _113_
rlabel metal2 9016 20272 9016 20272 0 _114_
rlabel metal3 7952 23688 7952 23688 0 _115_
rlabel metal3 11704 20552 11704 20552 0 _116_
rlabel metal2 16184 21728 16184 21728 0 _117_
rlabel metal2 16856 29624 16856 29624 0 _118_
rlabel metal2 16296 36848 16296 36848 0 _119_
rlabel metal3 11200 36568 11200 36568 0 _120_
rlabel metal2 15624 36904 15624 36904 0 _121_
rlabel metal3 14560 38808 14560 38808 0 _122_
rlabel metal2 10248 36008 10248 36008 0 _123_
rlabel metal2 10416 35448 10416 35448 0 _124_
rlabel metal2 11256 36568 11256 36568 0 _125_
rlabel metal2 16632 35448 16632 35448 0 _126_
rlabel metal2 19488 35000 19488 35000 0 _127_
rlabel metal3 17052 34664 17052 34664 0 _128_
rlabel metal2 12376 37128 12376 37128 0 _129_
rlabel metal2 12096 39368 12096 39368 0 _130_
rlabel metal2 18088 35896 18088 35896 0 _131_
rlabel metal2 14840 35616 14840 35616 0 _132_
rlabel metal2 13608 35952 13608 35952 0 _133_
rlabel metal3 14448 39480 14448 39480 0 _134_
rlabel metal3 11984 40488 11984 40488 0 _135_
rlabel metal3 22288 24024 22288 24024 0 _136_
rlabel metal2 10920 37464 10920 37464 0 _137_
rlabel metal2 14728 40320 14728 40320 0 _138_
rlabel metal2 12152 40432 12152 40432 0 _139_
rlabel metal2 12600 39984 12600 39984 0 _140_
rlabel metal2 15848 39088 15848 39088 0 _141_
rlabel metal3 15512 39368 15512 39368 0 _142_
rlabel metal2 16240 40600 16240 40600 0 _143_
rlabel metal3 8372 39480 8372 39480 0 _144_
rlabel metal2 25648 23128 25648 23128 0 _145_
rlabel metal2 26040 23296 26040 23296 0 _146_
rlabel metal3 27552 18984 27552 18984 0 _147_
rlabel metal2 31864 18704 31864 18704 0 _148_
rlabel metal2 31416 16352 31416 16352 0 _149_
rlabel metal2 25928 27104 25928 27104 0 _150_
rlabel metal3 21784 26936 21784 26936 0 _151_
rlabel metal2 24472 30968 24472 30968 0 _152_
rlabel metal2 31080 17192 31080 17192 0 _153_
rlabel metal2 31024 16296 31024 16296 0 _154_
rlabel metal2 35336 17584 35336 17584 0 _155_
rlabel metal2 35896 16408 35896 16408 0 _156_
rlabel metal2 24976 21784 24976 21784 0 _157_
rlabel metal2 34776 15960 34776 15960 0 _158_
rlabel metal3 35280 16072 35280 16072 0 _159_
rlabel metal2 36456 16912 36456 16912 0 _160_
rlabel metal2 36064 12824 36064 12824 0 _161_
rlabel metal2 7672 11088 7672 11088 0 _162_
rlabel metal2 35896 13216 35896 13216 0 _163_
rlabel metal2 34552 10080 34552 10080 0 _164_
rlabel metal2 30520 9352 30520 9352 0 _165_
rlabel metal2 35392 10696 35392 10696 0 _166_
rlabel metal3 32704 9128 32704 9128 0 _167_
rlabel metal2 30912 6104 30912 6104 0 _168_
rlabel metal2 33096 8960 33096 8960 0 _169_
rlabel metal3 30296 9800 30296 9800 0 _170_
rlabel metal2 29176 6048 29176 6048 0 _171_
rlabel metal3 29904 5880 29904 5880 0 _172_
rlabel metal2 25872 6104 25872 6104 0 _173_
rlabel metal2 28504 5824 28504 5824 0 _174_
rlabel metal3 26264 5768 26264 5768 0 _175_
rlabel metal3 33152 36232 33152 36232 0 _176_
rlabel metal3 24472 31640 24472 31640 0 _177_
rlabel metal2 24528 32088 24528 32088 0 _178_
rlabel metal2 34440 36680 34440 36680 0 _179_
rlabel metal2 35952 24024 35952 24024 0 _180_
rlabel metal2 28616 29232 28616 29232 0 _181_
rlabel metal2 37352 31780 37352 31780 0 _182_
rlabel metal2 37464 33880 37464 33880 0 _183_
rlabel metal2 36680 36120 36680 36120 0 _184_
rlabel metal2 35000 26768 35000 26768 0 _185_
rlabel metal2 37688 29624 37688 29624 0 _186_
rlabel metal2 34440 35952 34440 35952 0 _187_
rlabel metal2 37688 26656 37688 26656 0 _188_
rlabel metal2 20664 27104 20664 27104 0 _189_
rlabel metal2 37352 37688 37352 37688 0 _190_
rlabel metal2 37520 36568 37520 36568 0 _191_
rlabel metal3 33432 32648 33432 32648 0 _192_
rlabel metal2 40936 35560 40936 35560 0 _193_
rlabel metal2 28280 26992 28280 26992 0 _194_
rlabel metal2 28952 22400 28952 22400 0 _195_
rlabel metal2 28392 29904 28392 29904 0 _196_
rlabel metal2 28504 24136 28504 24136 0 _197_
rlabel metal2 41160 33320 41160 33320 0 _198_
rlabel metal2 40600 33992 40600 33992 0 _199_
rlabel metal2 39648 39368 39648 39368 0 _200_
rlabel metal4 39480 37296 39480 37296 0 _201_
rlabel metal2 37464 35560 37464 35560 0 _202_
rlabel metal2 29120 25256 29120 25256 0 _203_
rlabel metal3 34272 31528 34272 31528 0 _204_
rlabel metal2 33992 31696 33992 31696 0 _205_
rlabel metal2 33768 28896 33768 28896 0 _206_
rlabel metal2 34216 28896 34216 28896 0 _207_
rlabel metal3 40824 29960 40824 29960 0 _208_
rlabel metal2 37240 28000 37240 28000 0 _209_
rlabel metal2 38808 30632 38808 30632 0 _210_
rlabel metal2 41496 27384 41496 27384 0 _211_
rlabel metal2 41384 28112 41384 28112 0 _212_
rlabel metal3 26376 29288 26376 29288 0 _213_
rlabel metal2 41608 22456 41608 22456 0 _214_
rlabel metal2 40936 24864 40936 24864 0 _215_
rlabel metal2 40824 22792 40824 22792 0 _216_
rlabel metal2 41216 22568 41216 22568 0 _217_
rlabel metal2 35728 24136 35728 24136 0 _218_
rlabel metal2 36288 23240 36288 23240 0 _219_
rlabel metal2 37352 23576 37352 23576 0 _220_
rlabel metal2 33432 24024 33432 24024 0 _221_
rlabel metal2 33768 25088 33768 25088 0 _222_
rlabel metal2 35896 25816 35896 25816 0 _223_
rlabel metal2 20328 18984 20328 18984 0 _224_
rlabel metal2 15288 26432 15288 26432 0 _225_
rlabel metal2 16072 25592 16072 25592 0 _226_
rlabel metal2 22904 24584 22904 24584 0 _227_
rlabel metal2 19656 22792 19656 22792 0 _228_
rlabel metal2 21112 23016 21112 23016 0 _229_
rlabel metal2 28952 25256 28952 25256 0 _230_
rlabel metal2 19432 22848 19432 22848 0 _231_
rlabel metal2 19040 22344 19040 22344 0 _232_
rlabel metal2 19600 23688 19600 23688 0 _233_
rlabel metal2 19544 18424 19544 18424 0 _234_
rlabel metal2 10136 18088 10136 18088 0 _235_
rlabel metal2 21896 14056 21896 14056 0 _236_
rlabel metal2 6216 10976 6216 10976 0 _237_
rlabel metal2 18984 18760 18984 18760 0 _238_
rlabel metal2 12040 10976 12040 10976 0 _239_
rlabel metal2 5656 17976 5656 17976 0 _240_
rlabel metal2 5992 17976 5992 17976 0 _241_
rlabel metal2 11256 16856 11256 16856 0 _242_
rlabel metal2 10808 17472 10808 17472 0 _243_
rlabel metal2 10584 17360 10584 17360 0 _244_
rlabel metal2 11032 16856 11032 16856 0 _245_
rlabel metal3 21700 15400 21700 15400 0 _246_
rlabel metal2 17472 16632 17472 16632 0 _247_
rlabel metal3 11872 13944 11872 13944 0 _248_
rlabel metal3 15064 18424 15064 18424 0 _249_
rlabel metal2 6888 12040 6888 12040 0 _250_
rlabel metal2 7000 12992 7000 12992 0 _251_
rlabel metal2 5320 12600 5320 12600 0 _252_
rlabel metal3 5096 11256 5096 11256 0 _253_
rlabel metal3 5600 11368 5600 11368 0 _254_
rlabel metal2 4984 12768 4984 12768 0 _255_
rlabel metal3 5488 12824 5488 12824 0 _256_
rlabel metal3 13272 12824 13272 12824 0 _257_
rlabel metal2 7560 12488 7560 12488 0 _258_
rlabel metal2 8680 12656 8680 12656 0 _259_
rlabel metal3 23912 22960 23912 22960 0 _260_
rlabel metal2 10248 13384 10248 13384 0 _261_
rlabel metal2 9968 12152 9968 12152 0 _262_
rlabel metal2 14952 14056 14952 14056 0 _263_
rlabel metal2 14616 13832 14616 13832 0 _264_
rlabel metal3 13216 10584 13216 10584 0 _265_
rlabel metal2 14952 10472 14952 10472 0 _266_
rlabel metal2 12488 9296 12488 9296 0 _267_
rlabel metal2 11368 9968 11368 9968 0 _268_
rlabel metal3 11984 9688 11984 9688 0 _269_
rlabel metal2 15288 8372 15288 8372 0 _270_
rlabel metal2 14168 10304 14168 10304 0 _271_
rlabel metal2 14280 11536 14280 11536 0 _272_
rlabel metal2 23016 21532 23016 21532 0 _273_
rlabel metal2 13608 11032 13608 11032 0 _274_
rlabel metal2 18256 7784 18256 7784 0 _275_
rlabel metal3 16464 8120 16464 8120 0 _276_
rlabel metal2 22904 17864 22904 17864 0 _277_
rlabel metal2 18760 9744 18760 9744 0 _278_
rlabel metal3 18200 9016 18200 9016 0 _279_
rlabel metal2 18088 8624 18088 8624 0 _280_
rlabel metal3 23296 8344 23296 8344 0 _281_
rlabel metal2 20104 8316 20104 8316 0 _282_
rlabel metal2 19320 8904 19320 8904 0 _283_
rlabel metal3 19432 8232 19432 8232 0 _284_
rlabel metal3 16688 9800 16688 9800 0 _285_
rlabel metal2 20552 13328 20552 13328 0 _286_
rlabel metal2 23128 12544 23128 12544 0 _287_
rlabel metal2 23464 12488 23464 12488 0 _288_
rlabel metal2 22120 11816 22120 11816 0 _289_
rlabel metal3 23240 12152 23240 12152 0 _290_
rlabel metal2 23128 8372 23128 8372 0 _291_
rlabel metal2 24024 13664 24024 13664 0 _292_
rlabel metal2 24360 11760 24360 11760 0 _293_
rlabel metal2 23688 12320 23688 12320 0 _294_
rlabel metal2 23968 11368 23968 11368 0 _295_
rlabel metal3 25088 14728 25088 14728 0 _296_
rlabel metal2 24136 13552 24136 13552 0 _297_
rlabel metal2 23464 16072 23464 16072 0 _298_
rlabel metal3 23296 16296 23296 16296 0 _299_
rlabel metal2 23632 15400 23632 15400 0 _300_
rlabel metal2 24136 17640 24136 17640 0 _301_
rlabel metal2 23352 17864 23352 17864 0 _302_
rlabel metal3 23856 18424 23856 18424 0 _303_
rlabel metal2 24584 18704 24584 18704 0 _304_
rlabel metal2 18872 28560 18872 28560 0 _305_
rlabel metal3 7728 30408 7728 30408 0 _306_
rlabel metal3 9464 32648 9464 32648 0 _307_
rlabel metal2 8344 27048 8344 27048 0 _308_
rlabel metal3 7000 28616 7000 28616 0 _309_
rlabel metal3 5824 28392 5824 28392 0 _310_
rlabel metal2 5992 25592 5992 25592 0 _311_
rlabel metal2 15512 29456 15512 29456 0 _312_
rlabel metal2 4312 28056 4312 28056 0 _313_
rlabel metal2 4312 29120 4312 29120 0 _314_
rlabel metal2 3304 28896 3304 28896 0 _315_
rlabel metal2 4088 28392 4088 28392 0 _316_
rlabel metal2 4872 28728 4872 28728 0 _317_
rlabel metal2 5208 29120 5208 29120 0 _318_
rlabel metal2 10584 28336 10584 28336 0 _319_
rlabel metal2 15736 29064 15736 29064 0 _320_
rlabel metal3 17360 29288 17360 29288 0 _321_
rlabel metal2 3864 26544 3864 26544 0 _322_
rlabel metal2 19320 29624 19320 29624 0 _323_
rlabel metal3 18760 29400 18760 29400 0 _324_
rlabel metal2 17024 29288 17024 29288 0 _325_
rlabel metal2 17192 27664 17192 27664 0 _326_
rlabel metal3 17640 26824 17640 26824 0 _327_
rlabel metal2 15960 30464 15960 30464 0 _328_
rlabel metal3 18592 26264 18592 26264 0 _329_
rlabel metal2 18872 26712 18872 26712 0 _330_
rlabel metal2 29176 29792 29176 29792 0 _331_
rlabel metal2 24248 32592 24248 32592 0 _332_
rlabel metal2 24584 31472 24584 31472 0 _333_
rlabel metal2 24360 32312 24360 32312 0 _334_
rlabel metal2 25312 29512 25312 29512 0 _335_
rlabel metal3 28560 25368 28560 25368 0 _336_
rlabel metal2 9912 37464 9912 37464 0 bcd\[0\]
rlabel metal3 6440 36568 6440 36568 0 bcd\[1\]
rlabel metal3 8960 35784 8960 35784 0 bcd\[2\]
rlabel metal2 9016 33040 9016 33040 0 clkdiv\[0\]
rlabel metal2 6888 23968 6888 23968 0 clkdiv\[1\]
rlabel metal2 5656 30688 5656 30688 0 clkdiv\[2\]
rlabel metal3 8008 30184 8008 30184 0 clkdiv\[3\]
rlabel metal2 6888 22344 6888 22344 0 clkdiv\[4\]
rlabel metal2 18648 30240 18648 30240 0 clkdiv\[5\]
rlabel metal2 12768 25480 12768 25480 0 clkdiv\[6\]
rlabel metal2 23128 26096 23128 26096 0 clkdiv\[7\]
rlabel metal2 29400 30072 29400 30072 0 clknet_0_wb_clk_i
rlabel metal2 7112 8120 7112 8120 0 clknet_3_0__leaf_wb_clk_i
rlabel metal2 20664 18032 20664 18032 0 clknet_3_1__leaf_wb_clk_i
rlabel metal2 5936 40376 5936 40376 0 clknet_3_2__leaf_wb_clk_i
rlabel metal2 21448 40040 21448 40040 0 clknet_3_3__leaf_wb_clk_i
rlabel metal3 26880 7672 26880 7672 0 clknet_3_4__leaf_wb_clk_i
rlabel metal2 32648 5936 32648 5936 0 clknet_3_5__leaf_wb_clk_i
rlabel metal2 30072 25816 30072 25816 0 clknet_3_6__leaf_wb_clk_i
rlabel metal2 37016 30184 37016 30184 0 clknet_3_7__leaf_wb_clk_i
rlabel metal2 20216 18984 20216 18984 0 counter\[0\]
rlabel metal2 20328 5432 20328 5432 0 counter\[10\]
rlabel metal2 20216 9352 20216 9352 0 counter\[11\]
rlabel metal2 24696 7868 24696 7868 0 counter\[12\]
rlabel metal2 25704 14112 25704 14112 0 counter\[13\]
rlabel metal2 29064 15008 29064 15008 0 counter\[14\]
rlabel metal2 27608 17360 27608 17360 0 counter\[15\]
rlabel metal2 6104 19264 6104 19264 0 counter\[1\]
rlabel metal2 9632 16072 9632 16072 0 counter\[2\]
rlabel metal2 16856 17808 16856 17808 0 counter\[3\]
rlabel metal2 4872 11536 4872 11536 0 counter\[4\]
rlabel metal3 5544 14280 5544 14280 0 counter\[5\]
rlabel metal2 9912 8372 9912 8372 0 counter\[6\]
rlabel metal2 15120 14616 15120 14616 0 counter\[7\]
rlabel metal2 13048 6272 13048 6272 0 counter\[8\]
rlabel metal2 15288 4648 15288 4648 0 counter\[9\]
rlabel metal2 9464 44478 9464 44478 0 io_in
rlabel metal3 13888 41832 13888 41832 0 io_out[0]
rlabel metal2 17640 45304 17640 45304 0 io_out[1]
rlabel metal2 21448 45304 21448 45304 0 io_out[2]
rlabel metal3 25312 41832 25312 41832 0 io_out[3]
rlabel metal3 28504 42056 28504 42056 0 io_out[4]
rlabel metal2 32872 45304 32872 45304 0 io_out[5]
rlabel metal3 36736 41832 36736 41832 0 io_out[6]
rlabel metal3 40544 41832 40544 41832 0 io_out[7]
rlabel metal2 43736 43330 43736 43330 0 io_out[8]
rlabel metal3 28896 34888 28896 34888 0 lfsr\[0\]
rlabel metal2 44072 29680 44072 29680 0 lfsr\[10\]
rlabel metal3 43876 25592 43876 25592 0 lfsr\[11\]
rlabel metal2 43624 21168 43624 21168 0 lfsr\[12\]
rlabel metal3 38976 23128 38976 23128 0 lfsr\[13\]
rlabel metal2 33208 23184 33208 23184 0 lfsr\[14\]
rlabel metal2 36904 26488 36904 26488 0 lfsr\[15\]
rlabel metal2 28728 36904 28728 36904 0 lfsr\[1\]
rlabel metal2 34664 35672 34664 35672 0 lfsr\[2\]
rlabel metal2 41608 33488 41608 33488 0 lfsr\[4\]
rlabel metal3 41720 36456 41720 36456 0 lfsr\[5\]
rlabel metal2 41048 39704 41048 39704 0 lfsr\[6\]
rlabel metal3 36848 32424 36848 32424 0 lfsr\[7\]
rlabel metal2 33208 29960 33208 29960 0 lfsr\[8\]
rlabel metal2 37464 29960 37464 29960 0 lfsr\[9\]
rlabel metal2 33544 18872 33544 18872 0 m_clkdiv\[0\]
rlabel metal2 32424 17920 32424 17920 0 m_clkdiv\[1\]
rlabel metal3 30632 16856 30632 16856 0 m_clkdiv\[2\]
rlabel metal2 35896 17248 35896 17248 0 m_clkdiv\[3\]
rlabel metal2 36568 13832 36568 13832 0 m_clkdiv\[4\]
rlabel metal3 36624 11144 36624 11144 0 m_clkdiv\[5\]
rlabel metal2 33544 6216 33544 6216 0 m_clkdiv\[6\]
rlabel metal2 31080 9856 31080 9856 0 m_clkdiv\[7\]
rlabel metal2 30352 6104 30352 6104 0 m_clkdiv\[8\]
rlabel metal2 27496 6272 27496 6272 0 m_clkdiv\[9\]
rlabel metal2 15288 27104 15288 27104 0 net1
rlabel metal2 29736 25368 29736 25368 0 net10
rlabel metal2 43960 40712 43960 40712 0 net11
rlabel metal2 6384 40600 6384 40600 0 net2
rlabel metal3 6748 40264 6748 40264 0 net3
rlabel metal2 9016 40152 9016 40152 0 net4
rlabel metal2 20776 40824 20776 40824 0 net5
rlabel metal2 23240 41104 23240 41104 0 net6
rlabel metal2 28168 41104 28168 41104 0 net7
rlabel metal2 31416 41104 31416 41104 0 net8
rlabel metal2 33768 40824 33768 40824 0 net9
rlabel metal2 29400 33208 29400 33208 0 r_counter\[0\]
rlabel metal2 25200 37240 25200 37240 0 r_counter\[1\]
rlabel metal3 25928 30184 25928 30184 0 r_counter\[2\]
rlabel metal2 5656 44478 5656 44478 0 rst_n
rlabel metal2 21672 22344 21672 22344 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 46000 46000
<< end >>
