magic
tech gf180mcuD
magscale 1 5
timestamp 1699362620
<< obsm1 >>
rect 672 1471 64288 58785
<< metal2 >>
rect 4144 59600 4200 60000
rect 4592 59600 4648 60000
rect 5040 59600 5096 60000
rect 5488 59600 5544 60000
rect 5936 59600 5992 60000
rect 6384 59600 6440 60000
rect 6832 59600 6888 60000
rect 7280 59600 7336 60000
rect 7728 59600 7784 60000
rect 8176 59600 8232 60000
rect 8624 59600 8680 60000
rect 9072 59600 9128 60000
rect 9520 59600 9576 60000
rect 9968 59600 10024 60000
rect 10416 59600 10472 60000
rect 10864 59600 10920 60000
rect 11312 59600 11368 60000
rect 11760 59600 11816 60000
rect 12208 59600 12264 60000
rect 12656 59600 12712 60000
rect 13104 59600 13160 60000
rect 13552 59600 13608 60000
rect 14000 59600 14056 60000
rect 14448 59600 14504 60000
rect 14896 59600 14952 60000
rect 15344 59600 15400 60000
rect 15792 59600 15848 60000
rect 16240 59600 16296 60000
rect 16688 59600 16744 60000
rect 17136 59600 17192 60000
rect 17584 59600 17640 60000
rect 18032 59600 18088 60000
rect 18480 59600 18536 60000
rect 18928 59600 18984 60000
rect 19376 59600 19432 60000
rect 19824 59600 19880 60000
rect 20272 59600 20328 60000
rect 20720 59600 20776 60000
rect 21168 59600 21224 60000
rect 21616 59600 21672 60000
rect 22064 59600 22120 60000
rect 22512 59600 22568 60000
rect 22960 59600 23016 60000
rect 23408 59600 23464 60000
rect 23856 59600 23912 60000
rect 24304 59600 24360 60000
rect 24752 59600 24808 60000
rect 25200 59600 25256 60000
rect 25648 59600 25704 60000
rect 26096 59600 26152 60000
rect 26544 59600 26600 60000
rect 26992 59600 27048 60000
rect 27440 59600 27496 60000
rect 27888 59600 27944 60000
rect 28336 59600 28392 60000
rect 28784 59600 28840 60000
rect 29232 59600 29288 60000
rect 29680 59600 29736 60000
rect 30128 59600 30184 60000
rect 30576 59600 30632 60000
rect 31024 59600 31080 60000
rect 31472 59600 31528 60000
rect 31920 59600 31976 60000
rect 32368 59600 32424 60000
rect 32816 59600 32872 60000
rect 33264 59600 33320 60000
rect 33712 59600 33768 60000
rect 34160 59600 34216 60000
rect 34608 59600 34664 60000
rect 35056 59600 35112 60000
rect 35504 59600 35560 60000
rect 35952 59600 36008 60000
rect 36400 59600 36456 60000
rect 36848 59600 36904 60000
rect 37296 59600 37352 60000
rect 37744 59600 37800 60000
rect 38192 59600 38248 60000
rect 38640 59600 38696 60000
rect 39088 59600 39144 60000
rect 39536 59600 39592 60000
rect 39984 59600 40040 60000
rect 40432 59600 40488 60000
rect 40880 59600 40936 60000
rect 41328 59600 41384 60000
rect 41776 59600 41832 60000
rect 42224 59600 42280 60000
rect 42672 59600 42728 60000
rect 43120 59600 43176 60000
rect 43568 59600 43624 60000
rect 44016 59600 44072 60000
rect 44464 59600 44520 60000
rect 44912 59600 44968 60000
rect 45360 59600 45416 60000
rect 45808 59600 45864 60000
rect 46256 59600 46312 60000
rect 46704 59600 46760 60000
rect 47152 59600 47208 60000
rect 47600 59600 47656 60000
rect 48048 59600 48104 60000
rect 48496 59600 48552 60000
rect 48944 59600 49000 60000
rect 49392 59600 49448 60000
rect 49840 59600 49896 60000
rect 50288 59600 50344 60000
rect 50736 59600 50792 60000
rect 51184 59600 51240 60000
rect 51632 59600 51688 60000
rect 52080 59600 52136 60000
rect 52528 59600 52584 60000
rect 52976 59600 53032 60000
rect 53424 59600 53480 60000
rect 53872 59600 53928 60000
rect 54320 59600 54376 60000
rect 54768 59600 54824 60000
rect 55216 59600 55272 60000
rect 55664 59600 55720 60000
rect 56112 59600 56168 60000
rect 56560 59600 56616 60000
rect 57008 59600 57064 60000
rect 57456 59600 57512 60000
rect 57904 59600 57960 60000
rect 58352 59600 58408 60000
rect 58800 59600 58856 60000
rect 59248 59600 59304 60000
rect 59696 59600 59752 60000
rect 60144 59600 60200 60000
rect 60592 59600 60648 60000
rect 2576 0 2632 400
rect 3024 0 3080 400
rect 3472 0 3528 400
rect 3920 0 3976 400
rect 4368 0 4424 400
rect 4816 0 4872 400
rect 5264 0 5320 400
rect 5712 0 5768 400
rect 6160 0 6216 400
rect 6608 0 6664 400
rect 7056 0 7112 400
rect 7504 0 7560 400
rect 7952 0 8008 400
rect 8400 0 8456 400
rect 8848 0 8904 400
rect 9296 0 9352 400
rect 9744 0 9800 400
rect 10192 0 10248 400
rect 10640 0 10696 400
rect 11088 0 11144 400
rect 11536 0 11592 400
rect 11984 0 12040 400
rect 12432 0 12488 400
rect 12880 0 12936 400
rect 13328 0 13384 400
rect 13776 0 13832 400
rect 14224 0 14280 400
rect 14672 0 14728 400
rect 15120 0 15176 400
rect 15568 0 15624 400
rect 16016 0 16072 400
rect 16464 0 16520 400
rect 16912 0 16968 400
rect 17360 0 17416 400
rect 17808 0 17864 400
rect 18256 0 18312 400
rect 18704 0 18760 400
rect 19152 0 19208 400
rect 19600 0 19656 400
rect 20048 0 20104 400
rect 20496 0 20552 400
rect 20944 0 21000 400
rect 21392 0 21448 400
rect 21840 0 21896 400
rect 22288 0 22344 400
rect 22736 0 22792 400
rect 23184 0 23240 400
rect 23632 0 23688 400
rect 24080 0 24136 400
rect 24528 0 24584 400
rect 24976 0 25032 400
rect 25424 0 25480 400
rect 25872 0 25928 400
rect 26320 0 26376 400
rect 26768 0 26824 400
rect 27216 0 27272 400
rect 27664 0 27720 400
rect 28112 0 28168 400
rect 28560 0 28616 400
rect 29008 0 29064 400
rect 29456 0 29512 400
rect 29904 0 29960 400
rect 30352 0 30408 400
rect 30800 0 30856 400
rect 31248 0 31304 400
rect 31696 0 31752 400
rect 32144 0 32200 400
rect 32592 0 32648 400
rect 33040 0 33096 400
rect 33488 0 33544 400
rect 33936 0 33992 400
rect 34384 0 34440 400
rect 34832 0 34888 400
rect 35280 0 35336 400
rect 35728 0 35784 400
rect 36176 0 36232 400
rect 36624 0 36680 400
rect 37072 0 37128 400
rect 37520 0 37576 400
rect 37968 0 38024 400
rect 38416 0 38472 400
rect 38864 0 38920 400
rect 39312 0 39368 400
rect 39760 0 39816 400
rect 40208 0 40264 400
rect 40656 0 40712 400
rect 41104 0 41160 400
rect 41552 0 41608 400
rect 42000 0 42056 400
rect 42448 0 42504 400
rect 42896 0 42952 400
rect 43344 0 43400 400
rect 43792 0 43848 400
rect 44240 0 44296 400
rect 44688 0 44744 400
rect 45136 0 45192 400
rect 45584 0 45640 400
rect 46032 0 46088 400
rect 46480 0 46536 400
rect 46928 0 46984 400
rect 47376 0 47432 400
rect 47824 0 47880 400
rect 48272 0 48328 400
rect 48720 0 48776 400
rect 49168 0 49224 400
rect 49616 0 49672 400
rect 50064 0 50120 400
rect 50512 0 50568 400
rect 50960 0 51016 400
rect 51408 0 51464 400
rect 51856 0 51912 400
rect 52304 0 52360 400
rect 52752 0 52808 400
rect 53200 0 53256 400
rect 53648 0 53704 400
rect 54096 0 54152 400
rect 54544 0 54600 400
rect 54992 0 55048 400
rect 55440 0 55496 400
rect 55888 0 55944 400
rect 56336 0 56392 400
rect 56784 0 56840 400
rect 57232 0 57288 400
rect 57680 0 57736 400
rect 58128 0 58184 400
rect 58576 0 58632 400
rect 59024 0 59080 400
rect 59472 0 59528 400
rect 59920 0 59976 400
rect 60368 0 60424 400
rect 60816 0 60872 400
rect 61264 0 61320 400
rect 61712 0 61768 400
rect 62160 0 62216 400
<< obsm2 >>
rect 630 59570 4114 59682
rect 4230 59570 4562 59682
rect 4678 59570 5010 59682
rect 5126 59570 5458 59682
rect 5574 59570 5906 59682
rect 6022 59570 6354 59682
rect 6470 59570 6802 59682
rect 6918 59570 7250 59682
rect 7366 59570 7698 59682
rect 7814 59570 8146 59682
rect 8262 59570 8594 59682
rect 8710 59570 9042 59682
rect 9158 59570 9490 59682
rect 9606 59570 9938 59682
rect 10054 59570 10386 59682
rect 10502 59570 10834 59682
rect 10950 59570 11282 59682
rect 11398 59570 11730 59682
rect 11846 59570 12178 59682
rect 12294 59570 12626 59682
rect 12742 59570 13074 59682
rect 13190 59570 13522 59682
rect 13638 59570 13970 59682
rect 14086 59570 14418 59682
rect 14534 59570 14866 59682
rect 14982 59570 15314 59682
rect 15430 59570 15762 59682
rect 15878 59570 16210 59682
rect 16326 59570 16658 59682
rect 16774 59570 17106 59682
rect 17222 59570 17554 59682
rect 17670 59570 18002 59682
rect 18118 59570 18450 59682
rect 18566 59570 18898 59682
rect 19014 59570 19346 59682
rect 19462 59570 19794 59682
rect 19910 59570 20242 59682
rect 20358 59570 20690 59682
rect 20806 59570 21138 59682
rect 21254 59570 21586 59682
rect 21702 59570 22034 59682
rect 22150 59570 22482 59682
rect 22598 59570 22930 59682
rect 23046 59570 23378 59682
rect 23494 59570 23826 59682
rect 23942 59570 24274 59682
rect 24390 59570 24722 59682
rect 24838 59570 25170 59682
rect 25286 59570 25618 59682
rect 25734 59570 26066 59682
rect 26182 59570 26514 59682
rect 26630 59570 26962 59682
rect 27078 59570 27410 59682
rect 27526 59570 27858 59682
rect 27974 59570 28306 59682
rect 28422 59570 28754 59682
rect 28870 59570 29202 59682
rect 29318 59570 29650 59682
rect 29766 59570 30098 59682
rect 30214 59570 30546 59682
rect 30662 59570 30994 59682
rect 31110 59570 31442 59682
rect 31558 59570 31890 59682
rect 32006 59570 32338 59682
rect 32454 59570 32786 59682
rect 32902 59570 33234 59682
rect 33350 59570 33682 59682
rect 33798 59570 34130 59682
rect 34246 59570 34578 59682
rect 34694 59570 35026 59682
rect 35142 59570 35474 59682
rect 35590 59570 35922 59682
rect 36038 59570 36370 59682
rect 36486 59570 36818 59682
rect 36934 59570 37266 59682
rect 37382 59570 37714 59682
rect 37830 59570 38162 59682
rect 38278 59570 38610 59682
rect 38726 59570 39058 59682
rect 39174 59570 39506 59682
rect 39622 59570 39954 59682
rect 40070 59570 40402 59682
rect 40518 59570 40850 59682
rect 40966 59570 41298 59682
rect 41414 59570 41746 59682
rect 41862 59570 42194 59682
rect 42310 59570 42642 59682
rect 42758 59570 43090 59682
rect 43206 59570 43538 59682
rect 43654 59570 43986 59682
rect 44102 59570 44434 59682
rect 44550 59570 44882 59682
rect 44998 59570 45330 59682
rect 45446 59570 45778 59682
rect 45894 59570 46226 59682
rect 46342 59570 46674 59682
rect 46790 59570 47122 59682
rect 47238 59570 47570 59682
rect 47686 59570 48018 59682
rect 48134 59570 48466 59682
rect 48582 59570 48914 59682
rect 49030 59570 49362 59682
rect 49478 59570 49810 59682
rect 49926 59570 50258 59682
rect 50374 59570 50706 59682
rect 50822 59570 51154 59682
rect 51270 59570 51602 59682
rect 51718 59570 52050 59682
rect 52166 59570 52498 59682
rect 52614 59570 52946 59682
rect 53062 59570 53394 59682
rect 53510 59570 53842 59682
rect 53958 59570 54290 59682
rect 54406 59570 54738 59682
rect 54854 59570 55186 59682
rect 55302 59570 55634 59682
rect 55750 59570 56082 59682
rect 56198 59570 56530 59682
rect 56646 59570 56978 59682
rect 57094 59570 57426 59682
rect 57542 59570 57874 59682
rect 57990 59570 58322 59682
rect 58438 59570 58770 59682
rect 58886 59570 59218 59682
rect 59334 59570 59666 59682
rect 59782 59570 60114 59682
rect 60230 59570 60562 59682
rect 60678 59570 64498 59682
rect 630 430 64498 59570
rect 630 350 2546 430
rect 2662 350 2994 430
rect 3110 350 3442 430
rect 3558 350 3890 430
rect 4006 350 4338 430
rect 4454 350 4786 430
rect 4902 350 5234 430
rect 5350 350 5682 430
rect 5798 350 6130 430
rect 6246 350 6578 430
rect 6694 350 7026 430
rect 7142 350 7474 430
rect 7590 350 7922 430
rect 8038 350 8370 430
rect 8486 350 8818 430
rect 8934 350 9266 430
rect 9382 350 9714 430
rect 9830 350 10162 430
rect 10278 350 10610 430
rect 10726 350 11058 430
rect 11174 350 11506 430
rect 11622 350 11954 430
rect 12070 350 12402 430
rect 12518 350 12850 430
rect 12966 350 13298 430
rect 13414 350 13746 430
rect 13862 350 14194 430
rect 14310 350 14642 430
rect 14758 350 15090 430
rect 15206 350 15538 430
rect 15654 350 15986 430
rect 16102 350 16434 430
rect 16550 350 16882 430
rect 16998 350 17330 430
rect 17446 350 17778 430
rect 17894 350 18226 430
rect 18342 350 18674 430
rect 18790 350 19122 430
rect 19238 350 19570 430
rect 19686 350 20018 430
rect 20134 350 20466 430
rect 20582 350 20914 430
rect 21030 350 21362 430
rect 21478 350 21810 430
rect 21926 350 22258 430
rect 22374 350 22706 430
rect 22822 350 23154 430
rect 23270 350 23602 430
rect 23718 350 24050 430
rect 24166 350 24498 430
rect 24614 350 24946 430
rect 25062 350 25394 430
rect 25510 350 25842 430
rect 25958 350 26290 430
rect 26406 350 26738 430
rect 26854 350 27186 430
rect 27302 350 27634 430
rect 27750 350 28082 430
rect 28198 350 28530 430
rect 28646 350 28978 430
rect 29094 350 29426 430
rect 29542 350 29874 430
rect 29990 350 30322 430
rect 30438 350 30770 430
rect 30886 350 31218 430
rect 31334 350 31666 430
rect 31782 350 32114 430
rect 32230 350 32562 430
rect 32678 350 33010 430
rect 33126 350 33458 430
rect 33574 350 33906 430
rect 34022 350 34354 430
rect 34470 350 34802 430
rect 34918 350 35250 430
rect 35366 350 35698 430
rect 35814 350 36146 430
rect 36262 350 36594 430
rect 36710 350 37042 430
rect 37158 350 37490 430
rect 37606 350 37938 430
rect 38054 350 38386 430
rect 38502 350 38834 430
rect 38950 350 39282 430
rect 39398 350 39730 430
rect 39846 350 40178 430
rect 40294 350 40626 430
rect 40742 350 41074 430
rect 41190 350 41522 430
rect 41638 350 41970 430
rect 42086 350 42418 430
rect 42534 350 42866 430
rect 42982 350 43314 430
rect 43430 350 43762 430
rect 43878 350 44210 430
rect 44326 350 44658 430
rect 44774 350 45106 430
rect 45222 350 45554 430
rect 45670 350 46002 430
rect 46118 350 46450 430
rect 46566 350 46898 430
rect 47014 350 47346 430
rect 47462 350 47794 430
rect 47910 350 48242 430
rect 48358 350 48690 430
rect 48806 350 49138 430
rect 49254 350 49586 430
rect 49702 350 50034 430
rect 50150 350 50482 430
rect 50598 350 50930 430
rect 51046 350 51378 430
rect 51494 350 51826 430
rect 51942 350 52274 430
rect 52390 350 52722 430
rect 52838 350 53170 430
rect 53286 350 53618 430
rect 53734 350 54066 430
rect 54182 350 54514 430
rect 54630 350 54962 430
rect 55078 350 55410 430
rect 55526 350 55858 430
rect 55974 350 56306 430
rect 56422 350 56754 430
rect 56870 350 57202 430
rect 57318 350 57650 430
rect 57766 350 58098 430
rect 58214 350 58546 430
rect 58662 350 58994 430
rect 59110 350 59442 430
rect 59558 350 59890 430
rect 60006 350 60338 430
rect 60454 350 60786 430
rect 60902 350 61234 430
rect 61350 350 61682 430
rect 61798 350 62130 430
rect 62246 350 64498 430
<< metal3 >>
rect 0 56560 400 56616
rect 64600 56112 65000 56168
rect 0 56000 400 56056
rect 64600 55664 65000 55720
rect 0 55440 400 55496
rect 64600 55216 65000 55272
rect 0 54880 400 54936
rect 64600 54768 65000 54824
rect 0 54320 400 54376
rect 64600 54320 65000 54376
rect 64600 53872 65000 53928
rect 0 53760 400 53816
rect 64600 53424 65000 53480
rect 0 53200 400 53256
rect 64600 52976 65000 53032
rect 0 52640 400 52696
rect 64600 52528 65000 52584
rect 0 52080 400 52136
rect 64600 52080 65000 52136
rect 64600 51632 65000 51688
rect 0 51520 400 51576
rect 64600 51184 65000 51240
rect 0 50960 400 51016
rect 64600 50736 65000 50792
rect 0 50400 400 50456
rect 64600 50288 65000 50344
rect 0 49840 400 49896
rect 64600 49840 65000 49896
rect 64600 49392 65000 49448
rect 0 49280 400 49336
rect 64600 48944 65000 49000
rect 0 48720 400 48776
rect 64600 48496 65000 48552
rect 0 48160 400 48216
rect 64600 48048 65000 48104
rect 0 47600 400 47656
rect 64600 47600 65000 47656
rect 64600 47152 65000 47208
rect 0 47040 400 47096
rect 64600 46704 65000 46760
rect 0 46480 400 46536
rect 64600 46256 65000 46312
rect 0 45920 400 45976
rect 64600 45808 65000 45864
rect 0 45360 400 45416
rect 64600 45360 65000 45416
rect 64600 44912 65000 44968
rect 0 44800 400 44856
rect 64600 44464 65000 44520
rect 0 44240 400 44296
rect 64600 44016 65000 44072
rect 0 43680 400 43736
rect 64600 43568 65000 43624
rect 0 43120 400 43176
rect 64600 43120 65000 43176
rect 64600 42672 65000 42728
rect 0 42560 400 42616
rect 64600 42224 65000 42280
rect 0 42000 400 42056
rect 64600 41776 65000 41832
rect 0 41440 400 41496
rect 64600 41328 65000 41384
rect 0 40880 400 40936
rect 64600 40880 65000 40936
rect 64600 40432 65000 40488
rect 0 40320 400 40376
rect 64600 39984 65000 40040
rect 0 39760 400 39816
rect 64600 39536 65000 39592
rect 0 39200 400 39256
rect 64600 39088 65000 39144
rect 0 38640 400 38696
rect 64600 38640 65000 38696
rect 64600 38192 65000 38248
rect 0 38080 400 38136
rect 64600 37744 65000 37800
rect 0 37520 400 37576
rect 64600 37296 65000 37352
rect 0 36960 400 37016
rect 64600 36848 65000 36904
rect 0 36400 400 36456
rect 64600 36400 65000 36456
rect 64600 35952 65000 36008
rect 0 35840 400 35896
rect 64600 35504 65000 35560
rect 0 35280 400 35336
rect 64600 35056 65000 35112
rect 0 34720 400 34776
rect 64600 34608 65000 34664
rect 0 34160 400 34216
rect 64600 34160 65000 34216
rect 64600 33712 65000 33768
rect 0 33600 400 33656
rect 64600 33264 65000 33320
rect 0 33040 400 33096
rect 64600 32816 65000 32872
rect 0 32480 400 32536
rect 64600 32368 65000 32424
rect 0 31920 400 31976
rect 64600 31920 65000 31976
rect 64600 31472 65000 31528
rect 0 31360 400 31416
rect 64600 31024 65000 31080
rect 0 30800 400 30856
rect 64600 30576 65000 30632
rect 0 30240 400 30296
rect 64600 30128 65000 30184
rect 0 29680 400 29736
rect 64600 29680 65000 29736
rect 64600 29232 65000 29288
rect 0 29120 400 29176
rect 64600 28784 65000 28840
rect 0 28560 400 28616
rect 64600 28336 65000 28392
rect 0 28000 400 28056
rect 64600 27888 65000 27944
rect 0 27440 400 27496
rect 64600 27440 65000 27496
rect 64600 26992 65000 27048
rect 0 26880 400 26936
rect 64600 26544 65000 26600
rect 0 26320 400 26376
rect 64600 26096 65000 26152
rect 0 25760 400 25816
rect 64600 25648 65000 25704
rect 0 25200 400 25256
rect 64600 25200 65000 25256
rect 64600 24752 65000 24808
rect 0 24640 400 24696
rect 64600 24304 65000 24360
rect 0 24080 400 24136
rect 64600 23856 65000 23912
rect 0 23520 400 23576
rect 64600 23408 65000 23464
rect 0 22960 400 23016
rect 64600 22960 65000 23016
rect 64600 22512 65000 22568
rect 0 22400 400 22456
rect 64600 22064 65000 22120
rect 0 21840 400 21896
rect 64600 21616 65000 21672
rect 0 21280 400 21336
rect 64600 21168 65000 21224
rect 0 20720 400 20776
rect 64600 20720 65000 20776
rect 64600 20272 65000 20328
rect 0 20160 400 20216
rect 64600 19824 65000 19880
rect 0 19600 400 19656
rect 64600 19376 65000 19432
rect 0 19040 400 19096
rect 64600 18928 65000 18984
rect 0 18480 400 18536
rect 64600 18480 65000 18536
rect 64600 18032 65000 18088
rect 0 17920 400 17976
rect 64600 17584 65000 17640
rect 0 17360 400 17416
rect 64600 17136 65000 17192
rect 0 16800 400 16856
rect 64600 16688 65000 16744
rect 0 16240 400 16296
rect 64600 16240 65000 16296
rect 64600 15792 65000 15848
rect 0 15680 400 15736
rect 64600 15344 65000 15400
rect 0 15120 400 15176
rect 64600 14896 65000 14952
rect 0 14560 400 14616
rect 64600 14448 65000 14504
rect 0 14000 400 14056
rect 64600 14000 65000 14056
rect 64600 13552 65000 13608
rect 0 13440 400 13496
rect 64600 13104 65000 13160
rect 0 12880 400 12936
rect 64600 12656 65000 12712
rect 0 12320 400 12376
rect 64600 12208 65000 12264
rect 0 11760 400 11816
rect 64600 11760 65000 11816
rect 64600 11312 65000 11368
rect 0 11200 400 11256
rect 64600 10864 65000 10920
rect 0 10640 400 10696
rect 64600 10416 65000 10472
rect 0 10080 400 10136
rect 64600 9968 65000 10024
rect 0 9520 400 9576
rect 64600 9520 65000 9576
rect 64600 9072 65000 9128
rect 0 8960 400 9016
rect 64600 8624 65000 8680
rect 0 8400 400 8456
rect 64600 8176 65000 8232
rect 0 7840 400 7896
rect 64600 7728 65000 7784
rect 0 7280 400 7336
rect 64600 7280 65000 7336
rect 64600 6832 65000 6888
rect 0 6720 400 6776
rect 64600 6384 65000 6440
rect 0 6160 400 6216
rect 64600 5936 65000 5992
rect 0 5600 400 5656
rect 64600 5488 65000 5544
rect 0 5040 400 5096
rect 64600 5040 65000 5096
rect 64600 4592 65000 4648
rect 0 4480 400 4536
rect 64600 4144 65000 4200
rect 0 3920 400 3976
rect 64600 3696 65000 3752
rect 0 3360 400 3416
<< obsm3 >>
rect 400 56646 64666 59066
rect 430 56530 64666 56646
rect 400 56198 64666 56530
rect 400 56086 64570 56198
rect 430 56082 64570 56086
rect 430 55970 64666 56082
rect 400 55750 64666 55970
rect 400 55634 64570 55750
rect 400 55526 64666 55634
rect 430 55410 64666 55526
rect 400 55302 64666 55410
rect 400 55186 64570 55302
rect 400 54966 64666 55186
rect 430 54854 64666 54966
rect 430 54850 64570 54854
rect 400 54738 64570 54850
rect 400 54406 64666 54738
rect 430 54290 64570 54406
rect 400 53958 64666 54290
rect 400 53846 64570 53958
rect 430 53842 64570 53846
rect 430 53730 64666 53842
rect 400 53510 64666 53730
rect 400 53394 64570 53510
rect 400 53286 64666 53394
rect 430 53170 64666 53286
rect 400 53062 64666 53170
rect 400 52946 64570 53062
rect 400 52726 64666 52946
rect 430 52614 64666 52726
rect 430 52610 64570 52614
rect 400 52498 64570 52610
rect 400 52166 64666 52498
rect 430 52050 64570 52166
rect 400 51718 64666 52050
rect 400 51606 64570 51718
rect 430 51602 64570 51606
rect 430 51490 64666 51602
rect 400 51270 64666 51490
rect 400 51154 64570 51270
rect 400 51046 64666 51154
rect 430 50930 64666 51046
rect 400 50822 64666 50930
rect 400 50706 64570 50822
rect 400 50486 64666 50706
rect 430 50374 64666 50486
rect 430 50370 64570 50374
rect 400 50258 64570 50370
rect 400 49926 64666 50258
rect 430 49810 64570 49926
rect 400 49478 64666 49810
rect 400 49366 64570 49478
rect 430 49362 64570 49366
rect 430 49250 64666 49362
rect 400 49030 64666 49250
rect 400 48914 64570 49030
rect 400 48806 64666 48914
rect 430 48690 64666 48806
rect 400 48582 64666 48690
rect 400 48466 64570 48582
rect 400 48246 64666 48466
rect 430 48134 64666 48246
rect 430 48130 64570 48134
rect 400 48018 64570 48130
rect 400 47686 64666 48018
rect 430 47570 64570 47686
rect 400 47238 64666 47570
rect 400 47126 64570 47238
rect 430 47122 64570 47126
rect 430 47010 64666 47122
rect 400 46790 64666 47010
rect 400 46674 64570 46790
rect 400 46566 64666 46674
rect 430 46450 64666 46566
rect 400 46342 64666 46450
rect 400 46226 64570 46342
rect 400 46006 64666 46226
rect 430 45894 64666 46006
rect 430 45890 64570 45894
rect 400 45778 64570 45890
rect 400 45446 64666 45778
rect 430 45330 64570 45446
rect 400 44998 64666 45330
rect 400 44886 64570 44998
rect 430 44882 64570 44886
rect 430 44770 64666 44882
rect 400 44550 64666 44770
rect 400 44434 64570 44550
rect 400 44326 64666 44434
rect 430 44210 64666 44326
rect 400 44102 64666 44210
rect 400 43986 64570 44102
rect 400 43766 64666 43986
rect 430 43654 64666 43766
rect 430 43650 64570 43654
rect 400 43538 64570 43650
rect 400 43206 64666 43538
rect 430 43090 64570 43206
rect 400 42758 64666 43090
rect 400 42646 64570 42758
rect 430 42642 64570 42646
rect 430 42530 64666 42642
rect 400 42310 64666 42530
rect 400 42194 64570 42310
rect 400 42086 64666 42194
rect 430 41970 64666 42086
rect 400 41862 64666 41970
rect 400 41746 64570 41862
rect 400 41526 64666 41746
rect 430 41414 64666 41526
rect 430 41410 64570 41414
rect 400 41298 64570 41410
rect 400 40966 64666 41298
rect 430 40850 64570 40966
rect 400 40518 64666 40850
rect 400 40406 64570 40518
rect 430 40402 64570 40406
rect 430 40290 64666 40402
rect 400 40070 64666 40290
rect 400 39954 64570 40070
rect 400 39846 64666 39954
rect 430 39730 64666 39846
rect 400 39622 64666 39730
rect 400 39506 64570 39622
rect 400 39286 64666 39506
rect 430 39174 64666 39286
rect 430 39170 64570 39174
rect 400 39058 64570 39170
rect 400 38726 64666 39058
rect 430 38610 64570 38726
rect 400 38278 64666 38610
rect 400 38166 64570 38278
rect 430 38162 64570 38166
rect 430 38050 64666 38162
rect 400 37830 64666 38050
rect 400 37714 64570 37830
rect 400 37606 64666 37714
rect 430 37490 64666 37606
rect 400 37382 64666 37490
rect 400 37266 64570 37382
rect 400 37046 64666 37266
rect 430 36934 64666 37046
rect 430 36930 64570 36934
rect 400 36818 64570 36930
rect 400 36486 64666 36818
rect 430 36370 64570 36486
rect 400 36038 64666 36370
rect 400 35926 64570 36038
rect 430 35922 64570 35926
rect 430 35810 64666 35922
rect 400 35590 64666 35810
rect 400 35474 64570 35590
rect 400 35366 64666 35474
rect 430 35250 64666 35366
rect 400 35142 64666 35250
rect 400 35026 64570 35142
rect 400 34806 64666 35026
rect 430 34694 64666 34806
rect 430 34690 64570 34694
rect 400 34578 64570 34690
rect 400 34246 64666 34578
rect 430 34130 64570 34246
rect 400 33798 64666 34130
rect 400 33686 64570 33798
rect 430 33682 64570 33686
rect 430 33570 64666 33682
rect 400 33350 64666 33570
rect 400 33234 64570 33350
rect 400 33126 64666 33234
rect 430 33010 64666 33126
rect 400 32902 64666 33010
rect 400 32786 64570 32902
rect 400 32566 64666 32786
rect 430 32454 64666 32566
rect 430 32450 64570 32454
rect 400 32338 64570 32450
rect 400 32006 64666 32338
rect 430 31890 64570 32006
rect 400 31558 64666 31890
rect 400 31446 64570 31558
rect 430 31442 64570 31446
rect 430 31330 64666 31442
rect 400 31110 64666 31330
rect 400 30994 64570 31110
rect 400 30886 64666 30994
rect 430 30770 64666 30886
rect 400 30662 64666 30770
rect 400 30546 64570 30662
rect 400 30326 64666 30546
rect 430 30214 64666 30326
rect 430 30210 64570 30214
rect 400 30098 64570 30210
rect 400 29766 64666 30098
rect 430 29650 64570 29766
rect 400 29318 64666 29650
rect 400 29206 64570 29318
rect 430 29202 64570 29206
rect 430 29090 64666 29202
rect 400 28870 64666 29090
rect 400 28754 64570 28870
rect 400 28646 64666 28754
rect 430 28530 64666 28646
rect 400 28422 64666 28530
rect 400 28306 64570 28422
rect 400 28086 64666 28306
rect 430 27974 64666 28086
rect 430 27970 64570 27974
rect 400 27858 64570 27970
rect 400 27526 64666 27858
rect 430 27410 64570 27526
rect 400 27078 64666 27410
rect 400 26966 64570 27078
rect 430 26962 64570 26966
rect 430 26850 64666 26962
rect 400 26630 64666 26850
rect 400 26514 64570 26630
rect 400 26406 64666 26514
rect 430 26290 64666 26406
rect 400 26182 64666 26290
rect 400 26066 64570 26182
rect 400 25846 64666 26066
rect 430 25734 64666 25846
rect 430 25730 64570 25734
rect 400 25618 64570 25730
rect 400 25286 64666 25618
rect 430 25170 64570 25286
rect 400 24838 64666 25170
rect 400 24726 64570 24838
rect 430 24722 64570 24726
rect 430 24610 64666 24722
rect 400 24390 64666 24610
rect 400 24274 64570 24390
rect 400 24166 64666 24274
rect 430 24050 64666 24166
rect 400 23942 64666 24050
rect 400 23826 64570 23942
rect 400 23606 64666 23826
rect 430 23494 64666 23606
rect 430 23490 64570 23494
rect 400 23378 64570 23490
rect 400 23046 64666 23378
rect 430 22930 64570 23046
rect 400 22598 64666 22930
rect 400 22486 64570 22598
rect 430 22482 64570 22486
rect 430 22370 64666 22482
rect 400 22150 64666 22370
rect 400 22034 64570 22150
rect 400 21926 64666 22034
rect 430 21810 64666 21926
rect 400 21702 64666 21810
rect 400 21586 64570 21702
rect 400 21366 64666 21586
rect 430 21254 64666 21366
rect 430 21250 64570 21254
rect 400 21138 64570 21250
rect 400 20806 64666 21138
rect 430 20690 64570 20806
rect 400 20358 64666 20690
rect 400 20246 64570 20358
rect 430 20242 64570 20246
rect 430 20130 64666 20242
rect 400 19910 64666 20130
rect 400 19794 64570 19910
rect 400 19686 64666 19794
rect 430 19570 64666 19686
rect 400 19462 64666 19570
rect 400 19346 64570 19462
rect 400 19126 64666 19346
rect 430 19014 64666 19126
rect 430 19010 64570 19014
rect 400 18898 64570 19010
rect 400 18566 64666 18898
rect 430 18450 64570 18566
rect 400 18118 64666 18450
rect 400 18006 64570 18118
rect 430 18002 64570 18006
rect 430 17890 64666 18002
rect 400 17670 64666 17890
rect 400 17554 64570 17670
rect 400 17446 64666 17554
rect 430 17330 64666 17446
rect 400 17222 64666 17330
rect 400 17106 64570 17222
rect 400 16886 64666 17106
rect 430 16774 64666 16886
rect 430 16770 64570 16774
rect 400 16658 64570 16770
rect 400 16326 64666 16658
rect 430 16210 64570 16326
rect 400 15878 64666 16210
rect 400 15766 64570 15878
rect 430 15762 64570 15766
rect 430 15650 64666 15762
rect 400 15430 64666 15650
rect 400 15314 64570 15430
rect 400 15206 64666 15314
rect 430 15090 64666 15206
rect 400 14982 64666 15090
rect 400 14866 64570 14982
rect 400 14646 64666 14866
rect 430 14534 64666 14646
rect 430 14530 64570 14534
rect 400 14418 64570 14530
rect 400 14086 64666 14418
rect 430 13970 64570 14086
rect 400 13638 64666 13970
rect 400 13526 64570 13638
rect 430 13522 64570 13526
rect 430 13410 64666 13522
rect 400 13190 64666 13410
rect 400 13074 64570 13190
rect 400 12966 64666 13074
rect 430 12850 64666 12966
rect 400 12742 64666 12850
rect 400 12626 64570 12742
rect 400 12406 64666 12626
rect 430 12294 64666 12406
rect 430 12290 64570 12294
rect 400 12178 64570 12290
rect 400 11846 64666 12178
rect 430 11730 64570 11846
rect 400 11398 64666 11730
rect 400 11286 64570 11398
rect 430 11282 64570 11286
rect 430 11170 64666 11282
rect 400 10950 64666 11170
rect 400 10834 64570 10950
rect 400 10726 64666 10834
rect 430 10610 64666 10726
rect 400 10502 64666 10610
rect 400 10386 64570 10502
rect 400 10166 64666 10386
rect 430 10054 64666 10166
rect 430 10050 64570 10054
rect 400 9938 64570 10050
rect 400 9606 64666 9938
rect 430 9490 64570 9606
rect 400 9158 64666 9490
rect 400 9046 64570 9158
rect 430 9042 64570 9046
rect 430 8930 64666 9042
rect 400 8710 64666 8930
rect 400 8594 64570 8710
rect 400 8486 64666 8594
rect 430 8370 64666 8486
rect 400 8262 64666 8370
rect 400 8146 64570 8262
rect 400 7926 64666 8146
rect 430 7814 64666 7926
rect 430 7810 64570 7814
rect 400 7698 64570 7810
rect 400 7366 64666 7698
rect 430 7250 64570 7366
rect 400 6918 64666 7250
rect 400 6806 64570 6918
rect 430 6802 64570 6806
rect 430 6690 64666 6802
rect 400 6470 64666 6690
rect 400 6354 64570 6470
rect 400 6246 64666 6354
rect 430 6130 64666 6246
rect 400 6022 64666 6130
rect 400 5906 64570 6022
rect 400 5686 64666 5906
rect 430 5574 64666 5686
rect 430 5570 64570 5574
rect 400 5458 64570 5570
rect 400 5126 64666 5458
rect 430 5010 64570 5126
rect 400 4678 64666 5010
rect 400 4566 64570 4678
rect 430 4562 64570 4566
rect 430 4450 64666 4562
rect 400 4230 64666 4450
rect 400 4114 64570 4230
rect 400 4006 64666 4114
rect 430 3890 64666 4006
rect 400 3782 64666 3890
rect 400 3666 64570 3782
rect 400 3446 64666 3666
rect 430 3330 64666 3446
rect 400 630 64666 3330
<< metal4 >>
rect 2224 1538 2384 58438
rect 9904 1538 10064 58438
rect 17584 1538 17744 58438
rect 25264 1538 25424 58438
rect 32944 1538 33104 58438
rect 40624 1538 40784 58438
rect 48304 1538 48464 58438
rect 55984 1538 56144 58438
rect 63664 1538 63824 58438
<< obsm4 >>
rect 7406 1508 9874 58287
rect 10094 1508 17554 58287
rect 17774 1508 25234 58287
rect 25454 1508 32914 58287
rect 33134 1508 40594 58287
rect 40814 1508 48274 58287
rect 48494 1508 55954 58287
rect 56174 1508 63602 58287
rect 7406 1129 63602 1508
<< labels >>
rlabel metal2 s 48496 59600 48552 60000 6 ay8913_do[0]
port 1 nsew signal input
rlabel metal2 s 52976 59600 53032 60000 6 ay8913_do[10]
port 2 nsew signal input
rlabel metal2 s 53424 59600 53480 60000 6 ay8913_do[11]
port 3 nsew signal input
rlabel metal2 s 53872 59600 53928 60000 6 ay8913_do[12]
port 4 nsew signal input
rlabel metal2 s 54320 59600 54376 60000 6 ay8913_do[13]
port 5 nsew signal input
rlabel metal2 s 54768 59600 54824 60000 6 ay8913_do[14]
port 6 nsew signal input
rlabel metal2 s 55216 59600 55272 60000 6 ay8913_do[15]
port 7 nsew signal input
rlabel metal2 s 55664 59600 55720 60000 6 ay8913_do[16]
port 8 nsew signal input
rlabel metal2 s 56112 59600 56168 60000 6 ay8913_do[17]
port 9 nsew signal input
rlabel metal2 s 56560 59600 56616 60000 6 ay8913_do[18]
port 10 nsew signal input
rlabel metal2 s 57008 59600 57064 60000 6 ay8913_do[19]
port 11 nsew signal input
rlabel metal2 s 48944 59600 49000 60000 6 ay8913_do[1]
port 12 nsew signal input
rlabel metal2 s 57456 59600 57512 60000 6 ay8913_do[20]
port 13 nsew signal input
rlabel metal2 s 57904 59600 57960 60000 6 ay8913_do[21]
port 14 nsew signal input
rlabel metal2 s 58352 59600 58408 60000 6 ay8913_do[22]
port 15 nsew signal input
rlabel metal2 s 58800 59600 58856 60000 6 ay8913_do[23]
port 16 nsew signal input
rlabel metal2 s 59248 59600 59304 60000 6 ay8913_do[24]
port 17 nsew signal input
rlabel metal2 s 59696 59600 59752 60000 6 ay8913_do[25]
port 18 nsew signal input
rlabel metal2 s 60144 59600 60200 60000 6 ay8913_do[26]
port 19 nsew signal input
rlabel metal2 s 60592 59600 60648 60000 6 ay8913_do[27]
port 20 nsew signal input
rlabel metal2 s 49392 59600 49448 60000 6 ay8913_do[2]
port 21 nsew signal input
rlabel metal2 s 49840 59600 49896 60000 6 ay8913_do[3]
port 22 nsew signal input
rlabel metal2 s 50288 59600 50344 60000 6 ay8913_do[4]
port 23 nsew signal input
rlabel metal2 s 50736 59600 50792 60000 6 ay8913_do[5]
port 24 nsew signal input
rlabel metal2 s 51184 59600 51240 60000 6 ay8913_do[6]
port 25 nsew signal input
rlabel metal2 s 51632 59600 51688 60000 6 ay8913_do[7]
port 26 nsew signal input
rlabel metal2 s 52080 59600 52136 60000 6 ay8913_do[8]
port 27 nsew signal input
rlabel metal2 s 52528 59600 52584 60000 6 ay8913_do[9]
port 28 nsew signal input
rlabel metal2 s 39984 59600 40040 60000 6 blinker_do[0]
port 29 nsew signal input
rlabel metal2 s 40432 59600 40488 60000 6 blinker_do[1]
port 30 nsew signal input
rlabel metal2 s 40880 59600 40936 60000 6 blinker_do[2]
port 31 nsew signal input
rlabel metal3 s 64600 19824 65000 19880 6 custom_settings[0]
port 32 nsew signal output
rlabel metal3 s 64600 24304 65000 24360 6 custom_settings[10]
port 33 nsew signal output
rlabel metal3 s 64600 24752 65000 24808 6 custom_settings[11]
port 34 nsew signal output
rlabel metal3 s 64600 25200 65000 25256 6 custom_settings[12]
port 35 nsew signal output
rlabel metal3 s 64600 25648 65000 25704 6 custom_settings[13]
port 36 nsew signal output
rlabel metal3 s 64600 26096 65000 26152 6 custom_settings[14]
port 37 nsew signal output
rlabel metal3 s 64600 26544 65000 26600 6 custom_settings[15]
port 38 nsew signal output
rlabel metal3 s 64600 26992 65000 27048 6 custom_settings[16]
port 39 nsew signal output
rlabel metal3 s 64600 27440 65000 27496 6 custom_settings[17]
port 40 nsew signal output
rlabel metal3 s 64600 27888 65000 27944 6 custom_settings[18]
port 41 nsew signal output
rlabel metal3 s 64600 28336 65000 28392 6 custom_settings[19]
port 42 nsew signal output
rlabel metal3 s 64600 20272 65000 20328 6 custom_settings[1]
port 43 nsew signal output
rlabel metal3 s 64600 28784 65000 28840 6 custom_settings[20]
port 44 nsew signal output
rlabel metal3 s 64600 29232 65000 29288 6 custom_settings[21]
port 45 nsew signal output
rlabel metal3 s 64600 29680 65000 29736 6 custom_settings[22]
port 46 nsew signal output
rlabel metal3 s 64600 30128 65000 30184 6 custom_settings[23]
port 47 nsew signal output
rlabel metal3 s 64600 30576 65000 30632 6 custom_settings[24]
port 48 nsew signal output
rlabel metal3 s 64600 31024 65000 31080 6 custom_settings[25]
port 49 nsew signal output
rlabel metal3 s 64600 31472 65000 31528 6 custom_settings[26]
port 50 nsew signal output
rlabel metal3 s 64600 31920 65000 31976 6 custom_settings[27]
port 51 nsew signal output
rlabel metal3 s 64600 32368 65000 32424 6 custom_settings[28]
port 52 nsew signal output
rlabel metal3 s 64600 32816 65000 32872 6 custom_settings[29]
port 53 nsew signal output
rlabel metal3 s 64600 20720 65000 20776 6 custom_settings[2]
port 54 nsew signal output
rlabel metal3 s 64600 33264 65000 33320 6 custom_settings[30]
port 55 nsew signal output
rlabel metal3 s 64600 33712 65000 33768 6 custom_settings[31]
port 56 nsew signal output
rlabel metal3 s 64600 21168 65000 21224 6 custom_settings[3]
port 57 nsew signal output
rlabel metal3 s 64600 21616 65000 21672 6 custom_settings[4]
port 58 nsew signal output
rlabel metal3 s 64600 22064 65000 22120 6 custom_settings[5]
port 59 nsew signal output
rlabel metal3 s 64600 22512 65000 22568 6 custom_settings[6]
port 60 nsew signal output
rlabel metal3 s 64600 22960 65000 23016 6 custom_settings[7]
port 61 nsew signal output
rlabel metal3 s 64600 23408 65000 23464 6 custom_settings[8]
port 62 nsew signal output
rlabel metal3 s 64600 23856 65000 23912 6 custom_settings[9]
port 63 nsew signal output
rlabel metal3 s 0 56560 400 56616 6 hellorld_do
port 64 nsew signal input
rlabel metal2 s 4144 59600 4200 60000 6 io_in[0]
port 65 nsew signal input
rlabel metal2 s 8624 59600 8680 60000 6 io_in[10]
port 66 nsew signal input
rlabel metal2 s 9072 59600 9128 60000 6 io_in[11]
port 67 nsew signal input
rlabel metal2 s 9520 59600 9576 60000 6 io_in[12]
port 68 nsew signal input
rlabel metal2 s 9968 59600 10024 60000 6 io_in[13]
port 69 nsew signal input
rlabel metal2 s 10416 59600 10472 60000 6 io_in[14]
port 70 nsew signal input
rlabel metal2 s 10864 59600 10920 60000 6 io_in[15]
port 71 nsew signal input
rlabel metal2 s 11312 59600 11368 60000 6 io_in[16]
port 72 nsew signal input
rlabel metal2 s 11760 59600 11816 60000 6 io_in[17]
port 73 nsew signal input
rlabel metal2 s 12208 59600 12264 60000 6 io_in[18]
port 74 nsew signal input
rlabel metal2 s 12656 59600 12712 60000 6 io_in[19]
port 75 nsew signal input
rlabel metal2 s 4592 59600 4648 60000 6 io_in[1]
port 76 nsew signal input
rlabel metal2 s 13104 59600 13160 60000 6 io_in[20]
port 77 nsew signal input
rlabel metal2 s 13552 59600 13608 60000 6 io_in[21]
port 78 nsew signal input
rlabel metal2 s 14000 59600 14056 60000 6 io_in[22]
port 79 nsew signal input
rlabel metal2 s 14448 59600 14504 60000 6 io_in[23]
port 80 nsew signal input
rlabel metal2 s 14896 59600 14952 60000 6 io_in[24]
port 81 nsew signal input
rlabel metal2 s 15344 59600 15400 60000 6 io_in[25]
port 82 nsew signal input
rlabel metal2 s 15792 59600 15848 60000 6 io_in[26]
port 83 nsew signal input
rlabel metal2 s 16240 59600 16296 60000 6 io_in[27]
port 84 nsew signal input
rlabel metal2 s 16688 59600 16744 60000 6 io_in[28]
port 85 nsew signal input
rlabel metal2 s 17136 59600 17192 60000 6 io_in[29]
port 86 nsew signal input
rlabel metal2 s 5040 59600 5096 60000 6 io_in[2]
port 87 nsew signal input
rlabel metal2 s 17584 59600 17640 60000 6 io_in[30]
port 88 nsew signal input
rlabel metal2 s 18032 59600 18088 60000 6 io_in[31]
port 89 nsew signal input
rlabel metal2 s 18480 59600 18536 60000 6 io_in[32]
port 90 nsew signal input
rlabel metal2 s 18928 59600 18984 60000 6 io_in[33]
port 91 nsew signal input
rlabel metal2 s 19376 59600 19432 60000 6 io_in[34]
port 92 nsew signal input
rlabel metal2 s 19824 59600 19880 60000 6 io_in[35]
port 93 nsew signal input
rlabel metal2 s 20272 59600 20328 60000 6 io_in[36]
port 94 nsew signal input
rlabel metal2 s 20720 59600 20776 60000 6 io_in[37]
port 95 nsew signal input
rlabel metal2 s 5488 59600 5544 60000 6 io_in[3]
port 96 nsew signal input
rlabel metal2 s 5936 59600 5992 60000 6 io_in[4]
port 97 nsew signal input
rlabel metal2 s 6384 59600 6440 60000 6 io_in[5]
port 98 nsew signal input
rlabel metal2 s 6832 59600 6888 60000 6 io_in[6]
port 99 nsew signal input
rlabel metal2 s 7280 59600 7336 60000 6 io_in[7]
port 100 nsew signal input
rlabel metal2 s 7728 59600 7784 60000 6 io_in[8]
port 101 nsew signal input
rlabel metal2 s 8176 59600 8232 60000 6 io_in[9]
port 102 nsew signal input
rlabel metal3 s 0 3360 400 3416 6 io_oeb[0]
port 103 nsew signal output
rlabel metal3 s 0 8960 400 9016 6 io_oeb[10]
port 104 nsew signal output
rlabel metal3 s 0 9520 400 9576 6 io_oeb[11]
port 105 nsew signal output
rlabel metal3 s 0 10080 400 10136 6 io_oeb[12]
port 106 nsew signal output
rlabel metal3 s 0 10640 400 10696 6 io_oeb[13]
port 107 nsew signal output
rlabel metal3 s 0 11200 400 11256 6 io_oeb[14]
port 108 nsew signal output
rlabel metal3 s 0 11760 400 11816 6 io_oeb[15]
port 109 nsew signal output
rlabel metal3 s 0 12320 400 12376 6 io_oeb[16]
port 110 nsew signal output
rlabel metal3 s 0 12880 400 12936 6 io_oeb[17]
port 111 nsew signal output
rlabel metal3 s 0 13440 400 13496 6 io_oeb[18]
port 112 nsew signal output
rlabel metal3 s 0 14000 400 14056 6 io_oeb[19]
port 113 nsew signal output
rlabel metal3 s 0 3920 400 3976 6 io_oeb[1]
port 114 nsew signal output
rlabel metal3 s 0 14560 400 14616 6 io_oeb[20]
port 115 nsew signal output
rlabel metal3 s 0 15120 400 15176 6 io_oeb[21]
port 116 nsew signal output
rlabel metal3 s 0 15680 400 15736 6 io_oeb[22]
port 117 nsew signal output
rlabel metal3 s 0 16240 400 16296 6 io_oeb[23]
port 118 nsew signal output
rlabel metal3 s 0 16800 400 16856 6 io_oeb[24]
port 119 nsew signal output
rlabel metal3 s 0 17360 400 17416 6 io_oeb[25]
port 120 nsew signal output
rlabel metal3 s 0 17920 400 17976 6 io_oeb[26]
port 121 nsew signal output
rlabel metal3 s 0 18480 400 18536 6 io_oeb[27]
port 122 nsew signal output
rlabel metal3 s 0 19040 400 19096 6 io_oeb[28]
port 123 nsew signal output
rlabel metal3 s 0 19600 400 19656 6 io_oeb[29]
port 124 nsew signal output
rlabel metal3 s 0 4480 400 4536 6 io_oeb[2]
port 125 nsew signal output
rlabel metal3 s 0 20160 400 20216 6 io_oeb[30]
port 126 nsew signal output
rlabel metal3 s 0 20720 400 20776 6 io_oeb[31]
port 127 nsew signal output
rlabel metal3 s 0 21280 400 21336 6 io_oeb[32]
port 128 nsew signal output
rlabel metal3 s 0 21840 400 21896 6 io_oeb[33]
port 129 nsew signal output
rlabel metal3 s 0 22400 400 22456 6 io_oeb[34]
port 130 nsew signal output
rlabel metal3 s 0 22960 400 23016 6 io_oeb[35]
port 131 nsew signal output
rlabel metal3 s 0 23520 400 23576 6 io_oeb[36]
port 132 nsew signal output
rlabel metal3 s 0 24080 400 24136 6 io_oeb[37]
port 133 nsew signal output
rlabel metal3 s 0 5040 400 5096 6 io_oeb[3]
port 134 nsew signal output
rlabel metal3 s 0 5600 400 5656 6 io_oeb[4]
port 135 nsew signal output
rlabel metal3 s 0 6160 400 6216 6 io_oeb[5]
port 136 nsew signal output
rlabel metal3 s 0 6720 400 6776 6 io_oeb[6]
port 137 nsew signal output
rlabel metal3 s 0 7280 400 7336 6 io_oeb[7]
port 138 nsew signal output
rlabel metal3 s 0 7840 400 7896 6 io_oeb[8]
port 139 nsew signal output
rlabel metal3 s 0 8400 400 8456 6 io_oeb[9]
port 140 nsew signal output
rlabel metal2 s 21168 59600 21224 60000 6 io_out[0]
port 141 nsew signal output
rlabel metal2 s 25648 59600 25704 60000 6 io_out[10]
port 142 nsew signal output
rlabel metal2 s 26096 59600 26152 60000 6 io_out[11]
port 143 nsew signal output
rlabel metal2 s 26544 59600 26600 60000 6 io_out[12]
port 144 nsew signal output
rlabel metal2 s 26992 59600 27048 60000 6 io_out[13]
port 145 nsew signal output
rlabel metal2 s 27440 59600 27496 60000 6 io_out[14]
port 146 nsew signal output
rlabel metal2 s 27888 59600 27944 60000 6 io_out[15]
port 147 nsew signal output
rlabel metal2 s 28336 59600 28392 60000 6 io_out[16]
port 148 nsew signal output
rlabel metal2 s 28784 59600 28840 60000 6 io_out[17]
port 149 nsew signal output
rlabel metal2 s 29232 59600 29288 60000 6 io_out[18]
port 150 nsew signal output
rlabel metal2 s 29680 59600 29736 60000 6 io_out[19]
port 151 nsew signal output
rlabel metal2 s 21616 59600 21672 60000 6 io_out[1]
port 152 nsew signal output
rlabel metal2 s 30128 59600 30184 60000 6 io_out[20]
port 153 nsew signal output
rlabel metal2 s 30576 59600 30632 60000 6 io_out[21]
port 154 nsew signal output
rlabel metal2 s 31024 59600 31080 60000 6 io_out[22]
port 155 nsew signal output
rlabel metal2 s 31472 59600 31528 60000 6 io_out[23]
port 156 nsew signal output
rlabel metal2 s 31920 59600 31976 60000 6 io_out[24]
port 157 nsew signal output
rlabel metal2 s 32368 59600 32424 60000 6 io_out[25]
port 158 nsew signal output
rlabel metal2 s 32816 59600 32872 60000 6 io_out[26]
port 159 nsew signal output
rlabel metal2 s 33264 59600 33320 60000 6 io_out[27]
port 160 nsew signal output
rlabel metal2 s 33712 59600 33768 60000 6 io_out[28]
port 161 nsew signal output
rlabel metal2 s 34160 59600 34216 60000 6 io_out[29]
port 162 nsew signal output
rlabel metal2 s 22064 59600 22120 60000 6 io_out[2]
port 163 nsew signal output
rlabel metal2 s 34608 59600 34664 60000 6 io_out[30]
port 164 nsew signal output
rlabel metal2 s 35056 59600 35112 60000 6 io_out[31]
port 165 nsew signal output
rlabel metal2 s 35504 59600 35560 60000 6 io_out[32]
port 166 nsew signal output
rlabel metal2 s 35952 59600 36008 60000 6 io_out[33]
port 167 nsew signal output
rlabel metal2 s 36400 59600 36456 60000 6 io_out[34]
port 168 nsew signal output
rlabel metal2 s 36848 59600 36904 60000 6 io_out[35]
port 169 nsew signal output
rlabel metal2 s 37296 59600 37352 60000 6 io_out[36]
port 170 nsew signal output
rlabel metal2 s 37744 59600 37800 60000 6 io_out[37]
port 171 nsew signal output
rlabel metal2 s 22512 59600 22568 60000 6 io_out[3]
port 172 nsew signal output
rlabel metal2 s 22960 59600 23016 60000 6 io_out[4]
port 173 nsew signal output
rlabel metal2 s 23408 59600 23464 60000 6 io_out[5]
port 174 nsew signal output
rlabel metal2 s 23856 59600 23912 60000 6 io_out[6]
port 175 nsew signal output
rlabel metal2 s 24304 59600 24360 60000 6 io_out[7]
port 176 nsew signal output
rlabel metal2 s 24752 59600 24808 60000 6 io_out[8]
port 177 nsew signal output
rlabel metal2 s 25200 59600 25256 60000 6 io_out[9]
port 178 nsew signal output
rlabel metal2 s 38192 59600 38248 60000 6 irq[0]
port 179 nsew signal output
rlabel metal2 s 38640 59600 38696 60000 6 irq[1]
port 180 nsew signal output
rlabel metal2 s 39088 59600 39144 60000 6 irq[2]
port 181 nsew signal output
rlabel metal3 s 0 38640 400 38696 6 mc14500_do[0]
port 182 nsew signal input
rlabel metal3 s 0 44240 400 44296 6 mc14500_do[10]
port 183 nsew signal input
rlabel metal3 s 0 44800 400 44856 6 mc14500_do[11]
port 184 nsew signal input
rlabel metal3 s 0 45360 400 45416 6 mc14500_do[12]
port 185 nsew signal input
rlabel metal3 s 0 45920 400 45976 6 mc14500_do[13]
port 186 nsew signal input
rlabel metal3 s 0 46480 400 46536 6 mc14500_do[14]
port 187 nsew signal input
rlabel metal3 s 0 47040 400 47096 6 mc14500_do[15]
port 188 nsew signal input
rlabel metal3 s 0 47600 400 47656 6 mc14500_do[16]
port 189 nsew signal input
rlabel metal3 s 0 48160 400 48216 6 mc14500_do[17]
port 190 nsew signal input
rlabel metal3 s 0 48720 400 48776 6 mc14500_do[18]
port 191 nsew signal input
rlabel metal3 s 0 49280 400 49336 6 mc14500_do[19]
port 192 nsew signal input
rlabel metal3 s 0 39200 400 39256 6 mc14500_do[1]
port 193 nsew signal input
rlabel metal3 s 0 49840 400 49896 6 mc14500_do[20]
port 194 nsew signal input
rlabel metal3 s 0 50400 400 50456 6 mc14500_do[21]
port 195 nsew signal input
rlabel metal3 s 0 50960 400 51016 6 mc14500_do[22]
port 196 nsew signal input
rlabel metal3 s 0 51520 400 51576 6 mc14500_do[23]
port 197 nsew signal input
rlabel metal3 s 0 52080 400 52136 6 mc14500_do[24]
port 198 nsew signal input
rlabel metal3 s 0 52640 400 52696 6 mc14500_do[25]
port 199 nsew signal input
rlabel metal3 s 0 53200 400 53256 6 mc14500_do[26]
port 200 nsew signal input
rlabel metal3 s 0 53760 400 53816 6 mc14500_do[27]
port 201 nsew signal input
rlabel metal3 s 0 54320 400 54376 6 mc14500_do[28]
port 202 nsew signal input
rlabel metal3 s 0 54880 400 54936 6 mc14500_do[29]
port 203 nsew signal input
rlabel metal3 s 0 39760 400 39816 6 mc14500_do[2]
port 204 nsew signal input
rlabel metal3 s 0 55440 400 55496 6 mc14500_do[30]
port 205 nsew signal input
rlabel metal3 s 0 40320 400 40376 6 mc14500_do[3]
port 206 nsew signal input
rlabel metal3 s 0 40880 400 40936 6 mc14500_do[4]
port 207 nsew signal input
rlabel metal3 s 0 41440 400 41496 6 mc14500_do[5]
port 208 nsew signal input
rlabel metal3 s 0 42000 400 42056 6 mc14500_do[6]
port 209 nsew signal input
rlabel metal3 s 0 42560 400 42616 6 mc14500_do[7]
port 210 nsew signal input
rlabel metal3 s 0 43120 400 43176 6 mc14500_do[8]
port 211 nsew signal input
rlabel metal3 s 0 43680 400 43736 6 mc14500_do[9]
port 212 nsew signal input
rlabel metal2 s 41776 59600 41832 60000 6 mc14500_sram_addr[0]
port 213 nsew signal input
rlabel metal2 s 42224 59600 42280 60000 6 mc14500_sram_addr[1]
port 214 nsew signal input
rlabel metal2 s 42672 59600 42728 60000 6 mc14500_sram_addr[2]
port 215 nsew signal input
rlabel metal2 s 43120 59600 43176 60000 6 mc14500_sram_addr[3]
port 216 nsew signal input
rlabel metal2 s 43568 59600 43624 60000 6 mc14500_sram_addr[4]
port 217 nsew signal input
rlabel metal2 s 44016 59600 44072 60000 6 mc14500_sram_addr[5]
port 218 nsew signal input
rlabel metal2 s 48048 59600 48104 60000 6 mc14500_sram_gwe
port 219 nsew signal input
rlabel metal2 s 44464 59600 44520 60000 6 mc14500_sram_in[0]
port 220 nsew signal input
rlabel metal2 s 44912 59600 44968 60000 6 mc14500_sram_in[1]
port 221 nsew signal input
rlabel metal2 s 45360 59600 45416 60000 6 mc14500_sram_in[2]
port 222 nsew signal input
rlabel metal2 s 45808 59600 45864 60000 6 mc14500_sram_in[3]
port 223 nsew signal input
rlabel metal2 s 46256 59600 46312 60000 6 mc14500_sram_in[4]
port 224 nsew signal input
rlabel metal2 s 46704 59600 46760 60000 6 mc14500_sram_in[5]
port 225 nsew signal input
rlabel metal2 s 47152 59600 47208 60000 6 mc14500_sram_in[6]
port 226 nsew signal input
rlabel metal2 s 47600 59600 47656 60000 6 mc14500_sram_in[7]
port 227 nsew signal input
rlabel metal2 s 44688 0 44744 400 6 qcpu_do[0]
port 228 nsew signal input
rlabel metal2 s 49168 0 49224 400 6 qcpu_do[10]
port 229 nsew signal input
rlabel metal2 s 49616 0 49672 400 6 qcpu_do[11]
port 230 nsew signal input
rlabel metal2 s 50064 0 50120 400 6 qcpu_do[12]
port 231 nsew signal input
rlabel metal2 s 50512 0 50568 400 6 qcpu_do[13]
port 232 nsew signal input
rlabel metal2 s 50960 0 51016 400 6 qcpu_do[14]
port 233 nsew signal input
rlabel metal2 s 51408 0 51464 400 6 qcpu_do[15]
port 234 nsew signal input
rlabel metal2 s 51856 0 51912 400 6 qcpu_do[16]
port 235 nsew signal input
rlabel metal2 s 52304 0 52360 400 6 qcpu_do[17]
port 236 nsew signal input
rlabel metal2 s 52752 0 52808 400 6 qcpu_do[18]
port 237 nsew signal input
rlabel metal2 s 53200 0 53256 400 6 qcpu_do[19]
port 238 nsew signal input
rlabel metal2 s 45136 0 45192 400 6 qcpu_do[1]
port 239 nsew signal input
rlabel metal2 s 53648 0 53704 400 6 qcpu_do[20]
port 240 nsew signal input
rlabel metal2 s 54096 0 54152 400 6 qcpu_do[21]
port 241 nsew signal input
rlabel metal2 s 54544 0 54600 400 6 qcpu_do[22]
port 242 nsew signal input
rlabel metal2 s 54992 0 55048 400 6 qcpu_do[23]
port 243 nsew signal input
rlabel metal2 s 55440 0 55496 400 6 qcpu_do[24]
port 244 nsew signal input
rlabel metal2 s 55888 0 55944 400 6 qcpu_do[25]
port 245 nsew signal input
rlabel metal2 s 56336 0 56392 400 6 qcpu_do[26]
port 246 nsew signal input
rlabel metal2 s 56784 0 56840 400 6 qcpu_do[27]
port 247 nsew signal input
rlabel metal2 s 57232 0 57288 400 6 qcpu_do[28]
port 248 nsew signal input
rlabel metal2 s 57680 0 57736 400 6 qcpu_do[29]
port 249 nsew signal input
rlabel metal2 s 45584 0 45640 400 6 qcpu_do[2]
port 250 nsew signal input
rlabel metal2 s 58128 0 58184 400 6 qcpu_do[30]
port 251 nsew signal input
rlabel metal2 s 58576 0 58632 400 6 qcpu_do[31]
port 252 nsew signal input
rlabel metal2 s 59024 0 59080 400 6 qcpu_do[32]
port 253 nsew signal input
rlabel metal2 s 46032 0 46088 400 6 qcpu_do[3]
port 254 nsew signal input
rlabel metal2 s 46480 0 46536 400 6 qcpu_do[4]
port 255 nsew signal input
rlabel metal2 s 46928 0 46984 400 6 qcpu_do[5]
port 256 nsew signal input
rlabel metal2 s 47376 0 47432 400 6 qcpu_do[6]
port 257 nsew signal input
rlabel metal2 s 47824 0 47880 400 6 qcpu_do[7]
port 258 nsew signal input
rlabel metal2 s 48272 0 48328 400 6 qcpu_do[8]
port 259 nsew signal input
rlabel metal2 s 48720 0 48776 400 6 qcpu_do[9]
port 260 nsew signal input
rlabel metal3 s 64600 34160 65000 34216 6 qcpu_oeb[0]
port 261 nsew signal input
rlabel metal3 s 64600 38640 65000 38696 6 qcpu_oeb[10]
port 262 nsew signal input
rlabel metal3 s 64600 39088 65000 39144 6 qcpu_oeb[11]
port 263 nsew signal input
rlabel metal3 s 64600 39536 65000 39592 6 qcpu_oeb[12]
port 264 nsew signal input
rlabel metal3 s 64600 39984 65000 40040 6 qcpu_oeb[13]
port 265 nsew signal input
rlabel metal3 s 64600 40432 65000 40488 6 qcpu_oeb[14]
port 266 nsew signal input
rlabel metal3 s 64600 40880 65000 40936 6 qcpu_oeb[15]
port 267 nsew signal input
rlabel metal3 s 64600 41328 65000 41384 6 qcpu_oeb[16]
port 268 nsew signal input
rlabel metal3 s 64600 41776 65000 41832 6 qcpu_oeb[17]
port 269 nsew signal input
rlabel metal3 s 64600 42224 65000 42280 6 qcpu_oeb[18]
port 270 nsew signal input
rlabel metal3 s 64600 42672 65000 42728 6 qcpu_oeb[19]
port 271 nsew signal input
rlabel metal3 s 64600 34608 65000 34664 6 qcpu_oeb[1]
port 272 nsew signal input
rlabel metal3 s 64600 43120 65000 43176 6 qcpu_oeb[20]
port 273 nsew signal input
rlabel metal3 s 64600 43568 65000 43624 6 qcpu_oeb[21]
port 274 nsew signal input
rlabel metal3 s 64600 44016 65000 44072 6 qcpu_oeb[22]
port 275 nsew signal input
rlabel metal3 s 64600 44464 65000 44520 6 qcpu_oeb[23]
port 276 nsew signal input
rlabel metal3 s 64600 44912 65000 44968 6 qcpu_oeb[24]
port 277 nsew signal input
rlabel metal3 s 64600 45360 65000 45416 6 qcpu_oeb[25]
port 278 nsew signal input
rlabel metal3 s 64600 45808 65000 45864 6 qcpu_oeb[26]
port 279 nsew signal input
rlabel metal3 s 64600 46256 65000 46312 6 qcpu_oeb[27]
port 280 nsew signal input
rlabel metal3 s 64600 46704 65000 46760 6 qcpu_oeb[28]
port 281 nsew signal input
rlabel metal3 s 64600 47152 65000 47208 6 qcpu_oeb[29]
port 282 nsew signal input
rlabel metal3 s 64600 35056 65000 35112 6 qcpu_oeb[2]
port 283 nsew signal input
rlabel metal3 s 64600 47600 65000 47656 6 qcpu_oeb[30]
port 284 nsew signal input
rlabel metal3 s 64600 48048 65000 48104 6 qcpu_oeb[31]
port 285 nsew signal input
rlabel metal3 s 64600 48496 65000 48552 6 qcpu_oeb[32]
port 286 nsew signal input
rlabel metal3 s 64600 35504 65000 35560 6 qcpu_oeb[3]
port 287 nsew signal input
rlabel metal3 s 64600 35952 65000 36008 6 qcpu_oeb[4]
port 288 nsew signal input
rlabel metal3 s 64600 36400 65000 36456 6 qcpu_oeb[5]
port 289 nsew signal input
rlabel metal3 s 64600 36848 65000 36904 6 qcpu_oeb[6]
port 290 nsew signal input
rlabel metal3 s 64600 37296 65000 37352 6 qcpu_oeb[7]
port 291 nsew signal input
rlabel metal3 s 64600 37744 65000 37800 6 qcpu_oeb[8]
port 292 nsew signal input
rlabel metal3 s 64600 38192 65000 38248 6 qcpu_oeb[9]
port 293 nsew signal input
rlabel metal2 s 59472 0 59528 400 6 qcpu_sram_addr[0]
port 294 nsew signal input
rlabel metal2 s 59920 0 59976 400 6 qcpu_sram_addr[1]
port 295 nsew signal input
rlabel metal2 s 60368 0 60424 400 6 qcpu_sram_addr[2]
port 296 nsew signal input
rlabel metal2 s 60816 0 60872 400 6 qcpu_sram_addr[3]
port 297 nsew signal input
rlabel metal2 s 61264 0 61320 400 6 qcpu_sram_addr[4]
port 298 nsew signal input
rlabel metal2 s 61712 0 61768 400 6 qcpu_sram_addr[5]
port 299 nsew signal input
rlabel metal2 s 62160 0 62216 400 6 qcpu_sram_gwe
port 300 nsew signal input
rlabel metal3 s 64600 48944 65000 49000 6 qcpu_sram_in[0]
port 301 nsew signal input
rlabel metal3 s 64600 49392 65000 49448 6 qcpu_sram_in[1]
port 302 nsew signal input
rlabel metal3 s 64600 49840 65000 49896 6 qcpu_sram_in[2]
port 303 nsew signal input
rlabel metal3 s 64600 50288 65000 50344 6 qcpu_sram_in[3]
port 304 nsew signal input
rlabel metal3 s 64600 50736 65000 50792 6 qcpu_sram_in[4]
port 305 nsew signal input
rlabel metal3 s 64600 51184 65000 51240 6 qcpu_sram_in[5]
port 306 nsew signal input
rlabel metal3 s 64600 51632 65000 51688 6 qcpu_sram_in[6]
port 307 nsew signal input
rlabel metal3 s 64600 52080 65000 52136 6 qcpu_sram_in[7]
port 308 nsew signal input
rlabel metal3 s 64600 52528 65000 52584 6 qcpu_sram_out[0]
port 309 nsew signal output
rlabel metal3 s 64600 52976 65000 53032 6 qcpu_sram_out[1]
port 310 nsew signal output
rlabel metal3 s 64600 53424 65000 53480 6 qcpu_sram_out[2]
port 311 nsew signal output
rlabel metal3 s 64600 53872 65000 53928 6 qcpu_sram_out[3]
port 312 nsew signal output
rlabel metal3 s 64600 54320 65000 54376 6 qcpu_sram_out[4]
port 313 nsew signal output
rlabel metal3 s 64600 54768 65000 54824 6 qcpu_sram_out[5]
port 314 nsew signal output
rlabel metal3 s 64600 55216 65000 55272 6 qcpu_sram_out[6]
port 315 nsew signal output
rlabel metal3 s 64600 55664 65000 55720 6 qcpu_sram_out[7]
port 316 nsew signal output
rlabel metal3 s 64600 56112 65000 56168 6 rst_ay8913
port 317 nsew signal output
rlabel metal2 s 39536 59600 39592 60000 6 rst_blinker
port 318 nsew signal output
rlabel metal3 s 0 56000 400 56056 6 rst_hellorld
port 319 nsew signal output
rlabel metal3 s 0 38080 400 38136 6 rst_mc14500
port 320 nsew signal output
rlabel metal3 s 0 37520 400 37576 6 rst_qcpu
port 321 nsew signal output
rlabel metal3 s 0 24640 400 24696 6 rst_sid
port 322 nsew signal output
rlabel metal2 s 41328 59600 41384 60000 6 rst_sn76489
port 323 nsew signal output
rlabel metal3 s 0 25200 400 25256 6 sid_do[0]
port 324 nsew signal input
rlabel metal3 s 0 30800 400 30856 6 sid_do[10]
port 325 nsew signal input
rlabel metal3 s 0 31360 400 31416 6 sid_do[11]
port 326 nsew signal input
rlabel metal3 s 0 31920 400 31976 6 sid_do[12]
port 327 nsew signal input
rlabel metal3 s 0 32480 400 32536 6 sid_do[13]
port 328 nsew signal input
rlabel metal3 s 0 33040 400 33096 6 sid_do[14]
port 329 nsew signal input
rlabel metal3 s 0 33600 400 33656 6 sid_do[15]
port 330 nsew signal input
rlabel metal3 s 0 34160 400 34216 6 sid_do[16]
port 331 nsew signal input
rlabel metal3 s 0 34720 400 34776 6 sid_do[17]
port 332 nsew signal input
rlabel metal3 s 0 35280 400 35336 6 sid_do[18]
port 333 nsew signal input
rlabel metal3 s 0 35840 400 35896 6 sid_do[19]
port 334 nsew signal input
rlabel metal3 s 0 25760 400 25816 6 sid_do[1]
port 335 nsew signal input
rlabel metal3 s 0 36400 400 36456 6 sid_do[20]
port 336 nsew signal input
rlabel metal3 s 0 26320 400 26376 6 sid_do[2]
port 337 nsew signal input
rlabel metal3 s 0 26880 400 26936 6 sid_do[3]
port 338 nsew signal input
rlabel metal3 s 0 27440 400 27496 6 sid_do[4]
port 339 nsew signal input
rlabel metal3 s 0 28000 400 28056 6 sid_do[5]
port 340 nsew signal input
rlabel metal3 s 0 28560 400 28616 6 sid_do[6]
port 341 nsew signal input
rlabel metal3 s 0 29120 400 29176 6 sid_do[7]
port 342 nsew signal input
rlabel metal3 s 0 29680 400 29736 6 sid_do[8]
port 343 nsew signal input
rlabel metal3 s 0 30240 400 30296 6 sid_do[9]
port 344 nsew signal input
rlabel metal3 s 0 36960 400 37016 6 sid_oeb
port 345 nsew signal input
rlabel metal2 s 32144 0 32200 400 6 sn76489_do[0]
port 346 nsew signal input
rlabel metal2 s 36624 0 36680 400 6 sn76489_do[10]
port 347 nsew signal input
rlabel metal2 s 37072 0 37128 400 6 sn76489_do[11]
port 348 nsew signal input
rlabel metal2 s 37520 0 37576 400 6 sn76489_do[12]
port 349 nsew signal input
rlabel metal2 s 37968 0 38024 400 6 sn76489_do[13]
port 350 nsew signal input
rlabel metal2 s 38416 0 38472 400 6 sn76489_do[14]
port 351 nsew signal input
rlabel metal2 s 38864 0 38920 400 6 sn76489_do[15]
port 352 nsew signal input
rlabel metal2 s 39312 0 39368 400 6 sn76489_do[16]
port 353 nsew signal input
rlabel metal2 s 39760 0 39816 400 6 sn76489_do[17]
port 354 nsew signal input
rlabel metal2 s 40208 0 40264 400 6 sn76489_do[18]
port 355 nsew signal input
rlabel metal2 s 40656 0 40712 400 6 sn76489_do[19]
port 356 nsew signal input
rlabel metal2 s 32592 0 32648 400 6 sn76489_do[1]
port 357 nsew signal input
rlabel metal2 s 41104 0 41160 400 6 sn76489_do[20]
port 358 nsew signal input
rlabel metal2 s 41552 0 41608 400 6 sn76489_do[21]
port 359 nsew signal input
rlabel metal2 s 42000 0 42056 400 6 sn76489_do[22]
port 360 nsew signal input
rlabel metal2 s 42448 0 42504 400 6 sn76489_do[23]
port 361 nsew signal input
rlabel metal2 s 42896 0 42952 400 6 sn76489_do[24]
port 362 nsew signal input
rlabel metal2 s 43344 0 43400 400 6 sn76489_do[25]
port 363 nsew signal input
rlabel metal2 s 43792 0 43848 400 6 sn76489_do[26]
port 364 nsew signal input
rlabel metal2 s 44240 0 44296 400 6 sn76489_do[27]
port 365 nsew signal input
rlabel metal2 s 33040 0 33096 400 6 sn76489_do[2]
port 366 nsew signal input
rlabel metal2 s 33488 0 33544 400 6 sn76489_do[3]
port 367 nsew signal input
rlabel metal2 s 33936 0 33992 400 6 sn76489_do[4]
port 368 nsew signal input
rlabel metal2 s 34384 0 34440 400 6 sn76489_do[5]
port 369 nsew signal input
rlabel metal2 s 34832 0 34888 400 6 sn76489_do[6]
port 370 nsew signal input
rlabel metal2 s 35280 0 35336 400 6 sn76489_do[7]
port 371 nsew signal input
rlabel metal2 s 35728 0 35784 400 6 sn76489_do[8]
port 372 nsew signal input
rlabel metal2 s 36176 0 36232 400 6 sn76489_do[9]
port 373 nsew signal input
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 374 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58438 6 vdd
port 374 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58438 6 vdd
port 374 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58438 6 vdd
port 374 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 58438 6 vdd
port 374 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58438 6 vss
port 375 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58438 6 vss
port 375 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58438 6 vss
port 375 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 58438 6 vss
port 375 nsew ground bidirectional
rlabel metal2 s 2576 0 2632 400 6 wb_clk_i
port 376 nsew signal input
rlabel metal2 s 3024 0 3080 400 6 wb_rst_i
port 377 nsew signal input
rlabel metal3 s 64600 19376 65000 19432 6 wbs_ack_o
port 378 nsew signal output
rlabel metal2 s 3472 0 3528 400 6 wbs_adr_i[0]
port 379 nsew signal input
rlabel metal2 s 7952 0 8008 400 6 wbs_adr_i[10]
port 380 nsew signal input
rlabel metal2 s 8400 0 8456 400 6 wbs_adr_i[11]
port 381 nsew signal input
rlabel metal2 s 8848 0 8904 400 6 wbs_adr_i[12]
port 382 nsew signal input
rlabel metal2 s 9296 0 9352 400 6 wbs_adr_i[13]
port 383 nsew signal input
rlabel metal2 s 9744 0 9800 400 6 wbs_adr_i[14]
port 384 nsew signal input
rlabel metal2 s 10192 0 10248 400 6 wbs_adr_i[15]
port 385 nsew signal input
rlabel metal2 s 10640 0 10696 400 6 wbs_adr_i[16]
port 386 nsew signal input
rlabel metal2 s 11088 0 11144 400 6 wbs_adr_i[17]
port 387 nsew signal input
rlabel metal2 s 11536 0 11592 400 6 wbs_adr_i[18]
port 388 nsew signal input
rlabel metal2 s 11984 0 12040 400 6 wbs_adr_i[19]
port 389 nsew signal input
rlabel metal2 s 3920 0 3976 400 6 wbs_adr_i[1]
port 390 nsew signal input
rlabel metal2 s 12432 0 12488 400 6 wbs_adr_i[20]
port 391 nsew signal input
rlabel metal2 s 12880 0 12936 400 6 wbs_adr_i[21]
port 392 nsew signal input
rlabel metal2 s 13328 0 13384 400 6 wbs_adr_i[22]
port 393 nsew signal input
rlabel metal2 s 13776 0 13832 400 6 wbs_adr_i[23]
port 394 nsew signal input
rlabel metal2 s 14224 0 14280 400 6 wbs_adr_i[24]
port 395 nsew signal input
rlabel metal2 s 14672 0 14728 400 6 wbs_adr_i[25]
port 396 nsew signal input
rlabel metal2 s 15120 0 15176 400 6 wbs_adr_i[26]
port 397 nsew signal input
rlabel metal2 s 15568 0 15624 400 6 wbs_adr_i[27]
port 398 nsew signal input
rlabel metal2 s 16016 0 16072 400 6 wbs_adr_i[28]
port 399 nsew signal input
rlabel metal2 s 16464 0 16520 400 6 wbs_adr_i[29]
port 400 nsew signal input
rlabel metal2 s 4368 0 4424 400 6 wbs_adr_i[2]
port 401 nsew signal input
rlabel metal2 s 16912 0 16968 400 6 wbs_adr_i[30]
port 402 nsew signal input
rlabel metal2 s 17360 0 17416 400 6 wbs_adr_i[31]
port 403 nsew signal input
rlabel metal2 s 4816 0 4872 400 6 wbs_adr_i[3]
port 404 nsew signal input
rlabel metal2 s 5264 0 5320 400 6 wbs_adr_i[4]
port 405 nsew signal input
rlabel metal2 s 5712 0 5768 400 6 wbs_adr_i[5]
port 406 nsew signal input
rlabel metal2 s 6160 0 6216 400 6 wbs_adr_i[6]
port 407 nsew signal input
rlabel metal2 s 6608 0 6664 400 6 wbs_adr_i[7]
port 408 nsew signal input
rlabel metal2 s 7056 0 7112 400 6 wbs_adr_i[8]
port 409 nsew signal input
rlabel metal2 s 7504 0 7560 400 6 wbs_adr_i[9]
port 410 nsew signal input
rlabel metal3 s 64600 18480 65000 18536 6 wbs_cyc_i
port 411 nsew signal input
rlabel metal2 s 17808 0 17864 400 6 wbs_dat_i[0]
port 412 nsew signal input
rlabel metal2 s 22288 0 22344 400 6 wbs_dat_i[10]
port 413 nsew signal input
rlabel metal2 s 22736 0 22792 400 6 wbs_dat_i[11]
port 414 nsew signal input
rlabel metal2 s 23184 0 23240 400 6 wbs_dat_i[12]
port 415 nsew signal input
rlabel metal2 s 23632 0 23688 400 6 wbs_dat_i[13]
port 416 nsew signal input
rlabel metal2 s 24080 0 24136 400 6 wbs_dat_i[14]
port 417 nsew signal input
rlabel metal2 s 24528 0 24584 400 6 wbs_dat_i[15]
port 418 nsew signal input
rlabel metal2 s 24976 0 25032 400 6 wbs_dat_i[16]
port 419 nsew signal input
rlabel metal2 s 25424 0 25480 400 6 wbs_dat_i[17]
port 420 nsew signal input
rlabel metal2 s 25872 0 25928 400 6 wbs_dat_i[18]
port 421 nsew signal input
rlabel metal2 s 26320 0 26376 400 6 wbs_dat_i[19]
port 422 nsew signal input
rlabel metal2 s 18256 0 18312 400 6 wbs_dat_i[1]
port 423 nsew signal input
rlabel metal2 s 26768 0 26824 400 6 wbs_dat_i[20]
port 424 nsew signal input
rlabel metal2 s 27216 0 27272 400 6 wbs_dat_i[21]
port 425 nsew signal input
rlabel metal2 s 27664 0 27720 400 6 wbs_dat_i[22]
port 426 nsew signal input
rlabel metal2 s 28112 0 28168 400 6 wbs_dat_i[23]
port 427 nsew signal input
rlabel metal2 s 28560 0 28616 400 6 wbs_dat_i[24]
port 428 nsew signal input
rlabel metal2 s 29008 0 29064 400 6 wbs_dat_i[25]
port 429 nsew signal input
rlabel metal2 s 29456 0 29512 400 6 wbs_dat_i[26]
port 430 nsew signal input
rlabel metal2 s 29904 0 29960 400 6 wbs_dat_i[27]
port 431 nsew signal input
rlabel metal2 s 30352 0 30408 400 6 wbs_dat_i[28]
port 432 nsew signal input
rlabel metal2 s 30800 0 30856 400 6 wbs_dat_i[29]
port 433 nsew signal input
rlabel metal2 s 18704 0 18760 400 6 wbs_dat_i[2]
port 434 nsew signal input
rlabel metal2 s 31248 0 31304 400 6 wbs_dat_i[30]
port 435 nsew signal input
rlabel metal2 s 31696 0 31752 400 6 wbs_dat_i[31]
port 436 nsew signal input
rlabel metal2 s 19152 0 19208 400 6 wbs_dat_i[3]
port 437 nsew signal input
rlabel metal2 s 19600 0 19656 400 6 wbs_dat_i[4]
port 438 nsew signal input
rlabel metal2 s 20048 0 20104 400 6 wbs_dat_i[5]
port 439 nsew signal input
rlabel metal2 s 20496 0 20552 400 6 wbs_dat_i[6]
port 440 nsew signal input
rlabel metal2 s 20944 0 21000 400 6 wbs_dat_i[7]
port 441 nsew signal input
rlabel metal2 s 21392 0 21448 400 6 wbs_dat_i[8]
port 442 nsew signal input
rlabel metal2 s 21840 0 21896 400 6 wbs_dat_i[9]
port 443 nsew signal input
rlabel metal3 s 64600 3696 65000 3752 6 wbs_dat_o[0]
port 444 nsew signal output
rlabel metal3 s 64600 8176 65000 8232 6 wbs_dat_o[10]
port 445 nsew signal output
rlabel metal3 s 64600 8624 65000 8680 6 wbs_dat_o[11]
port 446 nsew signal output
rlabel metal3 s 64600 9072 65000 9128 6 wbs_dat_o[12]
port 447 nsew signal output
rlabel metal3 s 64600 9520 65000 9576 6 wbs_dat_o[13]
port 448 nsew signal output
rlabel metal3 s 64600 9968 65000 10024 6 wbs_dat_o[14]
port 449 nsew signal output
rlabel metal3 s 64600 10416 65000 10472 6 wbs_dat_o[15]
port 450 nsew signal output
rlabel metal3 s 64600 10864 65000 10920 6 wbs_dat_o[16]
port 451 nsew signal output
rlabel metal3 s 64600 11312 65000 11368 6 wbs_dat_o[17]
port 452 nsew signal output
rlabel metal3 s 64600 11760 65000 11816 6 wbs_dat_o[18]
port 453 nsew signal output
rlabel metal3 s 64600 12208 65000 12264 6 wbs_dat_o[19]
port 454 nsew signal output
rlabel metal3 s 64600 4144 65000 4200 6 wbs_dat_o[1]
port 455 nsew signal output
rlabel metal3 s 64600 12656 65000 12712 6 wbs_dat_o[20]
port 456 nsew signal output
rlabel metal3 s 64600 13104 65000 13160 6 wbs_dat_o[21]
port 457 nsew signal output
rlabel metal3 s 64600 13552 65000 13608 6 wbs_dat_o[22]
port 458 nsew signal output
rlabel metal3 s 64600 14000 65000 14056 6 wbs_dat_o[23]
port 459 nsew signal output
rlabel metal3 s 64600 14448 65000 14504 6 wbs_dat_o[24]
port 460 nsew signal output
rlabel metal3 s 64600 14896 65000 14952 6 wbs_dat_o[25]
port 461 nsew signal output
rlabel metal3 s 64600 15344 65000 15400 6 wbs_dat_o[26]
port 462 nsew signal output
rlabel metal3 s 64600 15792 65000 15848 6 wbs_dat_o[27]
port 463 nsew signal output
rlabel metal3 s 64600 16240 65000 16296 6 wbs_dat_o[28]
port 464 nsew signal output
rlabel metal3 s 64600 16688 65000 16744 6 wbs_dat_o[29]
port 465 nsew signal output
rlabel metal3 s 64600 4592 65000 4648 6 wbs_dat_o[2]
port 466 nsew signal output
rlabel metal3 s 64600 17136 65000 17192 6 wbs_dat_o[30]
port 467 nsew signal output
rlabel metal3 s 64600 17584 65000 17640 6 wbs_dat_o[31]
port 468 nsew signal output
rlabel metal3 s 64600 5040 65000 5096 6 wbs_dat_o[3]
port 469 nsew signal output
rlabel metal3 s 64600 5488 65000 5544 6 wbs_dat_o[4]
port 470 nsew signal output
rlabel metal3 s 64600 5936 65000 5992 6 wbs_dat_o[5]
port 471 nsew signal output
rlabel metal3 s 64600 6384 65000 6440 6 wbs_dat_o[6]
port 472 nsew signal output
rlabel metal3 s 64600 6832 65000 6888 6 wbs_dat_o[7]
port 473 nsew signal output
rlabel metal3 s 64600 7280 65000 7336 6 wbs_dat_o[8]
port 474 nsew signal output
rlabel metal3 s 64600 7728 65000 7784 6 wbs_dat_o[9]
port 475 nsew signal output
rlabel metal3 s 64600 18928 65000 18984 6 wbs_stb_i
port 476 nsew signal input
rlabel metal3 s 64600 18032 65000 18088 6 wbs_we_i
port 477 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 65000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8791238
string GDS_FILE /media/lucah/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1-multi/openlane/Multiplexer/runs/23_11_07_14_03/results/signoff/multiplexer.magic.gds
string GDS_START 395946
<< end >>

