magic
tech gf180mcuD
magscale 1 5
timestamp 1753965386
<< nwell >>
rect 629 1525 56827 58451
<< obsm1 >>
rect 672 1538 56784 58505
<< metal2 >>
rect 3248 59600 3304 60000
rect 4032 59600 4088 60000
rect 4816 59600 4872 60000
rect 5600 59600 5656 60000
rect 6384 59600 6440 60000
rect 7168 59600 7224 60000
rect 7952 59600 8008 60000
rect 8736 59600 8792 60000
rect 9520 59600 9576 60000
rect 10304 59600 10360 60000
rect 11088 59600 11144 60000
rect 11872 59600 11928 60000
rect 12656 59600 12712 60000
rect 13440 59600 13496 60000
rect 14224 59600 14280 60000
rect 15008 59600 15064 60000
rect 15792 59600 15848 60000
rect 16576 59600 16632 60000
rect 17360 59600 17416 60000
rect 18144 59600 18200 60000
rect 18928 59600 18984 60000
rect 19712 59600 19768 60000
rect 20496 59600 20552 60000
rect 21280 59600 21336 60000
rect 22064 59600 22120 60000
rect 22848 59600 22904 60000
rect 23632 59600 23688 60000
rect 24416 59600 24472 60000
rect 25200 59600 25256 60000
rect 25984 59600 26040 60000
rect 26768 59600 26824 60000
rect 27552 59600 27608 60000
rect 28336 59600 28392 60000
rect 29120 59600 29176 60000
rect 29904 59600 29960 60000
rect 30688 59600 30744 60000
rect 31472 59600 31528 60000
rect 32256 59600 32312 60000
rect 33040 59600 33096 60000
rect 33824 59600 33880 60000
rect 34608 59600 34664 60000
rect 35392 59600 35448 60000
rect 36176 59600 36232 60000
rect 36960 59600 37016 60000
rect 37744 59600 37800 60000
rect 38528 59600 38584 60000
rect 39312 59600 39368 60000
rect 40096 59600 40152 60000
rect 40880 59600 40936 60000
rect 41664 59600 41720 60000
rect 42448 59600 42504 60000
rect 43232 59600 43288 60000
rect 44016 59600 44072 60000
rect 44800 59600 44856 60000
rect 45584 59600 45640 60000
rect 46368 59600 46424 60000
rect 47152 59600 47208 60000
rect 47936 59600 47992 60000
rect 48720 59600 48776 60000
rect 49504 59600 49560 60000
rect 50288 59600 50344 60000
rect 51072 59600 51128 60000
rect 51856 59600 51912 60000
rect 52640 59600 52696 60000
rect 53424 59600 53480 60000
rect 54208 59600 54264 60000
<< obsm2 >>
rect 14 59570 3218 59682
rect 3334 59570 4002 59682
rect 4118 59570 4786 59682
rect 4902 59570 5570 59682
rect 5686 59570 6354 59682
rect 6470 59570 7138 59682
rect 7254 59570 7922 59682
rect 8038 59570 8706 59682
rect 8822 59570 9490 59682
rect 9606 59570 10274 59682
rect 10390 59570 11058 59682
rect 11174 59570 11842 59682
rect 11958 59570 12626 59682
rect 12742 59570 13410 59682
rect 13526 59570 14194 59682
rect 14310 59570 14978 59682
rect 15094 59570 15762 59682
rect 15878 59570 16546 59682
rect 16662 59570 17330 59682
rect 17446 59570 18114 59682
rect 18230 59570 18898 59682
rect 19014 59570 19682 59682
rect 19798 59570 20466 59682
rect 20582 59570 21250 59682
rect 21366 59570 22034 59682
rect 22150 59570 22818 59682
rect 22934 59570 23602 59682
rect 23718 59570 24386 59682
rect 24502 59570 25170 59682
rect 25286 59570 25954 59682
rect 26070 59570 26738 59682
rect 26854 59570 27522 59682
rect 27638 59570 28306 59682
rect 28422 59570 29090 59682
rect 29206 59570 29874 59682
rect 29990 59570 30658 59682
rect 30774 59570 31442 59682
rect 31558 59570 32226 59682
rect 32342 59570 33010 59682
rect 33126 59570 33794 59682
rect 33910 59570 34578 59682
rect 34694 59570 35362 59682
rect 35478 59570 36146 59682
rect 36262 59570 36930 59682
rect 37046 59570 37714 59682
rect 37830 59570 38498 59682
rect 38614 59570 39282 59682
rect 39398 59570 40066 59682
rect 40182 59570 40850 59682
rect 40966 59570 41634 59682
rect 41750 59570 42418 59682
rect 42534 59570 43202 59682
rect 43318 59570 43986 59682
rect 44102 59570 44770 59682
rect 44886 59570 45554 59682
rect 45670 59570 46338 59682
rect 46454 59570 47122 59682
rect 47238 59570 47906 59682
rect 48022 59570 48690 59682
rect 48806 59570 49474 59682
rect 49590 59570 50258 59682
rect 50374 59570 51042 59682
rect 51158 59570 51826 59682
rect 51942 59570 52610 59682
rect 52726 59570 53394 59682
rect 53510 59570 54178 59682
rect 54294 59570 56770 59682
rect 14 1549 56770 59570
<< metal3 >>
rect 0 57680 400 57736
rect 57100 57680 57500 57736
rect 57100 56672 57500 56728
rect 0 56000 400 56056
rect 57100 55664 57500 55720
rect 57100 54656 57500 54712
rect 0 54320 400 54376
rect 57100 53648 57500 53704
rect 0 52640 400 52696
rect 57100 52640 57500 52696
rect 57100 51632 57500 51688
rect 0 50960 400 51016
rect 57100 50624 57500 50680
rect 57100 49616 57500 49672
rect 0 49280 400 49336
rect 57100 48608 57500 48664
rect 0 47600 400 47656
rect 57100 47600 57500 47656
rect 57100 46592 57500 46648
rect 0 45920 400 45976
rect 57100 45584 57500 45640
rect 57100 44576 57500 44632
rect 0 44240 400 44296
rect 57100 43568 57500 43624
rect 0 42560 400 42616
rect 57100 42560 57500 42616
rect 57100 41552 57500 41608
rect 0 40880 400 40936
rect 57100 40544 57500 40600
rect 57100 39536 57500 39592
rect 0 39200 400 39256
rect 57100 38528 57500 38584
rect 0 37520 400 37576
rect 57100 37520 57500 37576
rect 57100 36512 57500 36568
rect 0 35840 400 35896
rect 57100 35504 57500 35560
rect 57100 34496 57500 34552
rect 0 34160 400 34216
rect 57100 33488 57500 33544
rect 0 32480 400 32536
rect 57100 32480 57500 32536
rect 57100 31472 57500 31528
rect 0 30800 400 30856
rect 57100 30464 57500 30520
rect 57100 29456 57500 29512
rect 0 29120 400 29176
rect 57100 28448 57500 28504
rect 0 27440 400 27496
rect 57100 27440 57500 27496
rect 57100 26432 57500 26488
rect 0 25760 400 25816
rect 57100 25424 57500 25480
rect 57100 24416 57500 24472
rect 0 24080 400 24136
rect 57100 23408 57500 23464
rect 0 22400 400 22456
rect 57100 22400 57500 22456
rect 57100 21392 57500 21448
rect 0 20720 400 20776
rect 57100 20384 57500 20440
rect 57100 19376 57500 19432
rect 0 19040 400 19096
rect 57100 18368 57500 18424
rect 0 17360 400 17416
rect 57100 17360 57500 17416
rect 57100 16352 57500 16408
rect 0 15680 400 15736
rect 57100 15344 57500 15400
rect 57100 14336 57500 14392
rect 0 14000 400 14056
rect 57100 13328 57500 13384
rect 0 12320 400 12376
rect 57100 12320 57500 12376
rect 57100 11312 57500 11368
rect 0 10640 400 10696
rect 57100 10304 57500 10360
rect 57100 9296 57500 9352
rect 0 8960 400 9016
rect 57100 8288 57500 8344
rect 0 7280 400 7336
rect 57100 7280 57500 7336
rect 57100 6272 57500 6328
rect 0 5600 400 5656
rect 57100 5264 57500 5320
rect 57100 4256 57500 4312
rect 0 3920 400 3976
rect 57100 3248 57500 3304
rect 0 2240 400 2296
rect 57100 2240 57500 2296
<< obsm3 >>
rect 9 57766 57162 59066
rect 430 57650 57070 57766
rect 9 56758 57162 57650
rect 9 56642 57070 56758
rect 9 56086 57162 56642
rect 430 55970 57162 56086
rect 9 55750 57162 55970
rect 9 55634 57070 55750
rect 9 54742 57162 55634
rect 9 54626 57070 54742
rect 9 54406 57162 54626
rect 430 54290 57162 54406
rect 9 53734 57162 54290
rect 9 53618 57070 53734
rect 9 52726 57162 53618
rect 430 52610 57070 52726
rect 9 51718 57162 52610
rect 9 51602 57070 51718
rect 9 51046 57162 51602
rect 430 50930 57162 51046
rect 9 50710 57162 50930
rect 9 50594 57070 50710
rect 9 49702 57162 50594
rect 9 49586 57070 49702
rect 9 49366 57162 49586
rect 430 49250 57162 49366
rect 9 48694 57162 49250
rect 9 48578 57070 48694
rect 9 47686 57162 48578
rect 430 47570 57070 47686
rect 9 46678 57162 47570
rect 9 46562 57070 46678
rect 9 46006 57162 46562
rect 430 45890 57162 46006
rect 9 45670 57162 45890
rect 9 45554 57070 45670
rect 9 44662 57162 45554
rect 9 44546 57070 44662
rect 9 44326 57162 44546
rect 430 44210 57162 44326
rect 9 43654 57162 44210
rect 9 43538 57070 43654
rect 9 42646 57162 43538
rect 430 42530 57070 42646
rect 9 41638 57162 42530
rect 9 41522 57070 41638
rect 9 40966 57162 41522
rect 430 40850 57162 40966
rect 9 40630 57162 40850
rect 9 40514 57070 40630
rect 9 39622 57162 40514
rect 9 39506 57070 39622
rect 9 39286 57162 39506
rect 430 39170 57162 39286
rect 9 38614 57162 39170
rect 9 38498 57070 38614
rect 9 37606 57162 38498
rect 430 37490 57070 37606
rect 9 36598 57162 37490
rect 9 36482 57070 36598
rect 9 35926 57162 36482
rect 430 35810 57162 35926
rect 9 35590 57162 35810
rect 9 35474 57070 35590
rect 9 34582 57162 35474
rect 9 34466 57070 34582
rect 9 34246 57162 34466
rect 430 34130 57162 34246
rect 9 33574 57162 34130
rect 9 33458 57070 33574
rect 9 32566 57162 33458
rect 430 32450 57070 32566
rect 9 31558 57162 32450
rect 9 31442 57070 31558
rect 9 30886 57162 31442
rect 430 30770 57162 30886
rect 9 30550 57162 30770
rect 9 30434 57070 30550
rect 9 29542 57162 30434
rect 9 29426 57070 29542
rect 9 29206 57162 29426
rect 430 29090 57162 29206
rect 9 28534 57162 29090
rect 9 28418 57070 28534
rect 9 27526 57162 28418
rect 430 27410 57070 27526
rect 9 26518 57162 27410
rect 9 26402 57070 26518
rect 9 25846 57162 26402
rect 430 25730 57162 25846
rect 9 25510 57162 25730
rect 9 25394 57070 25510
rect 9 24502 57162 25394
rect 9 24386 57070 24502
rect 9 24166 57162 24386
rect 430 24050 57162 24166
rect 9 23494 57162 24050
rect 9 23378 57070 23494
rect 9 22486 57162 23378
rect 430 22370 57070 22486
rect 9 21478 57162 22370
rect 9 21362 57070 21478
rect 9 20806 57162 21362
rect 430 20690 57162 20806
rect 9 20470 57162 20690
rect 9 20354 57070 20470
rect 9 19462 57162 20354
rect 9 19346 57070 19462
rect 9 19126 57162 19346
rect 430 19010 57162 19126
rect 9 18454 57162 19010
rect 9 18338 57070 18454
rect 9 17446 57162 18338
rect 430 17330 57070 17446
rect 9 16438 57162 17330
rect 9 16322 57070 16438
rect 9 15766 57162 16322
rect 430 15650 57162 15766
rect 9 15430 57162 15650
rect 9 15314 57070 15430
rect 9 14422 57162 15314
rect 9 14306 57070 14422
rect 9 14086 57162 14306
rect 430 13970 57162 14086
rect 9 13414 57162 13970
rect 9 13298 57070 13414
rect 9 12406 57162 13298
rect 430 12290 57070 12406
rect 9 11398 57162 12290
rect 9 11282 57070 11398
rect 9 10726 57162 11282
rect 430 10610 57162 10726
rect 9 10390 57162 10610
rect 9 10274 57070 10390
rect 9 9382 57162 10274
rect 9 9266 57070 9382
rect 9 9046 57162 9266
rect 430 8930 57162 9046
rect 9 8374 57162 8930
rect 9 8258 57070 8374
rect 9 7366 57162 8258
rect 430 7250 57070 7366
rect 9 6358 57162 7250
rect 9 6242 57070 6358
rect 9 5686 57162 6242
rect 430 5570 57162 5686
rect 9 5350 57162 5570
rect 9 5234 57070 5350
rect 9 4342 57162 5234
rect 9 4226 57070 4342
rect 9 4006 57162 4226
rect 430 3890 57162 4006
rect 9 3334 57162 3890
rect 9 3218 57070 3334
rect 9 2326 57162 3218
rect 430 2210 57070 2326
rect 9 1554 57162 2210
<< metal4 >>
rect 2224 1538 2384 58438
rect 9904 1538 10064 58438
rect 17584 1538 17744 58438
rect 25264 1538 25424 58438
rect 32944 1538 33104 58438
rect 40624 1538 40784 58438
rect 48304 1538 48464 58438
rect 55984 1538 56144 58438
<< obsm4 >>
rect 4270 58468 56266 58847
rect 4270 8073 9874 58468
rect 10094 8073 17554 58468
rect 17774 8073 25234 58468
rect 25454 8073 32914 58468
rect 33134 8073 40594 58468
rect 40814 8073 48274 58468
rect 48494 8073 55954 58468
rect 56174 8073 56266 58468
<< labels >>
rlabel metal3 s 0 5600 400 5656 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 0 22400 400 22456 6 custom_settings[10]
port 2 nsew signal input
rlabel metal3 s 0 24080 400 24136 6 custom_settings[11]
port 3 nsew signal input
rlabel metal3 s 0 25760 400 25816 6 custom_settings[12]
port 4 nsew signal input
rlabel metal3 s 0 27440 400 27496 6 custom_settings[13]
port 5 nsew signal input
rlabel metal3 s 0 29120 400 29176 6 custom_settings[14]
port 6 nsew signal input
rlabel metal3 s 0 30800 400 30856 6 custom_settings[15]
port 7 nsew signal input
rlabel metal3 s 0 32480 400 32536 6 custom_settings[16]
port 8 nsew signal input
rlabel metal3 s 0 34160 400 34216 6 custom_settings[17]
port 9 nsew signal input
rlabel metal3 s 0 35840 400 35896 6 custom_settings[18]
port 10 nsew signal input
rlabel metal3 s 0 37520 400 37576 6 custom_settings[19]
port 11 nsew signal input
rlabel metal3 s 0 7280 400 7336 6 custom_settings[1]
port 12 nsew signal input
rlabel metal3 s 0 39200 400 39256 6 custom_settings[20]
port 13 nsew signal input
rlabel metal3 s 0 40880 400 40936 6 custom_settings[21]
port 14 nsew signal input
rlabel metal3 s 0 42560 400 42616 6 custom_settings[22]
port 15 nsew signal input
rlabel metal3 s 0 44240 400 44296 6 custom_settings[23]
port 16 nsew signal input
rlabel metal3 s 0 45920 400 45976 6 custom_settings[24]
port 17 nsew signal input
rlabel metal3 s 0 47600 400 47656 6 custom_settings[25]
port 18 nsew signal input
rlabel metal3 s 0 49280 400 49336 6 custom_settings[26]
port 19 nsew signal input
rlabel metal3 s 0 50960 400 51016 6 custom_settings[27]
port 20 nsew signal input
rlabel metal3 s 0 52640 400 52696 6 custom_settings[28]
port 21 nsew signal input
rlabel metal3 s 0 54320 400 54376 6 custom_settings[29]
port 22 nsew signal input
rlabel metal3 s 0 8960 400 9016 6 custom_settings[2]
port 23 nsew signal input
rlabel metal3 s 0 56000 400 56056 6 custom_settings[30]
port 24 nsew signal input
rlabel metal3 s 0 57680 400 57736 6 custom_settings[31]
port 25 nsew signal input
rlabel metal3 s 0 10640 400 10696 6 custom_settings[3]
port 26 nsew signal input
rlabel metal3 s 0 12320 400 12376 6 custom_settings[4]
port 27 nsew signal input
rlabel metal3 s 0 14000 400 14056 6 custom_settings[5]
port 28 nsew signal input
rlabel metal3 s 0 15680 400 15736 6 custom_settings[6]
port 29 nsew signal input
rlabel metal3 s 0 17360 400 17416 6 custom_settings[7]
port 30 nsew signal input
rlabel metal3 s 0 19040 400 19096 6 custom_settings[8]
port 31 nsew signal input
rlabel metal3 s 0 20720 400 20776 6 custom_settings[9]
port 32 nsew signal input
rlabel metal2 s 3248 59600 3304 60000 6 io_in[0]
port 33 nsew signal input
rlabel metal2 s 11088 59600 11144 60000 6 io_in[10]
port 34 nsew signal input
rlabel metal2 s 11872 59600 11928 60000 6 io_in[11]
port 35 nsew signal input
rlabel metal2 s 12656 59600 12712 60000 6 io_in[12]
port 36 nsew signal input
rlabel metal2 s 13440 59600 13496 60000 6 io_in[13]
port 37 nsew signal input
rlabel metal2 s 14224 59600 14280 60000 6 io_in[14]
port 38 nsew signal input
rlabel metal2 s 15008 59600 15064 60000 6 io_in[15]
port 39 nsew signal input
rlabel metal2 s 15792 59600 15848 60000 6 io_in[16]
port 40 nsew signal input
rlabel metal2 s 16576 59600 16632 60000 6 io_in[17]
port 41 nsew signal input
rlabel metal2 s 17360 59600 17416 60000 6 io_in[18]
port 42 nsew signal input
rlabel metal2 s 18144 59600 18200 60000 6 io_in[19]
port 43 nsew signal input
rlabel metal2 s 4032 59600 4088 60000 6 io_in[1]
port 44 nsew signal input
rlabel metal2 s 18928 59600 18984 60000 6 io_in[20]
port 45 nsew signal input
rlabel metal2 s 19712 59600 19768 60000 6 io_in[21]
port 46 nsew signal input
rlabel metal2 s 20496 59600 20552 60000 6 io_in[22]
port 47 nsew signal input
rlabel metal2 s 21280 59600 21336 60000 6 io_in[23]
port 48 nsew signal input
rlabel metal2 s 22064 59600 22120 60000 6 io_in[24]
port 49 nsew signal input
rlabel metal2 s 22848 59600 22904 60000 6 io_in[25]
port 50 nsew signal input
rlabel metal2 s 23632 59600 23688 60000 6 io_in[26]
port 51 nsew signal input
rlabel metal2 s 24416 59600 24472 60000 6 io_in[27]
port 52 nsew signal input
rlabel metal2 s 25200 59600 25256 60000 6 io_in[28]
port 53 nsew signal input
rlabel metal2 s 25984 59600 26040 60000 6 io_in[29]
port 54 nsew signal input
rlabel metal2 s 4816 59600 4872 60000 6 io_in[2]
port 55 nsew signal input
rlabel metal2 s 26768 59600 26824 60000 6 io_in[30]
port 56 nsew signal input
rlabel metal2 s 27552 59600 27608 60000 6 io_in[31]
port 57 nsew signal input
rlabel metal2 s 28336 59600 28392 60000 6 io_in[32]
port 58 nsew signal input
rlabel metal2 s 5600 59600 5656 60000 6 io_in[3]
port 59 nsew signal input
rlabel metal2 s 6384 59600 6440 60000 6 io_in[4]
port 60 nsew signal input
rlabel metal2 s 7168 59600 7224 60000 6 io_in[5]
port 61 nsew signal input
rlabel metal2 s 7952 59600 8008 60000 6 io_in[6]
port 62 nsew signal input
rlabel metal2 s 8736 59600 8792 60000 6 io_in[7]
port 63 nsew signal input
rlabel metal2 s 9520 59600 9576 60000 6 io_in[8]
port 64 nsew signal input
rlabel metal2 s 10304 59600 10360 60000 6 io_in[9]
port 65 nsew signal input
rlabel metal3 s 57100 2240 57500 2296 6 io_oeb[0]
port 66 nsew signal output
rlabel metal3 s 57100 12320 57500 12376 6 io_oeb[10]
port 67 nsew signal output
rlabel metal3 s 57100 13328 57500 13384 6 io_oeb[11]
port 68 nsew signal output
rlabel metal3 s 57100 14336 57500 14392 6 io_oeb[12]
port 69 nsew signal output
rlabel metal3 s 57100 15344 57500 15400 6 io_oeb[13]
port 70 nsew signal output
rlabel metal3 s 57100 16352 57500 16408 6 io_oeb[14]
port 71 nsew signal output
rlabel metal3 s 57100 17360 57500 17416 6 io_oeb[15]
port 72 nsew signal output
rlabel metal3 s 57100 18368 57500 18424 6 io_oeb[16]
port 73 nsew signal output
rlabel metal3 s 57100 19376 57500 19432 6 io_oeb[17]
port 74 nsew signal output
rlabel metal3 s 57100 20384 57500 20440 6 io_oeb[18]
port 75 nsew signal output
rlabel metal3 s 57100 21392 57500 21448 6 io_oeb[19]
port 76 nsew signal output
rlabel metal3 s 57100 3248 57500 3304 6 io_oeb[1]
port 77 nsew signal output
rlabel metal3 s 57100 22400 57500 22456 6 io_oeb[20]
port 78 nsew signal output
rlabel metal3 s 57100 23408 57500 23464 6 io_oeb[21]
port 79 nsew signal output
rlabel metal3 s 57100 24416 57500 24472 6 io_oeb[22]
port 80 nsew signal output
rlabel metal3 s 57100 25424 57500 25480 6 io_oeb[23]
port 81 nsew signal output
rlabel metal3 s 57100 26432 57500 26488 6 io_oeb[24]
port 82 nsew signal output
rlabel metal3 s 57100 27440 57500 27496 6 io_oeb[25]
port 83 nsew signal output
rlabel metal3 s 57100 28448 57500 28504 6 io_oeb[26]
port 84 nsew signal output
rlabel metal3 s 57100 29456 57500 29512 6 io_oeb[27]
port 85 nsew signal output
rlabel metal3 s 57100 30464 57500 30520 6 io_oeb[28]
port 86 nsew signal output
rlabel metal3 s 57100 31472 57500 31528 6 io_oeb[29]
port 87 nsew signal output
rlabel metal3 s 57100 4256 57500 4312 6 io_oeb[2]
port 88 nsew signal output
rlabel metal3 s 57100 32480 57500 32536 6 io_oeb[30]
port 89 nsew signal output
rlabel metal3 s 57100 33488 57500 33544 6 io_oeb[31]
port 90 nsew signal output
rlabel metal3 s 57100 34496 57500 34552 6 io_oeb[32]
port 91 nsew signal output
rlabel metal3 s 57100 5264 57500 5320 6 io_oeb[3]
port 92 nsew signal output
rlabel metal3 s 57100 6272 57500 6328 6 io_oeb[4]
port 93 nsew signal output
rlabel metal3 s 57100 7280 57500 7336 6 io_oeb[5]
port 94 nsew signal output
rlabel metal3 s 57100 8288 57500 8344 6 io_oeb[6]
port 95 nsew signal output
rlabel metal3 s 57100 9296 57500 9352 6 io_oeb[7]
port 96 nsew signal output
rlabel metal3 s 57100 10304 57500 10360 6 io_oeb[8]
port 97 nsew signal output
rlabel metal3 s 57100 11312 57500 11368 6 io_oeb[9]
port 98 nsew signal output
rlabel metal2 s 29120 59600 29176 60000 6 io_out[0]
port 99 nsew signal output
rlabel metal2 s 36960 59600 37016 60000 6 io_out[10]
port 100 nsew signal output
rlabel metal2 s 37744 59600 37800 60000 6 io_out[11]
port 101 nsew signal output
rlabel metal2 s 38528 59600 38584 60000 6 io_out[12]
port 102 nsew signal output
rlabel metal2 s 39312 59600 39368 60000 6 io_out[13]
port 103 nsew signal output
rlabel metal2 s 40096 59600 40152 60000 6 io_out[14]
port 104 nsew signal output
rlabel metal2 s 40880 59600 40936 60000 6 io_out[15]
port 105 nsew signal output
rlabel metal2 s 41664 59600 41720 60000 6 io_out[16]
port 106 nsew signal output
rlabel metal2 s 42448 59600 42504 60000 6 io_out[17]
port 107 nsew signal output
rlabel metal2 s 43232 59600 43288 60000 6 io_out[18]
port 108 nsew signal output
rlabel metal2 s 44016 59600 44072 60000 6 io_out[19]
port 109 nsew signal output
rlabel metal2 s 29904 59600 29960 60000 6 io_out[1]
port 110 nsew signal output
rlabel metal2 s 44800 59600 44856 60000 6 io_out[20]
port 111 nsew signal output
rlabel metal2 s 45584 59600 45640 60000 6 io_out[21]
port 112 nsew signal output
rlabel metal2 s 46368 59600 46424 60000 6 io_out[22]
port 113 nsew signal output
rlabel metal2 s 47152 59600 47208 60000 6 io_out[23]
port 114 nsew signal output
rlabel metal2 s 47936 59600 47992 60000 6 io_out[24]
port 115 nsew signal output
rlabel metal2 s 48720 59600 48776 60000 6 io_out[25]
port 116 nsew signal output
rlabel metal2 s 49504 59600 49560 60000 6 io_out[26]
port 117 nsew signal output
rlabel metal2 s 50288 59600 50344 60000 6 io_out[27]
port 118 nsew signal output
rlabel metal2 s 51072 59600 51128 60000 6 io_out[28]
port 119 nsew signal output
rlabel metal2 s 51856 59600 51912 60000 6 io_out[29]
port 120 nsew signal output
rlabel metal2 s 30688 59600 30744 60000 6 io_out[2]
port 121 nsew signal output
rlabel metal2 s 52640 59600 52696 60000 6 io_out[30]
port 122 nsew signal output
rlabel metal2 s 53424 59600 53480 60000 6 io_out[31]
port 123 nsew signal output
rlabel metal2 s 54208 59600 54264 60000 6 io_out[32]
port 124 nsew signal output
rlabel metal2 s 31472 59600 31528 60000 6 io_out[3]
port 125 nsew signal output
rlabel metal2 s 32256 59600 32312 60000 6 io_out[4]
port 126 nsew signal output
rlabel metal2 s 33040 59600 33096 60000 6 io_out[5]
port 127 nsew signal output
rlabel metal2 s 33824 59600 33880 60000 6 io_out[6]
port 128 nsew signal output
rlabel metal2 s 34608 59600 34664 60000 6 io_out[7]
port 129 nsew signal output
rlabel metal2 s 35392 59600 35448 60000 6 io_out[8]
port 130 nsew signal output
rlabel metal2 s 36176 59600 36232 60000 6 io_out[9]
port 131 nsew signal output
rlabel metal3 s 0 3920 400 3976 6 rst_n
port 132 nsew signal input
rlabel metal3 s 57100 35504 57500 35560 6 sram_addr[0]
port 133 nsew signal output
rlabel metal3 s 57100 36512 57500 36568 6 sram_addr[1]
port 134 nsew signal output
rlabel metal3 s 57100 37520 57500 37576 6 sram_addr[2]
port 135 nsew signal output
rlabel metal3 s 57100 38528 57500 38584 6 sram_addr[3]
port 136 nsew signal output
rlabel metal3 s 57100 39536 57500 39592 6 sram_addr[4]
port 137 nsew signal output
rlabel metal3 s 57100 40544 57500 40600 6 sram_addr[5]
port 138 nsew signal output
rlabel metal3 s 57100 57680 57500 57736 6 sram_gwe
port 139 nsew signal output
rlabel metal3 s 57100 41552 57500 41608 6 sram_in[0]
port 140 nsew signal output
rlabel metal3 s 57100 42560 57500 42616 6 sram_in[1]
port 141 nsew signal output
rlabel metal3 s 57100 43568 57500 43624 6 sram_in[2]
port 142 nsew signal output
rlabel metal3 s 57100 44576 57500 44632 6 sram_in[3]
port 143 nsew signal output
rlabel metal3 s 57100 45584 57500 45640 6 sram_in[4]
port 144 nsew signal output
rlabel metal3 s 57100 46592 57500 46648 6 sram_in[5]
port 145 nsew signal output
rlabel metal3 s 57100 47600 57500 47656 6 sram_in[6]
port 146 nsew signal output
rlabel metal3 s 57100 48608 57500 48664 6 sram_in[7]
port 147 nsew signal output
rlabel metal3 s 57100 49616 57500 49672 6 sram_out[0]
port 148 nsew signal input
rlabel metal3 s 57100 50624 57500 50680 6 sram_out[1]
port 149 nsew signal input
rlabel metal3 s 57100 51632 57500 51688 6 sram_out[2]
port 150 nsew signal input
rlabel metal3 s 57100 52640 57500 52696 6 sram_out[3]
port 151 nsew signal input
rlabel metal3 s 57100 53648 57500 53704 6 sram_out[4]
port 152 nsew signal input
rlabel metal3 s 57100 54656 57500 54712 6 sram_out[5]
port 153 nsew signal input
rlabel metal3 s 57100 55664 57500 55720 6 sram_out[6]
port 154 nsew signal input
rlabel metal3 s 57100 56672 57500 56728 6 sram_out[7]
port 155 nsew signal input
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 156 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58438 6 vdd
port 156 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58438 6 vdd
port 156 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58438 6 vdd
port 156 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58438 6 vss
port 157 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58438 6 vss
port 157 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58438 6 vss
port 157 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 58438 6 vss
port 157 nsew ground bidirectional
rlabel metal3 s 0 2240 400 2296 6 wb_clk_i
port 158 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 57500 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 11220642
string GDS_FILE /home/lucah/gfmpw1-multi/openlane/wrapped_qcpu/runs/25_07_31_14_26/results/signoff/wrapped_qcpu.magic.gds
string GDS_START 272602
<< end >>

